$date
  Wed May 16 15:12:29 2018
$end
$version
  GHDL v0
$end
$timescale
  1 fs
$end
$var reg 1 ! clk $end
$var reg 1 " reset $end
$var reg 1 # detectedbit $end
$var reg 8 $ bitinput[7:0] $end
$scope module detector $end
$var reg 1 % clk $end
$var reg 1 & reset $end
$var reg 8 ' bitinput[7:0] $end
$var reg 1 ( detectedbit $end
$comment state is not handled $end
$var reg 1 ) auxbit1 $end
$var reg 1 * auxbit $end
$scope module memcompare1 $end
$var reg 8 + charinput[7:0] $end
$var integer 32 , address $end
$var reg 1 - iscorrect $end
$var reg 8 . auxdata[7:0] $end
$scope module rom $end
$var integer 32 / address $end
$var reg 8 0 data[7:0] $end
$upscope $end
$scope module comparador $end
$var reg 8 1 charinputa[7:0] $end
$var reg 8 2 charinputb[7:0] $end
$var reg 1 3 bitoutput $end
$var reg 1 4 a1 $end
$var reg 1 5 a2 $end
$var reg 1 6 a3 $end
$var reg 1 7 a4 $end
$var reg 1 8 a5 $end
$var reg 1 9 a6 $end
$var reg 1 : a7 $end
$var reg 1 ; a8 $end
$upscope $end
$upscope $end
$scope module memcompare2 $end
$var reg 8 < charinput[7:0] $end
$var integer 32 = address $end
$var reg 1 > iscorrect $end
$var reg 8 ? auxdata[7:0] $end
$scope module rom $end
$var integer 32 @ address $end
$var reg 8 A data[7:0] $end
$upscope $end
$scope module comparador $end
$var reg 8 B charinputa[7:0] $end
$var reg 8 C charinputb[7:0] $end
$var reg 1 D bitoutput $end
$var reg 1 E a1 $end
$var reg 1 F a2 $end
$var reg 1 G a3 $end
$var reg 1 H a4 $end
$var reg 1 I a5 $end
$var reg 1 J a6 $end
$var reg 1 K a7 $end
$var reg 1 L a8 $end
$upscope $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
0!
0"
U#
b00000000 $
0%
0&
b00000000 '
U(
0)
0*
b00000000 +
b1000 ,
0-
b01101001 .
b1000 /
b01101001 0
b00000000 1
b01101001 2
03
04
15
16
07
18
09
0:
1;
b00000000 <
b10010 =
0>
b01110011 ?
b10010 @
b01110011 A
b00000000 B
b01110011 C
0D
0E
0F
1G
1H
0I
0J
0K
1L
#5000000
1!
0#
1%
0(
#10000000
0!
b00010000 $
0%
b00010000 '
b00010000 +
b00010000 1
08
b00010000 <
b00010000 B
1I
#15000000
1!
1%
#20000000
0!
b01101001 $
0%
b01101001 '
1*
b01101001 +
1-
b01101001 1
13
14
17
18
19
1:
b01101001 <
b01101001 B
1E
0H
0I
1J
1K
#25000000
1!
1%
#30000000
0!
b01110011 $
0%
b01110011 '
1)
0*
b01110011 +
0-
b01110011 1
03
05
07
08
b01110011 <
1>
b01110011 B
1D
1F
1H
1I
#35000000
1!
1#
1%
1(
#40000000
0!
0%
#45000000
1!
0#
1%
0(
#50000000
0!
b00010001 $
0%
b00010001 '
0)
b00010001 +
b00010001 1
15
09
0:
b00010001 <
0>
b00010001 B
0D
0F
0J
0K
#55000000
1!
1%
#60000000
0!
b00010000 $
0%
b00010000 '
b00010000 +
b00010000 1
04
b00010000 <
b00010000 B
0E
#65000000
1!
1%
#70000000
0!
b01100001 $
0%
b01100001 '
b01100001 +
b01100001 1
14
18
19
1:
b01100001 <
b01100001 B
1E
0I
1J
1K
#75000000
1!
1%
#80000000
0!
b00000011 $
0%
b00000011 '
b00000011 +
b00000011 1
05
09
0:
b00000011 <
b00000011 B
1F
0J
0K
#85000000
1!
1%
#90000000
0!
b00000000 $
0%
b00000000 '
b00000000 +
b00000000 1
04
15
b00000000 <
b00000000 B
0E
0F
#95000000
1!
1%
#100000000
0!
0%
#105000000
1!
1%
#110000000
0!
0%
#115000000
1!
1%
#120000000
0!
0%
#125000000
1!
1%
#130000000
0!
0%
#135000000
1!
1%
#140000000
0!
0%
#145000000
1!
1%
#150000000
0!
0%
#155000000
1!
1%
#160000000
0!
0%
#165000000
1!
1%
#170000000
0!
0%
#175000000
1!
1%
#180000000
0!
0%
#185000000
1!
1%
#190000000
0!
0%
#195000000
1!
1%
#200000000
0!
0%
#205000000
1!
1%
#210000000
0!
0%
#215000000
1!
1%
#220000000
0!
0%
#225000000
1!
1%
#230000000
0!
0%
#235000000
1!
1%
#240000000
0!
0%
#245000000
1!
1%
#250000000
0!
0%
#255000000
1!
1%
#260000000
0!
0%
#265000000
1!
1%
#270000000
0!
0%
#275000000
1!
1%
#280000000
0!
0%
#285000000
1!
1%
#290000000
0!
0%
#295000000
1!
1%
#300000000
0!
0%
#305000000
1!
1%
#310000000
0!
0%
#315000000
1!
1%
#320000000
0!
0%
#325000000
1!
1%
#330000000
0!
0%
#335000000
1!
1%
#340000000
0!
0%
#345000000
1!
1%
#350000000
0!
0%
#355000000
1!
1%
#360000000
0!
0%
#365000000
1!
1%
#370000000
0!
0%
#375000000
1!
1%
#380000000
0!
0%
#385000000
1!
1%
#390000000
0!
0%
#395000000
1!
1%
#400000000
0!
0%
#405000000
1!
1%
#410000000
0!
0%
#415000000
1!
1%
#420000000
0!
0%
#425000000
1!
1%
#430000000
0!
0%
#435000000
1!
1%
#440000000
0!
0%
#445000000
1!
1%
#450000000
0!
0%
#455000000
1!
1%
#460000000
0!
0%
#465000000
1!
1%
#470000000
0!
0%
#475000000
1!
1%
#480000000
0!
0%
#485000000
1!
1%
#490000000
0!
0%
#495000000
1!
1%
#500000000
0!
0%
#505000000
1!
1%
#510000000
0!
0%
#515000000
1!
1%
#520000000
0!
0%
#525000000
1!
1%
#530000000
0!
0%
#535000000
1!
1%
#540000000
0!
0%
#545000000
1!
1%
#550000000
0!
0%
#555000000
1!
1%
#560000000
0!
0%
#565000000
1!
1%
#570000000
0!
0%
#575000000
1!
1%
#580000000
0!
0%
#585000000
1!
1%
#590000000
0!
0%
#595000000
1!
1%
#600000000
0!
0%
#605000000
1!
1%
#610000000
0!
0%
#615000000
1!
1%
#620000000
0!
0%
#625000000
1!
1%
#630000000
0!
0%
#635000000
1!
1%
#640000000
0!
0%
#645000000
1!
1%
#650000000
0!
0%
#655000000
1!
1%
#660000000
0!
0%
#665000000
1!
1%
#670000000
0!
0%
#675000000
1!
1%
#680000000
0!
0%
#685000000
1!
1%
#690000000
0!
0%
#695000000
1!
1%
#700000000
0!
0%
#705000000
1!
1%
#710000000
0!
0%
#715000000
1!
1%
#720000000
0!
0%
#725000000
1!
1%
#730000000
0!
0%
#735000000
1!
1%
#740000000
0!
0%
#745000000
1!
1%
#750000000
0!
0%
#755000000
1!
1%
#760000000
0!
0%
#765000000
1!
1%
#770000000
0!
0%
#775000000
1!
1%
#780000000
0!
0%
#785000000
1!
1%
#790000000
0!
0%
#795000000
1!
1%
#800000000
0!
0%
#805000000
1!
1%
#810000000
0!
0%
#815000000
1!
1%
#820000000
0!
0%
#825000000
1!
1%
#830000000
0!
0%
#835000000
1!
1%
#840000000
0!
0%
#845000000
1!
1%
#850000000
0!
0%
#855000000
1!
1%
#860000000
0!
0%
#865000000
1!
1%
#870000000
0!
0%
#875000000
1!
1%
#880000000
0!
0%
#885000000
1!
1%
#890000000
0!
0%
#895000000
1!
1%
#900000000
0!
0%
#905000000
1!
1%
#910000000
0!
0%
#915000000
1!
1%
#920000000
0!
0%
#925000000
1!
1%
#930000000
0!
0%
#935000000
1!
1%
#940000000
0!
0%
#945000000
1!
1%
#950000000
0!
0%
#955000000
1!
1%
#960000000
0!
0%
#965000000
1!
1%
#970000000
0!
0%
#975000000
1!
1%
#980000000
0!
0%
#985000000
1!
1%
#990000000
0!
0%
#995000000
1!
1%
#1000000000
0!
0%
#1005000000
1!
1%
#1010000000
0!
0%
#1015000000
1!
1%
#1020000000
0!
0%
#1025000000
1!
1%
#1030000000
0!
0%
#1035000000
1!
1%
#1040000000
0!
0%
#1045000000
1!
1%
#1050000000
0!
0%
#1055000000
1!
1%
#1060000000
0!
0%
#1065000000
1!
1%
#1070000000
0!
0%
#1075000000
1!
1%
#1080000000
0!
0%
#1085000000
1!
1%
#1090000000
0!
0%
#1095000000
1!
1%
#1100000000
0!
0%
#1105000000
1!
1%
#1110000000
0!
0%
#1115000000
1!
1%
#1120000000
0!
0%
#1125000000
1!
1%
#1130000000
0!
0%
#1135000000
1!
1%
#1140000000
0!
0%
#1145000000
1!
1%
#1150000000
0!
0%
#1155000000
1!
1%
#1160000000
0!
0%
#1165000000
1!
1%
#1170000000
0!
0%
#1175000000
1!
1%
#1180000000
0!
0%
#1185000000
1!
1%
#1190000000
0!
0%
#1195000000
1!
1%
#1200000000
0!
0%
#1205000000
1!
1%
#1210000000
0!
0%
#1215000000
1!
1%
#1220000000
0!
0%
#1225000000
1!
1%
#1230000000
0!
0%
#1235000000
1!
1%
#1240000000
0!
0%
#1245000000
1!
1%
#1250000000
0!
0%
#1255000000
1!
1%
#1260000000
0!
0%
#1265000000
1!
1%
#1270000000
0!
0%
#1275000000
1!
1%
#1280000000
0!
0%
#1285000000
1!
1%
#1290000000
0!
0%
#1295000000
1!
1%
#1300000000
0!
0%
#1305000000
1!
1%
#1310000000
0!
0%
#1315000000
1!
1%
#1320000000
0!
0%
#1325000000
1!
1%
#1330000000
0!
0%
#1335000000
1!
1%
#1340000000
0!
0%
#1345000000
1!
1%
#1350000000
0!
0%
#1355000000
1!
1%
#1360000000
0!
0%
#1365000000
1!
1%
#1370000000
0!
0%
#1375000000
1!
1%
#1380000000
0!
0%
#1385000000
1!
1%
#1390000000
0!
0%
#1395000000
1!
1%
#1400000000
0!
0%
#1405000000
1!
1%
#1410000000
0!
0%
#1415000000
1!
1%
#1420000000
0!
0%
#1425000000
1!
1%
#1430000000
0!
0%
#1435000000
1!
1%
#1440000000
0!
0%
#1445000000
1!
1%
#1450000000
0!
0%
#1455000000
1!
1%
#1460000000
0!
0%
#1465000000
1!
1%
#1470000000
0!
0%
#1475000000
1!
1%
#1480000000
0!
0%
#1485000000
1!
1%
#1490000000
0!
0%
#1495000000
1!
1%
#1500000000
0!
0%
#1505000000
1!
1%
#1510000000
0!
0%
#1515000000
1!
1%
#1520000000
0!
0%
#1525000000
1!
1%
#1530000000
0!
0%
#1535000000
1!
1%
#1540000000
0!
0%
#1545000000
1!
1%
#1550000000
0!
0%
#1555000000
1!
1%
#1560000000
0!
0%
#1565000000
1!
1%
#1570000000
0!
0%
#1575000000
1!
1%
#1580000000
0!
0%
#1585000000
1!
1%
#1590000000
0!
0%
#1595000000
1!
1%
#1600000000
0!
0%
#1605000000
1!
1%
#1610000000
0!
0%
#1615000000
1!
1%
#1620000000
0!
0%
#1625000000
1!
1%
#1630000000
0!
0%
#1635000000
1!
1%
#1640000000
0!
0%
#1645000000
1!
1%
#1650000000
0!
0%
#1655000000
1!
1%
#1660000000
0!
0%
#1665000000
1!
1%
#1670000000
0!
0%
#1675000000
1!
1%
#1680000000
0!
0%
#1685000000
1!
1%
#1690000000
0!
0%
#1695000000
1!
1%
#1700000000
0!
0%
#1705000000
1!
1%
#1710000000
0!
0%
#1715000000
1!
1%
#1720000000
0!
0%
#1725000000
1!
1%
#1730000000
0!
0%
#1735000000
1!
1%
#1740000000
0!
0%
#1745000000
1!
1%
#1750000000
0!
0%
#1755000000
1!
1%
#1760000000
0!
0%
#1765000000
1!
1%
#1770000000
0!
0%
#1775000000
1!
1%
#1780000000
0!
0%
#1785000000
1!
1%
#1790000000
0!
0%
#1795000000
1!
1%
#1800000000
0!
0%
#1805000000
1!
1%
#1810000000
0!
0%
#1815000000
1!
1%
#1820000000
0!
0%
#1825000000
1!
1%
#1830000000
0!
0%
#1835000000
1!
1%
#1840000000
0!
0%
#1845000000
1!
1%
#1850000000
0!
0%
#1855000000
1!
1%
#1860000000
0!
0%
#1865000000
1!
1%
#1870000000
0!
0%
#1875000000
1!
1%
#1880000000
0!
0%
#1885000000
1!
1%
#1890000000
0!
0%
#1895000000
1!
1%
#1900000000
0!
0%
#1905000000
1!
1%
#1910000000
0!
0%
#1915000000
1!
1%
#1920000000
0!
0%
#1925000000
1!
1%
#1930000000
0!
0%
#1935000000
1!
1%
#1940000000
0!
0%
#1945000000
1!
1%
#1950000000
0!
0%
#1955000000
1!
1%
#1960000000
0!
0%
#1965000000
1!
1%
#1970000000
0!
0%
#1975000000
1!
1%
#1980000000
0!
0%
#1985000000
1!
1%
#1990000000
0!
0%
#1995000000
1!
1%
#2000000000
0!
0%
#2005000000
1!
1%
#2010000000
0!
0%
#2015000000
1!
1%
#2020000000
0!
0%
#2025000000
1!
1%
#2030000000
0!
0%
#2035000000
1!
1%
#2040000000
0!
0%
#2045000000
1!
1%
#2050000000
0!
0%
#2055000000
1!
1%
#2060000000
0!
0%
#2065000000
1!
1%
#2070000000
0!
0%
#2075000000
1!
1%
#2080000000
0!
0%
#2085000000
1!
1%
#2090000000
0!
0%
#2095000000
1!
1%
#2100000000
0!
0%
#2105000000
1!
1%
#2110000000
0!
0%
#2115000000
1!
1%
#2120000000
0!
0%
#2125000000
1!
1%
#2130000000
0!
0%
#2135000000
1!
1%
#2140000000
0!
0%
#2145000000
1!
1%
#2150000000
0!
0%
#2155000000
1!
1%
#2160000000
0!
0%
#2165000000
1!
1%
#2170000000
0!
0%
#2175000000
1!
1%
#2180000000
0!
0%
#2185000000
1!
1%
#2190000000
0!
0%
#2195000000
1!
1%
#2200000000
0!
0%
#2205000000
1!
1%
#2210000000
0!
0%
#2215000000
1!
1%
#2220000000
0!
0%
#2225000000
1!
1%
#2230000000
0!
0%
#2235000000
1!
1%
#2240000000
0!
0%
#2245000000
1!
1%
#2250000000
0!
0%
#2255000000
1!
1%
#2260000000
0!
0%
#2265000000
1!
1%
#2270000000
0!
0%
#2275000000
1!
1%
#2280000000
0!
0%
#2285000000
1!
1%
#2290000000
0!
0%
#2295000000
1!
1%
#2300000000
0!
0%
#2305000000
1!
1%
#2310000000
0!
0%
#2315000000
1!
1%
#2320000000
0!
0%
#2325000000
1!
1%
#2330000000
0!
0%
#2335000000
1!
1%
#2340000000
0!
0%
#2345000000
1!
1%
#2350000000
0!
0%
#2355000000
1!
1%
#2360000000
0!
0%
#2365000000
1!
1%
#2370000000
0!
0%
#2375000000
1!
1%
#2380000000
0!
0%
#2385000000
1!
1%
#2390000000
0!
0%
#2395000000
1!
1%
#2400000000
0!
0%
#2405000000
1!
1%
#2410000000
0!
0%
#2415000000
1!
1%
#2420000000
0!
0%
#2425000000
1!
1%
#2430000000
0!
0%
#2435000000
1!
1%
#2440000000
0!
0%
#2445000000
1!
1%
#2450000000
0!
0%
#2455000000
1!
1%
#2460000000
0!
0%
#2465000000
1!
1%
#2470000000
0!
0%
#2475000000
1!
1%
#2480000000
0!
0%
#2485000000
1!
1%
#2490000000
0!
0%
#2495000000
1!
1%
#2500000000
0!
0%
#2505000000
1!
1%
#2510000000
0!
0%
#2515000000
1!
1%
#2520000000
0!
0%
#2525000000
1!
1%
#2530000000
0!
0%
#2535000000
1!
1%
#2540000000
0!
0%
#2545000000
1!
1%
#2550000000
0!
0%
#2555000000
1!
1%
#2560000000
0!
0%
#2565000000
1!
1%
#2570000000
0!
0%
#2575000000
1!
1%
#2580000000
0!
0%
#2585000000
1!
1%
#2590000000
0!
0%
#2595000000
1!
1%
#2600000000
0!
0%
#2605000000
1!
1%
#2610000000
0!
0%
#2615000000
1!
1%
#2620000000
0!
0%
#2625000000
1!
1%
#2630000000
0!
0%
#2635000000
1!
1%
#2640000000
0!
0%
#2645000000
1!
1%
#2650000000
0!
0%
#2655000000
1!
1%
#2660000000
0!
0%
#2665000000
1!
1%
#2670000000
0!
0%
#2675000000
1!
1%
#2680000000
0!
0%
#2685000000
1!
1%
#2690000000
0!
0%
#2695000000
1!
1%
#2700000000
0!
0%
#2705000000
1!
1%
#2710000000
0!
0%
#2715000000
1!
1%
#2720000000
0!
0%
#2725000000
1!
1%
#2730000000
0!
0%
#2735000000
1!
1%
#2740000000
0!
0%
#2745000000
1!
1%
#2750000000
0!
0%
#2755000000
1!
1%
#2760000000
0!
0%
#2765000000
1!
1%
#2770000000
0!
0%
#2775000000
1!
1%
#2780000000
0!
0%
#2785000000
1!
1%
#2790000000
0!
0%
#2795000000
1!
1%
#2800000000
0!
0%
#2805000000
1!
1%
#2810000000
0!
0%
#2815000000
1!
1%
#2820000000
0!
0%
#2825000000
1!
1%
#2830000000
0!
0%
#2835000000
1!
1%
#2840000000
0!
0%
#2845000000
1!
1%
#2850000000
0!
0%
#2855000000
1!
1%
#2860000000
0!
0%
#2865000000
1!
1%
#2870000000
0!
0%
#2875000000
1!
1%
#2880000000
0!
0%
#2885000000
1!
1%
#2890000000
0!
0%
#2895000000
1!
1%
#2900000000
0!
0%
#2905000000
1!
1%
#2910000000
0!
0%
#2915000000
1!
1%
#2920000000
0!
0%
#2925000000
1!
1%
#2930000000
0!
0%
#2935000000
1!
1%
#2940000000
0!
0%
#2945000000
1!
1%
#2950000000
0!
0%
#2955000000
1!
1%
#2960000000
0!
0%
#2965000000
1!
1%
#2970000000
0!
0%
#2975000000
1!
1%
#2980000000
0!
0%
#2985000000
1!
1%
#2990000000
0!
0%
#2995000000
1!
1%
#3000000000
0!
0%
#3005000000
1!
1%
#3010000000
0!
0%
#3015000000
1!
1%
#3020000000
0!
0%
#3025000000
1!
1%
#3030000000
0!
0%
#3035000000
1!
1%
#3040000000
0!
0%
#3045000000
1!
1%
#3050000000
0!
0%
#3055000000
1!
1%
#3060000000
0!
0%
#3065000000
1!
1%
#3070000000
0!
0%
#3075000000
1!
1%
#3080000000
0!
0%
#3085000000
1!
1%
#3090000000
0!
0%
#3095000000
1!
1%
#3100000000
0!
0%
#3105000000
1!
1%
#3110000000
0!
0%
#3115000000
1!
1%
#3120000000
0!
0%
#3125000000
1!
1%
#3130000000
0!
0%
#3135000000
1!
1%
#3140000000
0!
0%
#3145000000
1!
1%
#3150000000
0!
0%
#3155000000
1!
1%
#3160000000
0!
0%
#3165000000
1!
1%
#3170000000
0!
0%
#3175000000
1!
1%
#3180000000
0!
0%
#3185000000
1!
1%
#3190000000
0!
0%
#3195000000
1!
1%
#3200000000
0!
0%
#3205000000
1!
1%
#3210000000
0!
0%
#3215000000
1!
1%
#3220000000
0!
0%
#3225000000
1!
1%
#3230000000
0!
0%
#3235000000
1!
1%
#3240000000
0!
0%
#3245000000
1!
1%
#3250000000
0!
0%
#3255000000
1!
1%
#3260000000
0!
0%
#3265000000
1!
1%
#3270000000
0!
0%
#3275000000
1!
1%
#3280000000
0!
0%
#3285000000
1!
1%
#3290000000
0!
0%
#3295000000
1!
1%
#3300000000
0!
0%
#3305000000
1!
1%
#3310000000
0!
0%
#3315000000
1!
1%
#3320000000
0!
0%
#3325000000
1!
1%
#3330000000
0!
0%
#3335000000
1!
1%
#3340000000
0!
0%
#3345000000
1!
1%
#3350000000
0!
0%
#3355000000
1!
1%
#3360000000
0!
0%
#3365000000
1!
1%
#3370000000
0!
0%
#3375000000
1!
1%
#3380000000
0!
0%
#3385000000
1!
1%
#3390000000
0!
0%
#3395000000
1!
1%
#3400000000
0!
0%
#3405000000
1!
1%
#3410000000
0!
0%
#3415000000
1!
1%
#3420000000
0!
0%
#3425000000
1!
1%
#3430000000
0!
0%
#3435000000
1!
1%
#3440000000
0!
0%
#3445000000
1!
1%
#3450000000
0!
0%
#3455000000
1!
1%
#3460000000
0!
0%
#3465000000
1!
1%
#3470000000
0!
0%
#3475000000
1!
1%
#3480000000
0!
0%
#3485000000
1!
1%
#3490000000
0!
0%
#3495000000
1!
1%
#3500000000
0!
0%
#3505000000
1!
1%
#3510000000
0!
0%
#3515000000
1!
1%
#3520000000
0!
0%
#3525000000
1!
1%
#3530000000
0!
0%
#3535000000
1!
1%
#3540000000
0!
0%
#3545000000
1!
1%
#3550000000
0!
0%
#3555000000
1!
1%
#3560000000
0!
0%
#3565000000
1!
1%
#3570000000
0!
0%
#3575000000
1!
1%
#3580000000
0!
0%
#3585000000
1!
1%
#3590000000
0!
0%
#3595000000
1!
1%
#3600000000
0!
0%
#3605000000
1!
1%
#3610000000
0!
0%
#3615000000
1!
1%
#3620000000
0!
0%
#3625000000
1!
1%
#3630000000
0!
0%
#3635000000
1!
1%
#3640000000
0!
0%
#3645000000
1!
1%
#3650000000
0!
0%
#3655000000
1!
1%
#3660000000
0!
0%
#3665000000
1!
1%
#3670000000
0!
0%
#3675000000
1!
1%
#3680000000
0!
0%
#3685000000
1!
1%
#3690000000
0!
0%
#3695000000
1!
1%
#3700000000
0!
0%
#3705000000
1!
1%
#3710000000
0!
0%
#3715000000
1!
1%
#3720000000
0!
0%
#3725000000
1!
1%
#3730000000
0!
0%
#3735000000
1!
1%
#3740000000
0!
0%
#3745000000
1!
1%
#3750000000
0!
0%
#3755000000
1!
1%
#3760000000
0!
0%
#3765000000
1!
1%
#3770000000
0!
0%
#3775000000
1!
1%
#3780000000
0!
0%
#3785000000
1!
1%
#3790000000
0!
0%
#3795000000
1!
1%
#3800000000
0!
0%
#3805000000
1!
1%
#3810000000
0!
0%
#3815000000
1!
1%
#3820000000
0!
0%
#3825000000
1!
1%
#3830000000
0!
0%
#3835000000
1!
1%
#3840000000
0!
0%
#3845000000
1!
1%
#3850000000
0!
0%
#3855000000
1!
1%
#3860000000
0!
0%
#3865000000
1!
1%
#3870000000
0!
0%
#3875000000
1!
1%
#3880000000
0!
0%
#3885000000
1!
1%
#3890000000
0!
0%
#3895000000
1!
1%
#3900000000
0!
0%
#3905000000
1!
1%
#3910000000
0!
0%
#3915000000
1!
1%
#3920000000
0!
0%
#3925000000
1!
1%
#3930000000
0!
0%
#3935000000
1!
1%
#3940000000
0!
0%
#3945000000
1!
1%
#3950000000
0!
0%
#3955000000
1!
1%
#3960000000
0!
0%
#3965000000
1!
1%
#3970000000
0!
0%
#3975000000
1!
1%
#3980000000
0!
0%
#3985000000
1!
1%
#3990000000
0!
0%
#3995000000
1!
1%
#4000000000
0!
0%
#4005000000
1!
1%
#4010000000
0!
0%
#4015000000
1!
1%
#4020000000
0!
0%
#4025000000
1!
1%
#4030000000
0!
0%
#4035000000
1!
1%
#4040000000
0!
0%
#4045000000
1!
1%
#4050000000
0!
0%
#4055000000
1!
1%
#4060000000
0!
0%
#4065000000
1!
1%
#4070000000
0!
0%
#4075000000
1!
1%
#4080000000
0!
0%
#4085000000
1!
1%
#4090000000
0!
0%
#4095000000
1!
1%
#4100000000
0!
0%
#4105000000
1!
1%
#4110000000
0!
0%
#4115000000
1!
1%
#4120000000
0!
0%
#4125000000
1!
1%
#4130000000
0!
0%
#4135000000
1!
1%
#4140000000
0!
0%
#4145000000
1!
1%
#4150000000
0!
0%
#4155000000
1!
1%
#4160000000
0!
0%
#4165000000
1!
1%
#4170000000
0!
0%
#4175000000
1!
1%
#4180000000
0!
0%
#4185000000
1!
1%
#4190000000
0!
0%
#4195000000
1!
1%
#4200000000
0!
0%
#4205000000
1!
1%
#4210000000
0!
0%
#4215000000
1!
1%
#4220000000
0!
0%
#4225000000
1!
1%
#4230000000
0!
0%
#4235000000
1!
1%
#4240000000
0!
0%
#4245000000
1!
1%
#4250000000
0!
0%
#4255000000
1!
1%
#4260000000
0!
0%
#4265000000
1!
1%
#4270000000
0!
0%
#4275000000
1!
1%
#4280000000
0!
0%
#4285000000
1!
1%
#4290000000
0!
0%
#4295000000
1!
1%
#4300000000
0!
0%
#4305000000
1!
1%
#4310000000
0!
0%
#4315000000
1!
1%
#4320000000
0!
0%
#4325000000
1!
1%
#4330000000
0!
0%
#4335000000
1!
1%
#4340000000
0!
0%
#4345000000
1!
1%
#4350000000
0!
0%
#4355000000
1!
1%
#4360000000
0!
0%
#4365000000
1!
1%
#4370000000
0!
0%
#4375000000
1!
1%
#4380000000
0!
0%
#4385000000
1!
1%
#4390000000
0!
0%
#4395000000
1!
1%
#4400000000
0!
0%
#4405000000
1!
1%
#4410000000
0!
0%
#4415000000
1!
1%
#4420000000
0!
0%
#4425000000
1!
1%
#4430000000
0!
0%
#4435000000
1!
1%
#4440000000
0!
0%
#4445000000
1!
1%
#4450000000
0!
0%
#4455000000
1!
1%
#4460000000
0!
0%
#4465000000
1!
1%
#4470000000
0!
0%
#4475000000
1!
1%
#4480000000
0!
0%
#4485000000
1!
1%
#4490000000
0!
0%
#4495000000
1!
1%
#4500000000
0!
0%
#4505000000
1!
1%
#4510000000
0!
0%
#4515000000
1!
1%
#4520000000
0!
0%
#4525000000
1!
1%
#4530000000
0!
0%
#4535000000
1!
1%
#4540000000
0!
0%
#4545000000
1!
1%
#4550000000
0!
0%
#4555000000
1!
1%
#4560000000
0!
0%
#4565000000
1!
1%
#4570000000
0!
0%
#4575000000
1!
1%
#4580000000
0!
0%
#4585000000
1!
1%
#4590000000
0!
0%
#4595000000
1!
1%
#4600000000
0!
0%
#4605000000
1!
1%
#4610000000
0!
0%
#4615000000
1!
1%
#4620000000
0!
0%
#4625000000
1!
1%
#4630000000
0!
0%
#4635000000
1!
1%
#4640000000
0!
0%
#4645000000
1!
1%
#4650000000
0!
0%
#4655000000
1!
1%
#4660000000
0!
0%
#4665000000
1!
1%
#4670000000
0!
0%
#4675000000
1!
1%
#4680000000
0!
0%
#4685000000
1!
1%
#4690000000
0!
0%
#4695000000
1!
1%
#4700000000
0!
0%
#4705000000
1!
1%
#4710000000
0!
0%
#4715000000
1!
1%
#4720000000
0!
0%
#4725000000
1!
1%
#4730000000
0!
0%
#4735000000
1!
1%
#4740000000
0!
0%
#4745000000
1!
1%
#4750000000
0!
0%
#4755000000
1!
1%
#4760000000
0!
0%
#4765000000
1!
1%
#4770000000
0!
0%
#4775000000
1!
1%
#4780000000
0!
0%
#4785000000
1!
1%
#4790000000
0!
0%
#4795000000
1!
1%
#4800000000
0!
0%
#4805000000
1!
1%
#4810000000
0!
0%
#4815000000
1!
1%
#4820000000
0!
0%
#4825000000
1!
1%
#4830000000
0!
0%
#4835000000
1!
1%
#4840000000
0!
0%
#4845000000
1!
1%
#4850000000
0!
0%
#4855000000
1!
1%
#4860000000
0!
0%
#4865000000
1!
1%
#4870000000
0!
0%
#4875000000
1!
1%
#4880000000
0!
0%
#4885000000
1!
1%
#4890000000
0!
0%
#4895000000
1!
1%
#4900000000
0!
0%
#4905000000
1!
1%
#4910000000
0!
0%
#4915000000
1!
1%
#4920000000
0!
0%
#4925000000
1!
1%
#4930000000
0!
0%
#4935000000
1!
1%
#4940000000
0!
0%
#4945000000
1!
1%
#4950000000
0!
0%
#4955000000
1!
1%
#4960000000
0!
0%
#4965000000
1!
1%
#4970000000
0!
0%
#4975000000
1!
1%
#4980000000
0!
0%
#4985000000
1!
1%
#4990000000
0!
0%
#4995000000
1!
1%
#5000000000
0!
0%
#5005000000
1!
1%
#5010000000
0!
0%
#5015000000
1!
1%
#5020000000
0!
0%
#5025000000
1!
1%
#5030000000
0!
0%
#5035000000
1!
1%
#5040000000
0!
0%
#5045000000
1!
1%
#5050000000
0!
0%
#5055000000
1!
1%
#5060000000
0!
0%
#5065000000
1!
1%
#5070000000
0!
0%
#5075000000
1!
1%
#5080000000
0!
0%
#5085000000
1!
1%
#5090000000
0!
0%
#5095000000
1!
1%
#5100000000
0!
0%
#5105000000
1!
1%
#5110000000
0!
0%
#5115000000
1!
1%
#5120000000
0!
0%
#5125000000
1!
1%
#5130000000
0!
0%
#5135000000
1!
1%
#5140000000
0!
0%
#5145000000
1!
1%
#5150000000
0!
0%
#5155000000
1!
1%
#5160000000
0!
0%
#5165000000
1!
1%
#5170000000
0!
0%
#5175000000
1!
1%
#5180000000
0!
0%
#5185000000
1!
1%
#5190000000
0!
0%
#5195000000
1!
1%
#5200000000
0!
0%
#5205000000
1!
1%
#5210000000
0!
0%
#5215000000
1!
1%
#5220000000
0!
0%
#5225000000
1!
1%
#5230000000
0!
0%
#5235000000
1!
1%
#5240000000
0!
0%
#5245000000
1!
1%
#5250000000
0!
0%
#5255000000
1!
1%
#5260000000
0!
0%
#5265000000
1!
1%
#5270000000
0!
0%
#5275000000
1!
1%
#5280000000
0!
0%
#5285000000
1!
1%
#5290000000
0!
0%
#5295000000
1!
1%
#5300000000
0!
0%
#5305000000
1!
1%
#5310000000
0!
0%
#5315000000
1!
1%
#5320000000
0!
0%
#5325000000
1!
1%
#5330000000
0!
0%
#5335000000
1!
1%
#5340000000
0!
0%
#5345000000
1!
1%
#5350000000
0!
0%
#5355000000
1!
1%
#5360000000
0!
0%
#5365000000
1!
1%
#5370000000
0!
0%
#5375000000
1!
1%
#5380000000
0!
0%
#5385000000
1!
1%
#5390000000
0!
0%
#5395000000
1!
1%
#5400000000
0!
0%
#5405000000
1!
1%
#5410000000
0!
0%
#5415000000
1!
1%
#5420000000
0!
0%
#5425000000
1!
1%
#5430000000
0!
0%
#5435000000
1!
1%
#5440000000
0!
0%
#5445000000
1!
1%
#5450000000
0!
0%
#5455000000
1!
1%
#5460000000
0!
0%
#5465000000
1!
1%
#5470000000
0!
0%
#5475000000
1!
1%
#5480000000
0!
0%
#5485000000
1!
1%
#5490000000
0!
0%
#5495000000
1!
1%
#5500000000
0!
0%
#5505000000
1!
1%
#5510000000
0!
0%
#5515000000
1!
1%
#5520000000
0!
0%
#5525000000
1!
1%
#5530000000
0!
0%
#5535000000
1!
1%
#5540000000
0!
0%
#5545000000
1!
1%
#5550000000
0!
0%
#5555000000
1!
1%
#5560000000
0!
0%
#5565000000
1!
1%
#5570000000
0!
0%
#5575000000
1!
1%
#5580000000
0!
0%
#5585000000
1!
1%
#5590000000
0!
0%
#5595000000
1!
1%
#5600000000
0!
0%
#5605000000
1!
1%
#5610000000
0!
0%
#5615000000
1!
1%
#5620000000
0!
0%
#5625000000
1!
1%
#5630000000
0!
0%
#5635000000
1!
1%
#5640000000
0!
0%
#5645000000
1!
1%
#5650000000
0!
0%
#5655000000
1!
1%
#5660000000
0!
0%
#5665000000
1!
1%
#5670000000
0!
0%
#5675000000
1!
1%
#5680000000
0!
0%
#5685000000
1!
1%
#5690000000
0!
0%
#5695000000
1!
1%
#5700000000
0!
0%
#5705000000
1!
1%
#5710000000
0!
0%
#5715000000
1!
1%
#5720000000
0!
0%
#5725000000
1!
1%
#5730000000
0!
0%
#5735000000
1!
1%
#5740000000
0!
0%
#5745000000
1!
1%
#5750000000
0!
0%
#5755000000
1!
1%
#5760000000
0!
0%
#5765000000
1!
1%
#5770000000
0!
0%
#5775000000
1!
1%
#5780000000
0!
0%
#5785000000
1!
1%
#5790000000
0!
0%
#5795000000
1!
1%
#5800000000
0!
0%
#5805000000
1!
1%
#5810000000
0!
0%
#5815000000
1!
1%
#5820000000
0!
0%
#5825000000
1!
1%
#5830000000
0!
0%
#5835000000
1!
1%
#5840000000
0!
0%
#5845000000
1!
1%
#5850000000
0!
0%
#5855000000
1!
1%
#5860000000
0!
0%
#5865000000
1!
1%
#5870000000
0!
0%
#5875000000
1!
1%
#5880000000
0!
0%
#5885000000
1!
1%
#5890000000
0!
0%
#5895000000
1!
1%
#5900000000
0!
0%
#5905000000
1!
1%
#5910000000
0!
0%
#5915000000
1!
1%
#5920000000
0!
0%
#5925000000
1!
1%
#5930000000
0!
0%
#5935000000
1!
1%
#5940000000
0!
0%
#5945000000
1!
1%
#5950000000
0!
0%
#5955000000
1!
1%
#5960000000
0!
0%
#5965000000
1!
1%
#5970000000
0!
0%
#5975000000
1!
1%
#5980000000
0!
0%
#5985000000
1!
1%
#5990000000
0!
0%
#5995000000
1!
1%
#6000000000
0!
0%
#6005000000
1!
1%
#6010000000
0!
0%
#6015000000
1!
1%
#6020000000
0!
0%
#6025000000
1!
1%
#6030000000
0!
0%
#6035000000
1!
1%
#6040000000
0!
0%
#6045000000
1!
1%
#6050000000
0!
0%
#6055000000
1!
1%
#6060000000
0!
0%
#6065000000
1!
1%
#6070000000
0!
0%
#6075000000
1!
1%
#6080000000
0!
0%
#6085000000
1!
1%
#6090000000
0!
0%
#6095000000
1!
1%
#6100000000
0!
0%
#6105000000
1!
1%
#6110000000
0!
0%
#6115000000
1!
1%
#6120000000
0!
0%
#6125000000
1!
1%
#6130000000
0!
0%
#6135000000
1!
1%
#6140000000
0!
0%
#6145000000
1!
1%
#6150000000
0!
0%
#6155000000
1!
1%
#6160000000
0!
0%
#6165000000
1!
1%
#6170000000
0!
0%
#6175000000
1!
1%
#6180000000
0!
0%
#6185000000
1!
1%
#6190000000
0!
0%
#6195000000
1!
1%
#6200000000
0!
0%
#6205000000
1!
1%
#6210000000
0!
0%
#6215000000
1!
1%
#6220000000
0!
0%
#6225000000
1!
1%
#6230000000
0!
0%
#6235000000
1!
1%
#6240000000
0!
0%
#6245000000
1!
1%
#6250000000
0!
0%
#6255000000
1!
1%
#6260000000
0!
0%
#6265000000
1!
1%
#6270000000
0!
0%
#6275000000
1!
1%
#6280000000
0!
0%
#6285000000
1!
1%
#6290000000
0!
0%
#6295000000
1!
1%
#6300000000
0!
0%
#6305000000
1!
1%
#6310000000
0!
0%
#6315000000
1!
1%
#6320000000
0!
0%
#6325000000
1!
1%
#6330000000
0!
0%
#6335000000
1!
1%
#6340000000
0!
0%
#6345000000
1!
1%
#6350000000
0!
0%
#6355000000
1!
1%
#6360000000
0!
0%
#6365000000
1!
1%
#6370000000
0!
0%
#6375000000
1!
1%
#6380000000
0!
0%
#6385000000
1!
1%
#6390000000
0!
0%
#6395000000
1!
1%
#6400000000
0!
0%
#6405000000
1!
1%
#6410000000
0!
0%
#6415000000
1!
1%
#6420000000
0!
0%
#6425000000
1!
1%
#6430000000
0!
0%
#6435000000
1!
1%
#6440000000
0!
0%
#6445000000
1!
1%
#6450000000
0!
0%
#6455000000
1!
1%
#6460000000
0!
0%
#6465000000
1!
1%
#6470000000
0!
0%
#6475000000
1!
1%
#6480000000
0!
0%
#6485000000
1!
1%
#6490000000
0!
0%
#6495000000
1!
1%
#6500000000
0!
0%
#6505000000
1!
1%
#6510000000
0!
0%
#6515000000
1!
1%
#6520000000
0!
0%
#6525000000
1!
1%
#6530000000
0!
0%
#6535000000
1!
1%
#6540000000
0!
0%
#6545000000
1!
1%
#6550000000
0!
0%
#6555000000
1!
1%
#6560000000
0!
0%
#6565000000
1!
1%
#6570000000
0!
0%
#6575000000
1!
1%
#6580000000
0!
0%
#6585000000
1!
1%
#6590000000
0!
0%
#6595000000
1!
1%
#6600000000
0!
0%
#6605000000
1!
1%
#6610000000
0!
0%
#6615000000
1!
1%
#6620000000
0!
0%
#6625000000
1!
1%
#6630000000
0!
0%
#6635000000
1!
1%
#6640000000
0!
0%
#6645000000
1!
1%
#6650000000
0!
0%
#6655000000
1!
1%
#6660000000
0!
0%
#6665000000
1!
1%
#6670000000
0!
0%
#6675000000
1!
1%
#6680000000
0!
0%
#6685000000
1!
1%
#6690000000
0!
0%
#6695000000
1!
1%
#6700000000
0!
0%
#6705000000
1!
1%
#6710000000
0!
0%
#6715000000
1!
1%
#6720000000
0!
0%
#6725000000
1!
1%
#6730000000
0!
0%
#6735000000
1!
1%
#6740000000
0!
0%
#6745000000
1!
1%
#6750000000
0!
0%
#6755000000
1!
1%
#6760000000
0!
0%
#6765000000
1!
1%
#6770000000
0!
0%
#6775000000
1!
1%
#6780000000
0!
0%
#6785000000
1!
1%
#6790000000
0!
0%
#6795000000
1!
1%
#6800000000
0!
0%
#6805000000
1!
1%
#6810000000
0!
0%
#6815000000
1!
1%
#6820000000
0!
0%
#6825000000
1!
1%
#6830000000
0!
0%
#6835000000
1!
1%
#6840000000
0!
0%
#6845000000
1!
1%
#6850000000
0!
0%
#6855000000
1!
1%
#6860000000
0!
0%
#6865000000
1!
1%
#6870000000
0!
0%
#6875000000
1!
1%
#6880000000
0!
0%
#6885000000
1!
1%
#6890000000
0!
0%
#6895000000
1!
1%
#6900000000
0!
0%
#6905000000
1!
1%
#6910000000
0!
0%
#6915000000
1!
1%
#6920000000
0!
0%
#6925000000
1!
1%
#6930000000
0!
0%
#6935000000
1!
1%
#6940000000
0!
0%
#6945000000
1!
1%
#6950000000
0!
0%
#6955000000
1!
1%
#6960000000
0!
0%
#6965000000
1!
1%
#6970000000
0!
0%
#6975000000
1!
1%
#6980000000
0!
0%
#6985000000
1!
1%
#6990000000
0!
0%
#6995000000
1!
1%
#7000000000
0!
0%
#7005000000
1!
1%
#7010000000
0!
0%
#7015000000
1!
1%
#7020000000
0!
0%
#7025000000
1!
1%
#7030000000
0!
0%
#7035000000
1!
1%
#7040000000
0!
0%
#7045000000
1!
1%
#7050000000
0!
0%
#7055000000
1!
1%
#7060000000
0!
0%
#7065000000
1!
1%
#7070000000
0!
0%
#7075000000
1!
1%
#7080000000
0!
0%
#7085000000
1!
1%
#7090000000
0!
0%
#7095000000
1!
1%
#7100000000
0!
0%
#7105000000
1!
1%
#7110000000
0!
0%
#7115000000
1!
1%
#7120000000
0!
0%
#7125000000
1!
1%
#7130000000
0!
0%
#7135000000
1!
1%
#7140000000
0!
0%
#7145000000
1!
1%
#7150000000
0!
0%
#7155000000
1!
1%
#7160000000
0!
0%
#7165000000
1!
1%
#7170000000
0!
0%
#7175000000
1!
1%
#7180000000
0!
0%
#7185000000
1!
1%
#7190000000
0!
0%
#7195000000
1!
1%
#7200000000
0!
0%
#7205000000
1!
1%
#7210000000
0!
0%
#7215000000
1!
1%
#7220000000
0!
0%
#7225000000
1!
1%
#7230000000
0!
0%
#7235000000
1!
1%
#7240000000
0!
0%
#7245000000
1!
1%
#7250000000
0!
0%
#7255000000
1!
1%
#7260000000
0!
0%
#7265000000
1!
1%
#7270000000
0!
0%
#7275000000
1!
1%
#7280000000
0!
0%
#7285000000
1!
1%
#7290000000
0!
0%
#7295000000
1!
1%
#7300000000
0!
0%
#7305000000
1!
1%
#7310000000
0!
0%
#7315000000
1!
1%
#7320000000
0!
0%
#7325000000
1!
1%
#7330000000
0!
0%
#7335000000
1!
1%
#7340000000
0!
0%
#7345000000
1!
1%
#7350000000
0!
0%
#7355000000
1!
1%
#7360000000
0!
0%
#7365000000
1!
1%
#7370000000
0!
0%
#7375000000
1!
1%
#7380000000
0!
0%
#7385000000
1!
1%
#7390000000
0!
0%
#7395000000
1!
1%
#7400000000
0!
0%
#7405000000
1!
1%
#7410000000
0!
0%
#7415000000
1!
1%
#7420000000
0!
0%
#7425000000
1!
1%
#7430000000
0!
0%
#7435000000
1!
1%
#7440000000
0!
0%
#7445000000
1!
1%
#7450000000
0!
0%
#7455000000
1!
1%
#7460000000
0!
0%
#7465000000
1!
1%
#7470000000
0!
0%
#7475000000
1!
1%
#7480000000
0!
0%
#7485000000
1!
1%
#7490000000
0!
0%
#7495000000
1!
1%
#7500000000
0!
0%
#7505000000
1!
1%
#7510000000
0!
0%
#7515000000
1!
1%
#7520000000
0!
0%
#7525000000
1!
1%
#7530000000
0!
0%
#7535000000
1!
1%
#7540000000
0!
0%
#7545000000
1!
1%
#7550000000
0!
0%
#7555000000
1!
1%
#7560000000
0!
0%
#7565000000
1!
1%
#7570000000
0!
0%
#7575000000
1!
1%
#7580000000
0!
0%
#7585000000
1!
1%
#7590000000
0!
0%
#7595000000
1!
1%
#7600000000
0!
0%
#7605000000
1!
1%
#7610000000
0!
0%
#7615000000
1!
1%
#7620000000
0!
0%
#7625000000
1!
1%
#7630000000
0!
0%
#7635000000
1!
1%
#7640000000
0!
0%
#7645000000
1!
1%
#7650000000
0!
0%
#7655000000
1!
1%
#7660000000
0!
0%
#7665000000
1!
1%
#7670000000
0!
0%
#7675000000
1!
1%
#7680000000
0!
0%
#7685000000
1!
1%
#7690000000
0!
0%
#7695000000
1!
1%
#7700000000
0!
0%
#7705000000
1!
1%
#7710000000
0!
0%
#7715000000
1!
1%
#7720000000
0!
0%
#7725000000
1!
1%
#7730000000
0!
0%
#7735000000
1!
1%
#7740000000
0!
0%
#7745000000
1!
1%
#7750000000
0!
0%
#7755000000
1!
1%
#7760000000
0!
0%
#7765000000
1!
1%
#7770000000
0!
0%
#7775000000
1!
1%
#7780000000
0!
0%
#7785000000
1!
1%
#7790000000
0!
0%
#7795000000
1!
1%
#7800000000
0!
0%
#7805000000
1!
1%
#7810000000
0!
0%
#7815000000
1!
1%
#7820000000
0!
0%
#7825000000
1!
1%
#7830000000
0!
0%
#7835000000
1!
1%
#7840000000
0!
0%
#7845000000
1!
1%
#7850000000
0!
0%
#7855000000
1!
1%
#7860000000
0!
0%
#7865000000
1!
1%
#7870000000
0!
0%
#7875000000
1!
1%
#7880000000
0!
0%
#7885000000
1!
1%
#7890000000
0!
0%
#7895000000
1!
1%
#7900000000
0!
0%
#7905000000
1!
1%
#7910000000
0!
0%
#7915000000
1!
1%
#7920000000
0!
0%
#7925000000
1!
1%
#7930000000
0!
0%
#7935000000
1!
1%
#7940000000
0!
0%
#7945000000
1!
1%
#7950000000
0!
0%
#7955000000
1!
1%
#7960000000
0!
0%
#7965000000
1!
1%
#7970000000
0!
0%
#7975000000
1!
1%
#7980000000
0!
0%
#7985000000
1!
1%
#7990000000
0!
0%
#7995000000
1!
1%
#8000000000
0!
0%
#8005000000
1!
1%
#8010000000
0!
0%
#8015000000
1!
1%
#8020000000
0!
0%
#8025000000
1!
1%
#8030000000
0!
0%
#8035000000
1!
1%
#8040000000
0!
0%
#8045000000
1!
1%
#8050000000
0!
0%
#8055000000
1!
1%
#8060000000
0!
0%
#8065000000
1!
1%
#8070000000
0!
0%
#8075000000
1!
1%
#8080000000
0!
0%
#8085000000
1!
1%
#8090000000
0!
0%
#8095000000
1!
1%
#8100000000
0!
0%
#8105000000
1!
1%
#8110000000
0!
0%
#8115000000
1!
1%
#8120000000
0!
0%
#8125000000
1!
1%
#8130000000
0!
0%
#8135000000
1!
1%
#8140000000
0!
0%
#8145000000
1!
1%
#8150000000
0!
0%
#8155000000
1!
1%
#8160000000
0!
0%
#8165000000
1!
1%
#8170000000
0!
0%
#8175000000
1!
1%
#8180000000
0!
0%
#8185000000
1!
1%
#8190000000
0!
0%
#8195000000
1!
1%
#8200000000
0!
0%
#8205000000
1!
1%
#8210000000
0!
0%
#8215000000
1!
1%
#8220000000
0!
0%
#8225000000
1!
1%
#8230000000
0!
0%
#8235000000
1!
1%
#8240000000
0!
0%
#8245000000
1!
1%
#8250000000
0!
0%
#8255000000
1!
1%
#8260000000
0!
0%
#8265000000
1!
1%
#8270000000
0!
0%
#8275000000
1!
1%
#8280000000
0!
0%
#8285000000
1!
1%
#8290000000
0!
0%
#8295000000
1!
1%
#8300000000
0!
0%
#8305000000
1!
1%
#8310000000
0!
0%
#8315000000
1!
1%
#8320000000
0!
0%
#8325000000
1!
1%
#8330000000
0!
0%
#8335000000
1!
1%
#8340000000
0!
0%
#8345000000
1!
1%
#8350000000
0!
0%
#8355000000
1!
1%
#8360000000
0!
0%
#8365000000
1!
1%
#8370000000
0!
0%
#8375000000
1!
1%
#8380000000
0!
0%
#8385000000
1!
1%
#8390000000
0!
0%
#8395000000
1!
1%
#8400000000
0!
0%
#8405000000
1!
1%
#8410000000
0!
0%
#8415000000
1!
1%
#8420000000
0!
0%
#8425000000
1!
1%
#8430000000
0!
0%
#8435000000
1!
1%
#8440000000
0!
0%
#8445000000
1!
1%
#8450000000
0!
0%
#8455000000
1!
1%
#8460000000
0!
0%
#8465000000
1!
1%
#8470000000
0!
0%
#8475000000
1!
1%
#8480000000
0!
0%
#8485000000
1!
1%
#8490000000
0!
0%
#8495000000
1!
1%
#8500000000
0!
0%
#8505000000
1!
1%
#8510000000
0!
0%
#8515000000
1!
1%
#8520000000
0!
0%
#8525000000
1!
1%
#8530000000
0!
0%
#8535000000
1!
1%
#8540000000
0!
0%
#8545000000
1!
1%
#8550000000
0!
0%
#8555000000
1!
1%
#8560000000
0!
0%
#8565000000
1!
1%
#8570000000
0!
0%
#8575000000
1!
1%
#8580000000
0!
0%
#8585000000
1!
1%
#8590000000
0!
0%
#8595000000
1!
1%
#8600000000
0!
0%
#8605000000
1!
1%
#8610000000
0!
0%
#8615000000
1!
1%
#8620000000
0!
0%
#8625000000
1!
1%
#8630000000
0!
0%
#8635000000
1!
1%
#8640000000
0!
0%
#8645000000
1!
1%
#8650000000
0!
0%
#8655000000
1!
1%
#8660000000
0!
0%
#8665000000
1!
1%
#8670000000
0!
0%
#8675000000
1!
1%
#8680000000
0!
0%
#8685000000
1!
1%
#8690000000
0!
0%
#8695000000
1!
1%
#8700000000
0!
0%
#8705000000
1!
1%
#8710000000
0!
0%
#8715000000
1!
1%
#8720000000
0!
0%
#8725000000
1!
1%
#8730000000
0!
0%
#8735000000
1!
1%
#8740000000
0!
0%
#8745000000
1!
1%
#8750000000
0!
0%
#8755000000
1!
1%
#8760000000
0!
0%
#8765000000
1!
1%
#8770000000
0!
0%
#8775000000
1!
1%
#8780000000
0!
0%
#8785000000
1!
1%
#8790000000
0!
0%
#8795000000
1!
1%
#8800000000
0!
0%
#8805000000
1!
1%
#8810000000
0!
0%
#8815000000
1!
1%
#8820000000
0!
0%
#8825000000
1!
1%
#8830000000
0!
0%
#8835000000
1!
1%
#8840000000
0!
0%
#8845000000
1!
1%
#8850000000
0!
0%
#8855000000
1!
1%
#8860000000
0!
0%
#8865000000
1!
1%
#8870000000
0!
0%
#8875000000
1!
1%
#8880000000
0!
0%
#8885000000
1!
1%
#8890000000
0!
0%
#8895000000
1!
1%
#8900000000
0!
0%
#8905000000
1!
1%
#8910000000
0!
0%
#8915000000
1!
1%
#8920000000
0!
0%
#8925000000
1!
1%
#8930000000
0!
0%
#8935000000
1!
1%
#8940000000
0!
0%
#8945000000
1!
1%
#8950000000
0!
0%
#8955000000
1!
1%
#8960000000
0!
0%
#8965000000
1!
1%
#8970000000
0!
0%
#8975000000
1!
1%
#8980000000
0!
0%
#8985000000
1!
1%
#8990000000
0!
0%
#8995000000
1!
1%
#9000000000
0!
0%
#9005000000
1!
1%
#9010000000
0!
0%
#9015000000
1!
1%
#9020000000
0!
0%
#9025000000
1!
1%
#9030000000
0!
0%
#9035000000
1!
1%
#9040000000
0!
0%
#9045000000
1!
1%
#9050000000
0!
0%
#9055000000
1!
1%
#9060000000
0!
0%
#9065000000
1!
1%
#9070000000
0!
0%
#9075000000
1!
1%
#9080000000
0!
0%
#9085000000
1!
1%
#9090000000
0!
0%
#9095000000
1!
1%
#9100000000
0!
0%
#9105000000
1!
1%
#9110000000
0!
0%
#9115000000
1!
1%
#9120000000
0!
0%
#9125000000
1!
1%
#9130000000
0!
0%
#9135000000
1!
1%
#9140000000
0!
0%
#9145000000
1!
1%
#9150000000
0!
0%
#9155000000
1!
1%
#9160000000
0!
0%
#9165000000
1!
1%
#9170000000
0!
0%
#9175000000
1!
1%
#9180000000
0!
0%
#9185000000
1!
1%
#9190000000
0!
0%
#9195000000
1!
1%
#9200000000
0!
0%
#9205000000
1!
1%
#9210000000
0!
0%
#9215000000
1!
1%
#9220000000
0!
0%
#9225000000
1!
1%
#9230000000
0!
0%
#9235000000
1!
1%
#9240000000
0!
0%
#9245000000
1!
1%
#9250000000
0!
0%
#9255000000
1!
1%
#9260000000
0!
0%
#9265000000
1!
1%
#9270000000
0!
0%
#9275000000
1!
1%
#9280000000
0!
0%
#9285000000
1!
1%
#9290000000
0!
0%
#9295000000
1!
1%
#9300000000
0!
0%
#9305000000
1!
1%
#9310000000
0!
0%
#9315000000
1!
1%
#9320000000
0!
0%
#9325000000
1!
1%
#9330000000
0!
0%
#9335000000
1!
1%
#9340000000
0!
0%
#9345000000
1!
1%
#9350000000
0!
0%
#9355000000
1!
1%
#9360000000
0!
0%
#9365000000
1!
1%
#9370000000
0!
0%
#9375000000
1!
1%
#9380000000
0!
0%
#9385000000
1!
1%
#9390000000
0!
0%
#9395000000
1!
1%
#9400000000
0!
0%
#9405000000
1!
1%
#9410000000
0!
0%
#9415000000
1!
1%
#9420000000
0!
0%
#9425000000
1!
1%
#9430000000
0!
0%
#9435000000
1!
1%
#9440000000
0!
0%
#9445000000
1!
1%
#9450000000
0!
0%
#9455000000
1!
1%
#9460000000
0!
0%
#9465000000
1!
1%
#9470000000
0!
0%
#9475000000
1!
1%
#9480000000
0!
0%
#9485000000
1!
1%
#9490000000
0!
0%
#9495000000
1!
1%
#9500000000
0!
0%
#9505000000
1!
1%
#9510000000
0!
0%
#9515000000
1!
1%
#9520000000
0!
0%
#9525000000
1!
1%
#9530000000
0!
0%
#9535000000
1!
1%
#9540000000
0!
0%
#9545000000
1!
1%
#9550000000
0!
0%
#9555000000
1!
1%
#9560000000
0!
0%
#9565000000
1!
1%
#9570000000
0!
0%
#9575000000
1!
1%
#9580000000
0!
0%
#9585000000
1!
1%
#9590000000
0!
0%
#9595000000
1!
1%
#9600000000
0!
0%
#9605000000
1!
1%
#9610000000
0!
0%
#9615000000
1!
1%
#9620000000
0!
0%
#9625000000
1!
1%
#9630000000
0!
0%
#9635000000
1!
1%
#9640000000
0!
0%
#9645000000
1!
1%
#9650000000
0!
0%
#9655000000
1!
1%
#9660000000
0!
0%
#9665000000
1!
1%
#9670000000
0!
0%
#9675000000
1!
1%
#9680000000
0!
0%
#9685000000
1!
1%
#9690000000
0!
0%
#9695000000
1!
1%
#9700000000
0!
0%
#9705000000
1!
1%
#9710000000
0!
0%
#9715000000
1!
1%
#9720000000
0!
0%
#9725000000
1!
1%
#9730000000
0!
0%
#9735000000
1!
1%
#9740000000
0!
0%
#9745000000
1!
1%
#9750000000
0!
0%
#9755000000
1!
1%
#9760000000
0!
0%
#9765000000
1!
1%
#9770000000
0!
0%
#9775000000
1!
1%
#9780000000
0!
0%
#9785000000
1!
1%
#9790000000
0!
0%
#9795000000
1!
1%
#9800000000
0!
0%
#9805000000
1!
1%
#9810000000
0!
0%
#9815000000
1!
1%
#9820000000
0!
0%
#9825000000
1!
1%
#9830000000
0!
0%
#9835000000
1!
1%
#9840000000
0!
0%
#9845000000
1!
1%
#9850000000
0!
0%
#9855000000
1!
1%
#9860000000
0!
0%
#9865000000
1!
1%
#9870000000
0!
0%
#9875000000
1!
1%
#9880000000
0!
0%
#9885000000
1!
1%
#9890000000
0!
0%
#9895000000
1!
1%
#9900000000
0!
0%
#9905000000
1!
1%
#9910000000
0!
0%
#9915000000
1!
1%
#9920000000
0!
0%
#9925000000
1!
1%
#9930000000
0!
0%
#9935000000
1!
1%
#9940000000
0!
0%
#9945000000
1!
1%
#9950000000
0!
0%
#9955000000
1!
1%
#9960000000
0!
0%
#9965000000
1!
1%
#9970000000
0!
0%
#9975000000
1!
1%
#9980000000
0!
0%
#9985000000
1!
1%
#9990000000
0!
0%
#9995000000
1!
1%
#10000000000
0!
0%
#10005000000
1!
1%
#10010000000
0!
0%
#10015000000
1!
1%
#10020000000
0!
0%
#10025000000
1!
1%
#10030000000
0!
0%
#10035000000
1!
1%
#10040000000
0!
0%
#10045000000
1!
1%
#10050000000
0!
0%
#10055000000
1!
1%
#10060000000
0!
0%
#10065000000
1!
1%
#10070000000
0!
0%
#10075000000
1!
1%
#10080000000
0!
0%
#10085000000
1!
1%
#10090000000
0!
0%
#10095000000
1!
1%
#10100000000
0!
0%
#10105000000
1!
1%
#10110000000
0!
0%
#10115000000
1!
1%
#10120000000
0!
0%
#10125000000
1!
1%
#10130000000
0!
0%
#10135000000
1!
1%
#10140000000
0!
0%
#10145000000
1!
1%
#10150000000
0!
0%
#10155000000
1!
1%
#10160000000
0!
0%
#10165000000
1!
1%
#10170000000
0!
0%
#10175000000
1!
1%
#10180000000
0!
0%
#10185000000
1!
1%
#10190000000
0!
0%
#10195000000
1!
1%
#10200000000
0!
0%
#10205000000
1!
1%
#10210000000
0!
0%
#10215000000
1!
1%
#10220000000
0!
0%
#10225000000
1!
1%
#10230000000
0!
0%
#10235000000
1!
1%
#10240000000
0!
0%
#10245000000
1!
1%
#10250000000
0!
0%
#10255000000
1!
1%
#10260000000
0!
0%
#10265000000
1!
1%
#10270000000
0!
0%
#10275000000
1!
1%
#10280000000
0!
0%
#10285000000
1!
1%
#10290000000
0!
0%
#10295000000
1!
1%
#10300000000
0!
0%
#10305000000
1!
1%
#10310000000
0!
0%
#10315000000
1!
1%
#10320000000
0!
0%
#10325000000
1!
1%
#10330000000
0!
0%
#10335000000
1!
1%
#10340000000
0!
0%
#10345000000
1!
1%
#10350000000
0!
0%
#10355000000
1!
1%
#10360000000
0!
0%
#10365000000
1!
1%
#10370000000
0!
0%
#10375000000
1!
1%
#10380000000
0!
0%
#10385000000
1!
1%
#10390000000
0!
0%
#10395000000
1!
1%
#10400000000
0!
0%
#10405000000
1!
1%
#10410000000
0!
0%
#10415000000
1!
1%
#10420000000
0!
0%
#10425000000
1!
1%
#10430000000
0!
0%
#10435000000
1!
1%
#10440000000
0!
0%
#10445000000
1!
1%
#10450000000
0!
0%
#10455000000
1!
1%
#10460000000
0!
0%
#10465000000
1!
1%
#10470000000
0!
0%
#10475000000
1!
1%
#10480000000
0!
0%
#10485000000
1!
1%
#10490000000
0!
0%
#10495000000
1!
1%
#10500000000
0!
0%
#10505000000
1!
1%
#10510000000
0!
0%
#10515000000
1!
1%
#10520000000
0!
0%
#10525000000
1!
1%
#10530000000
0!
0%
#10535000000
1!
1%
#10540000000
0!
0%
#10545000000
1!
1%
#10550000000
0!
0%
#10555000000
1!
1%
#10560000000
0!
0%
#10565000000
1!
1%
#10570000000
0!
0%
#10575000000
1!
1%
#10580000000
0!
0%
#10585000000
1!
1%
#10590000000
0!
0%
#10595000000
1!
1%
#10600000000
0!
0%
#10605000000
1!
1%
#10610000000
0!
0%
#10615000000
1!
1%
#10620000000
0!
0%
#10625000000
1!
1%
#10630000000
0!
0%
#10635000000
1!
1%
#10640000000
0!
0%
#10645000000
1!
1%
#10650000000
0!
0%
#10655000000
1!
1%
#10660000000
0!
0%
#10665000000
1!
1%
#10670000000
0!
0%
#10675000000
1!
1%
#10680000000
0!
0%
#10685000000
1!
1%
#10690000000
0!
0%
#10695000000
1!
1%
#10700000000
0!
0%
#10705000000
1!
1%
#10710000000
0!
0%
#10715000000
1!
1%
#10720000000
0!
0%
#10725000000
1!
1%
#10730000000
0!
0%
#10735000000
1!
1%
#10740000000
0!
0%
#10745000000
1!
1%
#10750000000
0!
0%
#10755000000
1!
1%
#10760000000
0!
0%
#10765000000
1!
1%
#10770000000
0!
0%
#10775000000
1!
1%
#10780000000
0!
0%
#10785000000
1!
1%
#10790000000
0!
0%
#10795000000
1!
1%
#10800000000
0!
0%
#10805000000
1!
1%
#10810000000
0!
0%
#10815000000
1!
1%
#10820000000
0!
0%
#10825000000
1!
1%
#10830000000
0!
0%
#10835000000
1!
1%
#10840000000
0!
0%
#10845000000
1!
1%
#10850000000
0!
0%
#10855000000
1!
1%
#10860000000
0!
0%
#10865000000
1!
1%
#10870000000
0!
0%
#10875000000
1!
1%
#10880000000
0!
0%
#10885000000
1!
1%
#10890000000
0!
0%
#10895000000
1!
1%
#10900000000
0!
0%
#10905000000
1!
1%
#10910000000
0!
0%
#10915000000
1!
1%
#10920000000
0!
0%
#10925000000
1!
1%
#10930000000
0!
0%
#10935000000
1!
1%
#10940000000
0!
0%
#10945000000
1!
1%
#10950000000
0!
0%
#10955000000
1!
1%
#10960000000
0!
0%
#10965000000
1!
1%
#10970000000
0!
0%
#10975000000
1!
1%
#10980000000
0!
0%
#10985000000
1!
1%
#10990000000
0!
0%
#10995000000
1!
1%
#11000000000
0!
0%
#11005000000
1!
1%
#11010000000
0!
0%
#11015000000
1!
1%
#11020000000
0!
0%
#11025000000
1!
1%
#11030000000
0!
0%
#11035000000
1!
1%
#11040000000
0!
0%
#11045000000
1!
1%
#11050000000
0!
0%
#11055000000
1!
1%
#11060000000
0!
0%
#11065000000
1!
1%
#11070000000
0!
0%
#11075000000
1!
1%
#11080000000
0!
0%
#11085000000
1!
1%
#11090000000
0!
0%
#11095000000
1!
1%
#11100000000
0!
0%
#11105000000
1!
1%
#11110000000
0!
0%
#11115000000
1!
1%
#11120000000
0!
0%
#11125000000
1!
1%
#11130000000
0!
0%
#11135000000
1!
1%
#11140000000
0!
0%
#11145000000
1!
1%
#11150000000
0!
0%
#11155000000
1!
1%
#11160000000
0!
0%
#11165000000
1!
1%
#11170000000
0!
0%
#11175000000
1!
1%
#11180000000
0!
0%
#11185000000
1!
1%
#11190000000
0!
0%
#11195000000
1!
1%
#11200000000
0!
0%
#11205000000
1!
1%
#11210000000
0!
0%
#11215000000
1!
1%
#11220000000
0!
0%
#11225000000
1!
1%
#11230000000
0!
0%
#11235000000
1!
1%
#11240000000
0!
0%
#11245000000
1!
1%
#11250000000
0!
0%
#11255000000
1!
1%
#11260000000
0!
0%
#11265000000
1!
1%
#11270000000
0!
0%
#11275000000
1!
1%
#11280000000
0!
0%
#11285000000
1!
1%
#11290000000
0!
0%
#11295000000
1!
1%
#11300000000
0!
0%
#11305000000
1!
1%
#11310000000
0!
0%
#11315000000
1!
1%
#11320000000
0!
0%
#11325000000
1!
1%
#11330000000
0!
0%
#11335000000
1!
1%
#11340000000
0!
0%
#11345000000
1!
1%
#11350000000
0!
0%
#11355000000
1!
1%
#11360000000
0!
0%
#11365000000
1!
1%
#11370000000
0!
0%
#11375000000
1!
1%
#11380000000
0!
0%
#11385000000
1!
1%
#11390000000
0!
0%
#11395000000
1!
1%
#11400000000
0!
0%
#11405000000
1!
1%
#11410000000
0!
0%
#11415000000
1!
1%
#11420000000
0!
0%
#11425000000
1!
1%
#11430000000
0!
0%
#11435000000
1!
1%
#11440000000
0!
0%
#11445000000
1!
1%
#11450000000
0!
0%
#11455000000
1!
1%
#11460000000
0!
0%
#11465000000
1!
1%
#11470000000
0!
0%
#11475000000
1!
1%
#11480000000
0!
0%
#11485000000
1!
1%
#11490000000
0!
0%
#11495000000
1!
1%
#11500000000
0!
0%
#11505000000
1!
1%
#11510000000
0!
0%
#11515000000
1!
1%
#11520000000
0!
0%
#11525000000
1!
1%
#11530000000
0!
0%
#11535000000
1!
1%
#11540000000
0!
0%
#11545000000
1!
1%
#11550000000
0!
0%
#11555000000
1!
1%
#11560000000
0!
0%
#11565000000
1!
1%
#11570000000
0!
0%
#11575000000
1!
1%
#11580000000
0!
0%
#11585000000
1!
1%
#11590000000
0!
0%
#11595000000
1!
1%
#11600000000
0!
0%
#11605000000
1!
1%
#11610000000
0!
0%
#11615000000
1!
1%
#11620000000
0!
0%
#11625000000
1!
1%
#11630000000
0!
0%
#11635000000
1!
1%
#11640000000
0!
0%
#11645000000
1!
1%
#11650000000
0!
0%
#11655000000
1!
1%
#11660000000
0!
0%
#11665000000
1!
1%
#11670000000
0!
0%
#11675000000
1!
1%
#11680000000
0!
0%
#11685000000
1!
1%
#11690000000
0!
0%
#11695000000
1!
1%
#11700000000
0!
0%
#11705000000
1!
1%
#11710000000
0!
0%
#11715000000
1!
1%
#11720000000
0!
0%
#11725000000
1!
1%
#11730000000
0!
0%
#11735000000
1!
1%
#11740000000
0!
0%
#11745000000
1!
1%
#11750000000
0!
0%
#11755000000
1!
1%
#11760000000
0!
0%
#11765000000
1!
1%
#11770000000
0!
0%
#11775000000
1!
1%
#11780000000
0!
0%
#11785000000
1!
1%
#11790000000
0!
0%
#11795000000
1!
1%
#11800000000
0!
0%
#11805000000
1!
1%
#11810000000
0!
0%
#11815000000
1!
1%
#11820000000
0!
0%
#11825000000
1!
1%
#11830000000
0!
0%
#11835000000
1!
1%
#11840000000
0!
0%
#11845000000
1!
1%
#11850000000
0!
0%
#11855000000
1!
1%
#11860000000
0!
0%
#11865000000
1!
1%
#11870000000
0!
0%
#11875000000
1!
1%
#11880000000
0!
0%
#11885000000
1!
1%
#11890000000
0!
0%
#11895000000
1!
1%
#11900000000
0!
0%
#11905000000
1!
1%
#11910000000
0!
0%
#11915000000
1!
1%
#11920000000
0!
0%
#11925000000
1!
1%
#11930000000
0!
0%
#11935000000
1!
1%
#11940000000
0!
0%
#11945000000
1!
1%
#11950000000
0!
0%
#11955000000
1!
1%
#11960000000
0!
0%
#11965000000
1!
1%
#11970000000
0!
0%
#11975000000
1!
1%
#11980000000
0!
0%
#11985000000
1!
1%
#11990000000
0!
0%
#11995000000
1!
1%
#12000000000
0!
0%
#12005000000
1!
1%
#12010000000
0!
0%
#12015000000
1!
1%
#12020000000
0!
0%
#12025000000
1!
1%
#12030000000
0!
0%
#12035000000
1!
1%
#12040000000
0!
0%
#12045000000
1!
1%
#12050000000
0!
0%
#12055000000
1!
1%
#12060000000
0!
0%
#12065000000
1!
1%
#12070000000
0!
0%
#12075000000
1!
1%
#12080000000
0!
0%
#12085000000
1!
1%
#12090000000
0!
0%
#12095000000
1!
1%
#12100000000
0!
0%
#12105000000
1!
1%
#12110000000
0!
0%
#12115000000
1!
1%
#12120000000
0!
0%
#12125000000
1!
1%
#12130000000
0!
0%
#12135000000
1!
1%
#12140000000
0!
0%
#12145000000
1!
1%
#12150000000
0!
0%
#12155000000
1!
1%
#12160000000
0!
0%
#12165000000
1!
1%
#12170000000
0!
0%
#12175000000
1!
1%
#12180000000
0!
0%
#12185000000
1!
1%
#12190000000
0!
0%
#12195000000
1!
1%
#12200000000
0!
0%
#12205000000
1!
1%
#12210000000
0!
0%
#12215000000
1!
1%
#12220000000
0!
0%
#12225000000
1!
1%
#12230000000
0!
0%
#12235000000
1!
1%
#12240000000
0!
0%
#12245000000
1!
1%
#12250000000
0!
0%
#12255000000
1!
1%
#12260000000
0!
0%
#12265000000
1!
1%
#12270000000
0!
0%
#12275000000
1!
1%
#12280000000
0!
0%
#12285000000
1!
1%
#12290000000
0!
0%
#12295000000
1!
1%
#12300000000
0!
0%
#12305000000
1!
1%
#12310000000
0!
0%
#12315000000
1!
1%
#12320000000
0!
0%
#12325000000
1!
1%
#12330000000
0!
0%
#12335000000
1!
1%
#12340000000
0!
0%
#12345000000
1!
1%
#12350000000
0!
0%
#12355000000
1!
1%
#12360000000
0!
0%
#12365000000
1!
1%
#12370000000
0!
0%
#12375000000
1!
1%
#12380000000
0!
0%
#12385000000
1!
1%
#12390000000
0!
0%
#12395000000
1!
1%
#12400000000
0!
0%
#12405000000
1!
1%
#12410000000
0!
0%
#12415000000
1!
1%
#12420000000
0!
0%
#12425000000
1!
1%
#12430000000
0!
0%
#12435000000
1!
1%
#12440000000
0!
0%
#12445000000
1!
1%
#12450000000
0!
0%
#12455000000
1!
1%
#12460000000
0!
0%
#12465000000
1!
1%
#12470000000
0!
0%
#12475000000
1!
1%
#12480000000
0!
0%
#12485000000
1!
1%
#12490000000
0!
0%
#12495000000
1!
1%
#12500000000
0!
0%
#12505000000
1!
1%
#12510000000
0!
0%
#12515000000
1!
1%
#12520000000
0!
0%
#12525000000
1!
1%
#12530000000
0!
0%
#12535000000
1!
1%
#12540000000
0!
0%
#12545000000
1!
1%
#12550000000
0!
0%
#12555000000
1!
1%
#12560000000
0!
0%
#12565000000
1!
1%
#12570000000
0!
0%
#12575000000
1!
1%
#12580000000
0!
0%
#12585000000
1!
1%
#12590000000
0!
0%
#12595000000
1!
1%
#12600000000
0!
0%
#12605000000
1!
1%
#12610000000
0!
0%
#12615000000
1!
1%
#12620000000
0!
0%
#12625000000
1!
1%
#12630000000
0!
0%
#12635000000
1!
1%
#12640000000
0!
0%
#12645000000
1!
1%
#12650000000
0!
0%
#12655000000
1!
1%
#12660000000
0!
0%
#12665000000
1!
1%
#12670000000
0!
0%
#12675000000
1!
1%
#12680000000
0!
0%
#12685000000
1!
1%
#12690000000
0!
0%
#12695000000
1!
1%
#12700000000
0!
0%
#12705000000
1!
1%
#12710000000
0!
0%
#12715000000
1!
1%
#12720000000
0!
0%
#12725000000
1!
1%
#12730000000
0!
0%
#12735000000
1!
1%
#12740000000
0!
0%
#12745000000
1!
1%
#12750000000
0!
0%
#12755000000
1!
1%
#12760000000
0!
0%
#12765000000
1!
1%
#12770000000
0!
0%
#12775000000
1!
1%
#12780000000
0!
0%
#12785000000
1!
1%
#12790000000
0!
0%
#12795000000
1!
1%
#12800000000
0!
0%
#12805000000
1!
1%
#12810000000
0!
0%
#12815000000
1!
1%
#12820000000
0!
0%
#12825000000
1!
1%
#12830000000
0!
0%
#12835000000
1!
1%
#12840000000
0!
0%
#12845000000
1!
1%
#12850000000
0!
0%
#12855000000
1!
1%
#12860000000
0!
0%
#12865000000
1!
1%
#12870000000
0!
0%
#12875000000
1!
1%
#12880000000
0!
0%
#12885000000
1!
1%
#12890000000
0!
0%
#12895000000
1!
1%
#12900000000
0!
0%
#12905000000
1!
1%
#12910000000
0!
0%
#12915000000
1!
1%
#12920000000
0!
0%
#12925000000
1!
1%
#12930000000
0!
0%
#12935000000
1!
1%
#12940000000
0!
0%
#12945000000
1!
1%
#12950000000
0!
0%
#12955000000
1!
1%
#12960000000
0!
0%
#12965000000
1!
1%
#12970000000
0!
0%
#12975000000
1!
1%
#12980000000
0!
0%
#12985000000
1!
1%
#12990000000
0!
0%
#12995000000
1!
1%
#13000000000
0!
0%
#13005000000
1!
1%
#13010000000
0!
0%
#13015000000
1!
1%
#13020000000
0!
0%
#13025000000
1!
1%
#13030000000
0!
0%
#13035000000
1!
1%
#13040000000
0!
0%
#13045000000
1!
1%
#13050000000
0!
0%
#13055000000
1!
1%
#13060000000
0!
0%
#13065000000
1!
1%
#13070000000
0!
0%
#13075000000
1!
1%
#13080000000
0!
0%
#13085000000
1!
1%
#13090000000
0!
0%
#13095000000
1!
1%
#13100000000
0!
0%
#13105000000
1!
1%
#13110000000
0!
0%
#13115000000
1!
1%
#13120000000
0!
0%
#13125000000
1!
1%
#13130000000
0!
0%
#13135000000
1!
1%
#13140000000
0!
0%
#13145000000
1!
1%
#13150000000
0!
0%
#13155000000
1!
1%
#13160000000
0!
0%
#13165000000
1!
1%
#13170000000
0!
0%
#13175000000
1!
1%
#13180000000
0!
0%
#13185000000
1!
1%
#13190000000
0!
0%
#13195000000
1!
1%
#13200000000
0!
0%
#13205000000
1!
1%
#13210000000
0!
0%
#13215000000
1!
1%
#13220000000
0!
0%
#13225000000
1!
1%
#13230000000
0!
0%
#13235000000
1!
1%
#13240000000
0!
0%
#13245000000
1!
1%
#13250000000
0!
0%
#13255000000
1!
1%
#13260000000
0!
0%
#13265000000
1!
1%
#13270000000
0!
0%
#13275000000
1!
1%
#13280000000
0!
0%
#13285000000
1!
1%
#13290000000
0!
0%
#13295000000
1!
1%
#13300000000
0!
0%
#13305000000
1!
1%
#13310000000
0!
0%
#13315000000
1!
1%
#13320000000
0!
0%
#13325000000
1!
1%
#13330000000
0!
0%
#13335000000
1!
1%
#13340000000
0!
0%
#13345000000
1!
1%
#13350000000
0!
0%
#13355000000
1!
1%
#13360000000
0!
0%
#13365000000
1!
1%
#13370000000
0!
0%
#13375000000
1!
1%
#13380000000
0!
0%
#13385000000
1!
1%
#13390000000
0!
0%
#13395000000
1!
1%
#13400000000
0!
0%
#13405000000
1!
1%
#13410000000
0!
0%
#13415000000
1!
1%
#13420000000
0!
0%
#13425000000
1!
1%
#13430000000
0!
0%
#13435000000
1!
1%
#13440000000
0!
0%
#13445000000
1!
1%
#13450000000
0!
0%
#13455000000
1!
1%
#13460000000
0!
0%
#13465000000
1!
1%
#13470000000
0!
0%
#13475000000
1!
1%
#13480000000
0!
0%
#13485000000
1!
1%
#13490000000
0!
0%
#13495000000
1!
1%
#13500000000
0!
0%
#13505000000
1!
1%
#13510000000
0!
0%
#13515000000
1!
1%
#13520000000
0!
0%
#13525000000
1!
1%
#13530000000
0!
0%
#13535000000
1!
1%
#13540000000
0!
0%
#13545000000
1!
1%
#13550000000
0!
0%
#13555000000
1!
1%
#13560000000
0!
0%
#13565000000
1!
1%
#13570000000
0!
0%
#13575000000
1!
1%
#13580000000
0!
0%
#13585000000
1!
1%
#13590000000
0!
0%
#13595000000
1!
1%
#13600000000
0!
0%
#13605000000
1!
1%
#13610000000
0!
0%
#13615000000
1!
1%
#13620000000
0!
0%
#13625000000
1!
1%
#13630000000
0!
0%
#13635000000
1!
1%
#13640000000
0!
0%
#13645000000
1!
1%
#13650000000
0!
0%
#13655000000
1!
1%
#13660000000
0!
0%
#13665000000
1!
1%
#13670000000
0!
0%
#13675000000
1!
1%
#13680000000
0!
0%
#13685000000
1!
1%
#13690000000
0!
0%
#13695000000
1!
1%
#13700000000
0!
0%
#13705000000
1!
1%
#13710000000
0!
0%
#13715000000
1!
1%
#13720000000
0!
0%
#13725000000
1!
1%
#13730000000
0!
0%
#13735000000
1!
1%
#13740000000
0!
0%
#13745000000
1!
1%
#13750000000
0!
0%
#13755000000
1!
1%
#13760000000
0!
0%
#13765000000
1!
1%
#13770000000
0!
0%
#13775000000
1!
1%
#13780000000
0!
0%
#13785000000
1!
1%
#13790000000
0!
0%
#13795000000
1!
1%
#13800000000
0!
0%
#13805000000
1!
1%
#13810000000
0!
0%
#13815000000
1!
1%
#13820000000
0!
0%
#13825000000
1!
1%
#13830000000
0!
0%
#13835000000
1!
1%
#13840000000
0!
0%
#13845000000
1!
1%
#13850000000
0!
0%
#13855000000
1!
1%
#13860000000
0!
0%
#13865000000
1!
1%
#13870000000
0!
0%
#13875000000
1!
1%
#13880000000
0!
0%
#13885000000
1!
1%
#13890000000
0!
0%
#13895000000
1!
1%
#13900000000
0!
0%
#13905000000
1!
1%
#13910000000
0!
0%
#13915000000
1!
1%
#13920000000
0!
0%
#13925000000
1!
1%
#13930000000
0!
0%
#13935000000
1!
1%
#13940000000
0!
0%
#13945000000
1!
1%
#13950000000
0!
0%
#13955000000
1!
1%
#13960000000
0!
0%
#13965000000
1!
1%
#13970000000
0!
0%
#13975000000
1!
1%
#13980000000
0!
0%
#13985000000
1!
1%
#13990000000
0!
0%
#13995000000
1!
1%
#14000000000
0!
0%
#14005000000
1!
1%
#14010000000
0!
0%
#14015000000
1!
1%
#14020000000
0!
0%
#14025000000
1!
1%
#14030000000
0!
0%
#14035000000
1!
1%
#14040000000
0!
0%
#14045000000
1!
1%
#14050000000
0!
0%
#14055000000
1!
1%
#14060000000
0!
0%
#14065000000
1!
1%
#14070000000
0!
0%
#14075000000
1!
1%
#14080000000
0!
0%
#14085000000
1!
1%
#14090000000
0!
0%
#14095000000
1!
1%
#14100000000
0!
0%
#14105000000
1!
1%
#14110000000
0!
0%
#14115000000
1!
1%
#14120000000
0!
0%
#14125000000
1!
1%
#14130000000
0!
0%
#14135000000
1!
1%
#14140000000
0!
0%
#14145000000
1!
1%
#14150000000
0!
0%
#14155000000
1!
1%
#14160000000
0!
0%
#14165000000
1!
1%
#14170000000
0!
0%
#14175000000
1!
1%
#14180000000
0!
0%
#14185000000
1!
1%
#14190000000
0!
0%
#14195000000
1!
1%
#14200000000
0!
0%
#14205000000
1!
1%
#14210000000
0!
0%
#14215000000
1!
1%
#14220000000
0!
0%
#14225000000
1!
1%
#14230000000
0!
0%
#14235000000
1!
1%
#14240000000
0!
0%
#14245000000
1!
1%
#14250000000
0!
0%
#14255000000
1!
1%
#14260000000
0!
0%
#14265000000
1!
1%
#14270000000
0!
0%
#14275000000
1!
1%
#14280000000
0!
0%
#14285000000
1!
1%
#14290000000
0!
0%
#14295000000
1!
1%
#14300000000
0!
0%
#14305000000
1!
1%
#14310000000
0!
0%
#14315000000
1!
1%
#14320000000
0!
0%
#14325000000
1!
1%
#14330000000
0!
0%
#14335000000
1!
1%
#14340000000
0!
0%
#14345000000
1!
1%
#14350000000
0!
0%
#14355000000
1!
1%
#14360000000
0!
0%
#14365000000
1!
1%
#14370000000
0!
0%
#14375000000
1!
1%
#14380000000
0!
0%
#14385000000
1!
1%
#14390000000
0!
0%
#14395000000
1!
1%
#14400000000
0!
0%
#14405000000
1!
1%
#14410000000
0!
0%
#14415000000
1!
1%
#14420000000
0!
0%
#14425000000
1!
1%
#14430000000
0!
0%
#14435000000
1!
1%
#14440000000
0!
0%
#14445000000
1!
1%
#14450000000
0!
0%
#14455000000
1!
1%
#14460000000
0!
0%
#14465000000
1!
1%
#14470000000
0!
0%
#14475000000
1!
1%
#14480000000
0!
0%
#14485000000
1!
1%
#14490000000
0!
0%
#14495000000
1!
1%
#14500000000
0!
0%
#14505000000
1!
1%
#14510000000
0!
0%
#14515000000
1!
1%
#14520000000
0!
0%
#14525000000
1!
1%
#14530000000
0!
0%
#14535000000
1!
1%
#14540000000
0!
0%
#14545000000
1!
1%
#14550000000
0!
0%
#14555000000
1!
1%
#14560000000
0!
0%
#14565000000
1!
1%
#14570000000
0!
0%
#14575000000
1!
1%
#14580000000
0!
0%
#14585000000
1!
1%
#14590000000
0!
0%
#14595000000
1!
1%
#14600000000
0!
0%
#14605000000
1!
1%
#14610000000
0!
0%
#14615000000
1!
1%
#14620000000
0!
0%
#14625000000
1!
1%
#14630000000
0!
0%
#14635000000
1!
1%
#14640000000
0!
0%
#14645000000
1!
1%
#14650000000
0!
0%
#14655000000
1!
1%
#14660000000
0!
0%
#14665000000
1!
1%
#14670000000
0!
0%
#14675000000
1!
1%
#14680000000
0!
0%
#14685000000
1!
1%
#14690000000
0!
0%
#14695000000
1!
1%
#14700000000
0!
0%
#14705000000
1!
1%
#14710000000
0!
0%
#14715000000
1!
1%
#14720000000
0!
0%
#14725000000
1!
1%
#14730000000
0!
0%
#14735000000
1!
1%
#14740000000
0!
0%
#14745000000
1!
1%
#14750000000
0!
0%
#14755000000
1!
1%
#14760000000
0!
0%
#14765000000
1!
1%
#14770000000
0!
0%
#14775000000
1!
1%
#14780000000
0!
0%
#14785000000
1!
1%
#14790000000
0!
0%
#14795000000
1!
1%
#14800000000
0!
0%
#14805000000
1!
1%
#14810000000
0!
0%
#14815000000
1!
1%
#14820000000
0!
0%
#14825000000
1!
1%
#14830000000
0!
0%
#14835000000
1!
1%
#14840000000
0!
0%
#14845000000
1!
1%
#14850000000
0!
0%
#14855000000
1!
1%
#14860000000
0!
0%
#14865000000
1!
1%
#14870000000
0!
0%
#14875000000
1!
1%
#14880000000
0!
0%
#14885000000
1!
1%
#14890000000
0!
0%
#14895000000
1!
1%
#14900000000
0!
0%
#14905000000
1!
1%
#14910000000
0!
0%
#14915000000
1!
1%
#14920000000
0!
0%
#14925000000
1!
1%
#14930000000
0!
0%
#14935000000
1!
1%
#14940000000
0!
0%
#14945000000
1!
1%
#14950000000
0!
0%
#14955000000
1!
1%
#14960000000
0!
0%
#14965000000
1!
1%
#14970000000
0!
0%
#14975000000
1!
1%
#14980000000
0!
0%
#14985000000
1!
1%
#14990000000
0!
0%
#14995000000
1!
1%
#15000000000
0!
0%
#15005000000
1!
1%
#15010000000
0!
0%
#15015000000
1!
1%
#15020000000
0!
0%
#15025000000
1!
1%
#15030000000
0!
0%
#15035000000
1!
1%
#15040000000
0!
0%
#15045000000
1!
1%
#15050000000
0!
0%
#15055000000
1!
1%
#15060000000
0!
0%
#15065000000
1!
1%
#15070000000
0!
0%
#15075000000
1!
1%
#15080000000
0!
0%
#15085000000
1!
1%
#15090000000
0!
0%
#15095000000
1!
1%
#15100000000
0!
0%
#15105000000
1!
1%
#15110000000
0!
0%
#15115000000
1!
1%
#15120000000
0!
0%
#15125000000
1!
1%
#15130000000
0!
0%
#15135000000
1!
1%
#15140000000
0!
0%
#15145000000
1!
1%
#15150000000
0!
0%
#15155000000
1!
1%
#15160000000
0!
0%
#15165000000
1!
1%
#15170000000
0!
0%
#15175000000
1!
1%
#15180000000
0!
0%
#15185000000
1!
1%
#15190000000
0!
0%
#15195000000
1!
1%
#15200000000
0!
0%
#15205000000
1!
1%
#15210000000
0!
0%
#15215000000
1!
1%
#15220000000
0!
0%
#15225000000
1!
1%
#15230000000
0!
0%
#15235000000
1!
1%
#15240000000
0!
0%
#15245000000
1!
1%
#15250000000
0!
0%
#15255000000
1!
1%
#15260000000
0!
0%
#15265000000
1!
1%
#15270000000
0!
0%
#15275000000
1!
1%
#15280000000
0!
0%
#15285000000
1!
1%
#15290000000
0!
0%
#15295000000
1!
1%
#15300000000
0!
0%
#15305000000
1!
1%
#15310000000
0!
0%
#15315000000
1!
1%
#15320000000
0!
0%
#15325000000
1!
1%
#15330000000
0!
0%
#15335000000
1!
1%
#15340000000
0!
0%
#15345000000
1!
1%
#15350000000
0!
0%
#15355000000
1!
1%
#15360000000
0!
0%
#15365000000
1!
1%
#15370000000
0!
0%
#15375000000
1!
1%
#15380000000
0!
0%
#15385000000
1!
1%
#15390000000
0!
0%
#15395000000
1!
1%
#15400000000
0!
0%
#15405000000
1!
1%
#15410000000
0!
0%
#15415000000
1!
1%
#15420000000
0!
0%
#15425000000
1!
1%
#15430000000
0!
0%
#15435000000
1!
1%
#15440000000
0!
0%
#15445000000
1!
1%
#15450000000
0!
0%
#15455000000
1!
1%
#15460000000
0!
0%
#15465000000
1!
1%
#15470000000
0!
0%
#15475000000
1!
1%
#15480000000
0!
0%
#15485000000
1!
1%
#15490000000
0!
0%
#15495000000
1!
1%
#15500000000
0!
0%
#15505000000
1!
1%
#15510000000
0!
0%
#15515000000
1!
1%
#15520000000
0!
0%
#15525000000
1!
1%
#15530000000
0!
0%
#15535000000
1!
1%
#15540000000
0!
0%
#15545000000
1!
1%
#15550000000
0!
0%
#15555000000
1!
1%
#15560000000
0!
0%
#15565000000
1!
1%
#15570000000
0!
0%
#15575000000
1!
1%
#15580000000
0!
0%
#15585000000
1!
1%
#15590000000
0!
0%
#15595000000
1!
1%
#15600000000
0!
0%
#15605000000
1!
1%
#15610000000
0!
0%
#15615000000
1!
1%
#15620000000
0!
0%
#15625000000
1!
1%
#15630000000
0!
0%
#15635000000
1!
1%
#15640000000
0!
0%
#15645000000
1!
1%
#15650000000
0!
0%
#15655000000
1!
1%
#15660000000
0!
0%
#15665000000
1!
1%
#15670000000
0!
0%
#15675000000
1!
1%
#15680000000
0!
0%
#15685000000
1!
1%
#15690000000
0!
0%
#15695000000
1!
1%
#15700000000
0!
0%
#15705000000
1!
1%
#15710000000
0!
0%
#15715000000
1!
1%
#15720000000
0!
0%
#15725000000
1!
1%
#15730000000
0!
0%
#15735000000
1!
1%
#15740000000
0!
0%
#15745000000
1!
1%
#15750000000
0!
0%
#15755000000
1!
1%
#15760000000
0!
0%
#15765000000
1!
1%
#15770000000
0!
0%
#15775000000
1!
1%
#15780000000
0!
0%
#15785000000
1!
1%
#15790000000
0!
0%
#15795000000
1!
1%
#15800000000
0!
0%
#15805000000
1!
1%
#15810000000
0!
0%
#15815000000
1!
1%
#15820000000
0!
0%
#15825000000
1!
1%
#15830000000
0!
0%
#15835000000
1!
1%
#15840000000
0!
0%
#15845000000
1!
1%
#15850000000
0!
0%
#15855000000
1!
1%
#15860000000
0!
0%
#15865000000
1!
1%
#15870000000
0!
0%
#15875000000
1!
1%
#15880000000
0!
0%
#15885000000
1!
1%
#15890000000
0!
0%
#15895000000
1!
1%
#15900000000
0!
0%
#15905000000
1!
1%
#15910000000
0!
0%
#15915000000
1!
1%
#15920000000
0!
0%
#15925000000
1!
1%
#15930000000
0!
0%
#15935000000
1!
1%
#15940000000
0!
0%
#15945000000
1!
1%
#15950000000
0!
0%
#15955000000
1!
1%
#15960000000
0!
0%
#15965000000
1!
1%
#15970000000
0!
0%
#15975000000
1!
1%
#15980000000
0!
0%
#15985000000
1!
1%
#15990000000
0!
0%
#15995000000
1!
1%
#16000000000
0!
0%
#16005000000
1!
1%
#16010000000
0!
0%
#16015000000
1!
1%
#16020000000
0!
0%
#16025000000
1!
1%
#16030000000
0!
0%
#16035000000
1!
1%
#16040000000
0!
0%
#16045000000
1!
1%
#16050000000
0!
0%
#16055000000
1!
1%
#16060000000
0!
0%
#16065000000
1!
1%
#16070000000
0!
0%
#16075000000
1!
1%
#16080000000
0!
0%
#16085000000
1!
1%
#16090000000
0!
0%
#16095000000
1!
1%
#16100000000
0!
0%
#16105000000
1!
1%
#16110000000
0!
0%
#16115000000
1!
1%
#16120000000
0!
0%
#16125000000
1!
1%
#16130000000
0!
0%
#16135000000
1!
1%
#16140000000
0!
0%
#16145000000
1!
1%
#16150000000
0!
0%
#16155000000
1!
1%
#16160000000
0!
0%
#16165000000
1!
1%
#16170000000
0!
0%
#16175000000
1!
1%
#16180000000
0!
0%
#16185000000
1!
1%
#16190000000
0!
0%
#16195000000
1!
1%
#16200000000
0!
0%
#16205000000
1!
1%
#16210000000
0!
0%
#16215000000
1!
1%
#16220000000
0!
0%
#16225000000
1!
1%
#16230000000
0!
0%
#16235000000
1!
1%
#16240000000
0!
0%
#16245000000
1!
1%
#16250000000
0!
0%
#16255000000
1!
1%
#16260000000
0!
0%
#16265000000
1!
1%
#16270000000
0!
0%
#16275000000
1!
1%
#16280000000
0!
0%
#16285000000
1!
1%
#16290000000
0!
0%
#16295000000
1!
1%
#16300000000
0!
0%
#16305000000
1!
1%
#16310000000
0!
0%
#16315000000
1!
1%
#16320000000
0!
0%
#16325000000
1!
1%
#16330000000
0!
0%
#16335000000
1!
1%
#16340000000
0!
0%
#16345000000
1!
1%
#16350000000
0!
0%
#16355000000
1!
1%
#16360000000
0!
0%
#16365000000
1!
1%
#16370000000
0!
0%
#16375000000
1!
1%
#16380000000
0!
0%
#16385000000
1!
1%
#16390000000
0!
0%
#16395000000
1!
1%
#16400000000
0!
0%
#16405000000
1!
1%
#16410000000
0!
0%
#16415000000
1!
1%
#16420000000
0!
0%
#16425000000
1!
1%
#16430000000
0!
0%
#16435000000
1!
1%
#16440000000
0!
0%
#16445000000
1!
1%
#16450000000
0!
0%
#16455000000
1!
1%
#16460000000
0!
0%
#16465000000
1!
1%
#16470000000
0!
0%
#16475000000
1!
1%
#16480000000
0!
0%
#16485000000
1!
1%
#16490000000
0!
0%
#16495000000
1!
1%
#16500000000
0!
0%
#16505000000
1!
1%
#16510000000
0!
0%
#16515000000
1!
1%
#16520000000
0!
0%
#16525000000
1!
1%
#16530000000
0!
0%
#16535000000
1!
1%
#16540000000
0!
0%
#16545000000
1!
1%
#16550000000
0!
0%
#16555000000
1!
1%
#16560000000
0!
0%
#16565000000
1!
1%
#16570000000
0!
0%
#16575000000
1!
1%
#16580000000
0!
0%
#16585000000
1!
1%
#16590000000
0!
0%
#16595000000
1!
1%
#16600000000
0!
0%
#16605000000
1!
1%
#16610000000
0!
0%
#16615000000
1!
1%
#16620000000
0!
0%
#16625000000
1!
1%
#16630000000
0!
0%
#16635000000
1!
1%
#16640000000
0!
0%
#16645000000
1!
1%
#16650000000
0!
0%
#16655000000
1!
1%
#16660000000
0!
0%
#16665000000
1!
1%
#16670000000
0!
0%
#16675000000
1!
1%
#16680000000
0!
0%
#16685000000
1!
1%
#16690000000
0!
0%
#16695000000
1!
1%
#16700000000
0!
0%
#16705000000
1!
1%
#16710000000
0!
0%
#16715000000
1!
1%
#16720000000
0!
0%
#16725000000
1!
1%
#16730000000
0!
0%
#16735000000
1!
1%
#16740000000
0!
0%
#16745000000
1!
1%
#16750000000
0!
0%
#16755000000
1!
1%
#16760000000
0!
0%
#16765000000
1!
1%
#16770000000
0!
0%
#16775000000
1!
1%
#16780000000
0!
0%
#16785000000
1!
1%
#16790000000
0!
0%
#16795000000
1!
1%
#16800000000
0!
0%
#16805000000
1!
1%
#16810000000
0!
0%
#16815000000
1!
1%
#16820000000
0!
0%
#16825000000
1!
1%
#16830000000
0!
0%
#16835000000
1!
1%
#16840000000
0!
0%
#16845000000
1!
1%
#16850000000
0!
0%
#16855000000
1!
1%
#16860000000
0!
0%
#16865000000
1!
1%
#16870000000
0!
0%
#16875000000
1!
1%
#16880000000
0!
0%
#16885000000
1!
1%
#16890000000
0!
0%
#16895000000
1!
1%
#16900000000
0!
0%
#16905000000
1!
1%
#16910000000
0!
0%
#16915000000
1!
1%
#16920000000
0!
0%
#16925000000
1!
1%
#16930000000
0!
0%
#16935000000
1!
1%
#16940000000
0!
0%
#16945000000
1!
1%
#16950000000
0!
0%
#16955000000
1!
1%
#16960000000
0!
0%
#16965000000
1!
1%
#16970000000
0!
0%
#16975000000
1!
1%
#16980000000
0!
0%
#16985000000
1!
1%
#16990000000
0!
0%
#16995000000
1!
1%
#17000000000
0!
0%
#17005000000
1!
1%
#17010000000
0!
0%
#17015000000
1!
1%
#17020000000
0!
0%
#17025000000
1!
1%
#17030000000
0!
0%
#17035000000
1!
1%
#17040000000
0!
0%
#17045000000
1!
1%
#17050000000
0!
0%
#17055000000
1!
1%
#17060000000
0!
0%
#17065000000
1!
1%
#17070000000
0!
0%
#17075000000
1!
1%
#17080000000
0!
0%
#17085000000
1!
1%
#17090000000
0!
0%
#17095000000
1!
1%
#17100000000
0!
0%
#17105000000
1!
1%
#17110000000
0!
0%
#17115000000
1!
1%
#17120000000
0!
0%
#17125000000
1!
1%
#17130000000
0!
0%
#17135000000
1!
1%
#17140000000
0!
0%
#17145000000
1!
1%
#17150000000
0!
0%
#17155000000
1!
1%
#17160000000
0!
0%
#17165000000
1!
1%
#17170000000
0!
0%
#17175000000
1!
1%
#17180000000
0!
0%
#17185000000
1!
1%
#17190000000
0!
0%
#17195000000
1!
1%
#17200000000
0!
0%
#17205000000
1!
1%
#17210000000
0!
0%
#17215000000
1!
1%
#17220000000
0!
0%
#17225000000
1!
1%
#17230000000
0!
0%
#17235000000
1!
1%
#17240000000
0!
0%
#17245000000
1!
1%
#17250000000
0!
0%
#17255000000
1!
1%
#17260000000
0!
0%
#17265000000
1!
1%
#17270000000
0!
0%
#17275000000
1!
1%
#17280000000
0!
0%
#17285000000
1!
1%
#17290000000
0!
0%
#17295000000
1!
1%
#17300000000
0!
0%
#17305000000
1!
1%
#17310000000
0!
0%
#17315000000
1!
1%
#17320000000
0!
0%
#17325000000
1!
1%
#17330000000
0!
0%
#17335000000
1!
1%
#17340000000
0!
0%
#17345000000
1!
1%
#17350000000
0!
0%
#17355000000
1!
1%
#17360000000
0!
0%
#17365000000
1!
1%
#17370000000
0!
0%
#17375000000
1!
1%
#17380000000
0!
0%
#17385000000
1!
1%
#17390000000
0!
0%
#17395000000
1!
1%
#17400000000
0!
0%
#17405000000
1!
1%
#17410000000
0!
0%
#17415000000
1!
1%
#17420000000
0!
0%
#17425000000
1!
1%
#17430000000
0!
0%
#17435000000
1!
1%
#17440000000
0!
0%
#17445000000
1!
1%
#17450000000
0!
0%
#17455000000
1!
1%
#17460000000
0!
0%
#17465000000
1!
1%
#17470000000
0!
0%
#17475000000
1!
1%
#17480000000
0!
0%
#17485000000
1!
1%
#17490000000
0!
0%
#17495000000
1!
1%
#17500000000
0!
0%
#17505000000
1!
1%
#17510000000
0!
0%
#17515000000
1!
1%
#17520000000
0!
0%
#17525000000
1!
1%
#17530000000
0!
0%
#17535000000
1!
1%
#17540000000
0!
0%
#17545000000
1!
1%
#17550000000
0!
0%
#17555000000
1!
1%
#17560000000
0!
0%
#17565000000
1!
1%
#17570000000
0!
0%
#17575000000
1!
1%
#17580000000
0!
0%
#17585000000
1!
1%
#17590000000
0!
0%
#17595000000
1!
1%
#17600000000
0!
0%
#17605000000
1!
1%
#17610000000
0!
0%
#17615000000
1!
1%
#17620000000
0!
0%
#17625000000
1!
1%
#17630000000
0!
0%
#17635000000
1!
1%
#17640000000
0!
0%
#17645000000
1!
1%
#17650000000
0!
0%
#17655000000
1!
1%
#17660000000
0!
0%
#17665000000
1!
1%
#17670000000
0!
0%
#17675000000
1!
1%
#17680000000
0!
0%
#17685000000
1!
1%
#17690000000
0!
0%
#17695000000
1!
1%
#17700000000
0!
0%
#17705000000
1!
1%
#17710000000
0!
0%
#17715000000
1!
1%
#17720000000
0!
0%
#17725000000
1!
1%
#17730000000
0!
0%
#17735000000
1!
1%
#17740000000
0!
0%
#17745000000
1!
1%
#17750000000
0!
0%
#17755000000
1!
1%
#17760000000
0!
0%
#17765000000
1!
1%
#17770000000
0!
0%
#17775000000
1!
1%
#17780000000
0!
0%
#17785000000
1!
1%
#17790000000
0!
0%
#17795000000
1!
1%
#17800000000
0!
0%
#17805000000
1!
1%
#17810000000
0!
0%
#17815000000
1!
1%
#17820000000
0!
0%
#17825000000
1!
1%
#17830000000
0!
0%
#17835000000
1!
1%
#17840000000
0!
0%
#17845000000
1!
1%
#17850000000
0!
0%
#17855000000
1!
1%
#17860000000
0!
0%
#17865000000
1!
1%
#17870000000
0!
0%
#17875000000
1!
1%
#17880000000
0!
0%
#17885000000
1!
1%
#17890000000
0!
0%
#17895000000
1!
1%
#17900000000
0!
0%
#17905000000
1!
1%
#17910000000
0!
0%
#17915000000
1!
1%
#17920000000
0!
0%
#17925000000
1!
1%
#17930000000
0!
0%
#17935000000
1!
1%
#17940000000
0!
0%
#17945000000
1!
1%
#17950000000
0!
0%
#17955000000
1!
1%
#17960000000
0!
0%
#17965000000
1!
1%
#17970000000
0!
0%
#17975000000
1!
1%
#17980000000
0!
0%
#17985000000
1!
1%
#17990000000
0!
0%
#17995000000
1!
1%
#18000000000
0!
0%
#18005000000
1!
1%
#18010000000
0!
0%
#18015000000
1!
1%
#18020000000
0!
0%
#18025000000
1!
1%
#18030000000
0!
0%
#18035000000
1!
1%
#18040000000
0!
0%
#18045000000
1!
1%
#18050000000
0!
0%
#18055000000
1!
1%
#18060000000
0!
0%
#18065000000
1!
1%
#18070000000
0!
0%
#18075000000
1!
1%
#18080000000
0!
0%
#18085000000
1!
1%
#18090000000
0!
0%
#18095000000
1!
1%
#18100000000
0!
0%
#18105000000
1!
1%
#18110000000
0!
0%
#18115000000
1!
1%
#18120000000
0!
0%
#18125000000
1!
1%
#18130000000
0!
0%
#18135000000
1!
1%
#18140000000
0!
0%
#18145000000
1!
1%
#18150000000
0!
0%
#18155000000
1!
1%
#18160000000
0!
0%
#18165000000
1!
1%
#18170000000
0!
0%
#18175000000
1!
1%
#18180000000
0!
0%
#18185000000
1!
1%
#18190000000
0!
0%
#18195000000
1!
1%
#18200000000
0!
0%
#18205000000
1!
1%
#18210000000
0!
0%
#18215000000
1!
1%
#18220000000
0!
0%
#18225000000
1!
1%
#18230000000
0!
0%
#18235000000
1!
1%
#18240000000
0!
0%
#18245000000
1!
1%
#18250000000
0!
0%
#18255000000
1!
1%
#18260000000
0!
0%
#18265000000
1!
1%
#18270000000
0!
0%
#18275000000
1!
1%
#18280000000
0!
0%
#18285000000
1!
1%
#18290000000
0!
0%
#18295000000
1!
1%
#18300000000
0!
0%
#18305000000
1!
1%
#18310000000
0!
0%
#18315000000
1!
1%
#18320000000
0!
0%
#18325000000
1!
1%
#18330000000
0!
0%
#18335000000
1!
1%
#18340000000
0!
0%
#18345000000
1!
1%
#18350000000
0!
0%
#18355000000
1!
1%
#18360000000
0!
0%
#18365000000
1!
1%
#18370000000
0!
0%
#18375000000
1!
1%
#18380000000
0!
0%
#18385000000
1!
1%
#18390000000
0!
0%
#18395000000
1!
1%
#18400000000
0!
0%
#18405000000
1!
1%
#18410000000
0!
0%
#18415000000
1!
1%
#18420000000
0!
0%
#18425000000
1!
1%
#18430000000
0!
0%
#18435000000
1!
1%
#18440000000
0!
0%
#18445000000
1!
1%
#18450000000
0!
0%
#18455000000
1!
1%
#18460000000
0!
0%
#18465000000
1!
1%
#18470000000
0!
0%
#18475000000
1!
1%
#18480000000
0!
0%
#18485000000
1!
1%
#18490000000
0!
0%
#18495000000
1!
1%
#18500000000
0!
0%
#18505000000
1!
1%
#18510000000
0!
0%
#18515000000
1!
1%
#18520000000
0!
0%
#18525000000
1!
1%
#18530000000
0!
0%
#18535000000
1!
1%
#18540000000
0!
0%
#18545000000
1!
1%
#18550000000
0!
0%
#18555000000
1!
1%
#18560000000
0!
0%
#18565000000
1!
1%
#18570000000
0!
0%
#18575000000
1!
1%
#18580000000
0!
0%
#18585000000
1!
1%
#18590000000
0!
0%
#18595000000
1!
1%
#18600000000
0!
0%
#18605000000
1!
1%
#18610000000
0!
0%
#18615000000
1!
1%
#18620000000
0!
0%
#18625000000
1!
1%
#18630000000
0!
0%
#18635000000
1!
1%
#18640000000
0!
0%
#18645000000
1!
1%
#18650000000
0!
0%
#18655000000
1!
1%
#18660000000
0!
0%
#18665000000
1!
1%
#18670000000
0!
0%
#18675000000
1!
1%
#18680000000
0!
0%
#18685000000
1!
1%
#18690000000
0!
0%
#18695000000
1!
1%
#18700000000
0!
0%
#18705000000
1!
1%
#18710000000
0!
0%
#18715000000
1!
1%
#18720000000
0!
0%
#18725000000
1!
1%
#18730000000
0!
0%
#18735000000
1!
1%
#18740000000
0!
0%
#18745000000
1!
1%
#18750000000
0!
0%
#18755000000
1!
1%
#18760000000
0!
0%
#18765000000
1!
1%
#18770000000
0!
0%
#18775000000
1!
1%
#18780000000
0!
0%
#18785000000
1!
1%
#18790000000
0!
0%
#18795000000
1!
1%
#18800000000
0!
0%
#18805000000
1!
1%
#18810000000
0!
0%
#18815000000
1!
1%
#18820000000
0!
0%
#18825000000
1!
1%
#18830000000
0!
0%
#18835000000
1!
1%
#18840000000
0!
0%
#18845000000
1!
1%
#18850000000
0!
0%
#18855000000
1!
1%
#18860000000
0!
0%
#18865000000
1!
1%
#18870000000
0!
0%
#18875000000
1!
1%
#18880000000
0!
0%
#18885000000
1!
1%
#18890000000
0!
0%
#18895000000
1!
1%
#18900000000
0!
0%
#18905000000
1!
1%
#18910000000
0!
0%
#18915000000
1!
1%
#18920000000
0!
0%
#18925000000
1!
1%
#18930000000
0!
0%
#18935000000
1!
1%
#18940000000
0!
0%
#18945000000
1!
1%
#18950000000
0!
0%
#18955000000
1!
1%
#18960000000
0!
0%
#18965000000
1!
1%
#18970000000
0!
0%
#18975000000
1!
1%
#18980000000
0!
0%
#18985000000
1!
1%
#18990000000
0!
0%
#18995000000
1!
1%
#19000000000
0!
0%
#19005000000
1!
1%
#19010000000
0!
0%
#19015000000
1!
1%
#19020000000
0!
0%
#19025000000
1!
1%
#19030000000
0!
0%
#19035000000
1!
1%
#19040000000
0!
0%
#19045000000
1!
1%
#19050000000
0!
0%
#19055000000
1!
1%
#19060000000
0!
0%
#19065000000
1!
1%
#19070000000
0!
0%
#19075000000
1!
1%
#19080000000
0!
0%
#19085000000
1!
1%
#19090000000
0!
0%
#19095000000
1!
1%
#19100000000
0!
0%
#19105000000
1!
1%
#19110000000
0!
0%
#19115000000
1!
1%
#19120000000
0!
0%
#19125000000
1!
1%
#19130000000
0!
0%
#19135000000
1!
1%
#19140000000
0!
0%
#19145000000
1!
1%
#19150000000
0!
0%
#19155000000
1!
1%
#19160000000
0!
0%
#19165000000
1!
1%
#19170000000
0!
0%
#19175000000
1!
1%
#19180000000
0!
0%
#19185000000
1!
1%
#19190000000
0!
0%
#19195000000
1!
1%
#19200000000
0!
0%
#19205000000
1!
1%
#19210000000
0!
0%
#19215000000
1!
1%
#19220000000
0!
0%
#19225000000
1!
1%
#19230000000
0!
0%
#19235000000
1!
1%
#19240000000
0!
0%
#19245000000
1!
1%
#19250000000
0!
0%
#19255000000
1!
1%
#19260000000
0!
0%
#19265000000
1!
1%
#19270000000
0!
0%
#19275000000
1!
1%
#19280000000
0!
0%
#19285000000
1!
1%
#19290000000
0!
0%
#19295000000
1!
1%
#19300000000
0!
0%
#19305000000
1!
1%
#19310000000
0!
0%
#19315000000
1!
1%
#19320000000
0!
0%
#19325000000
1!
1%
#19330000000
0!
0%
#19335000000
1!
1%
#19340000000
0!
0%
#19345000000
1!
1%
#19350000000
0!
0%
#19355000000
1!
1%
#19360000000
0!
0%
#19365000000
1!
1%
#19370000000
0!
0%
#19375000000
1!
1%
#19380000000
0!
0%
#19385000000
1!
1%
#19390000000
0!
0%
#19395000000
1!
1%
#19400000000
0!
0%
#19405000000
1!
1%
#19410000000
0!
0%
#19415000000
1!
1%
#19420000000
0!
0%
#19425000000
1!
1%
#19430000000
0!
0%
#19435000000
1!
1%
#19440000000
0!
0%
#19445000000
1!
1%
#19450000000
0!
0%
#19455000000
1!
1%
#19460000000
0!
0%
#19465000000
1!
1%
#19470000000
0!
0%
#19475000000
1!
1%
#19480000000
0!
0%
#19485000000
1!
1%
#19490000000
0!
0%
#19495000000
1!
1%
#19500000000
0!
0%
#19505000000
1!
1%
#19510000000
0!
0%
#19515000000
1!
1%
#19520000000
0!
0%
#19525000000
1!
1%
#19530000000
0!
0%
#19535000000
1!
1%
#19540000000
0!
0%
#19545000000
1!
1%
#19550000000
0!
0%
#19555000000
1!
1%
#19560000000
0!
0%
#19565000000
1!
1%
#19570000000
0!
0%
#19575000000
1!
1%
#19580000000
0!
0%
#19585000000
1!
1%
#19590000000
0!
0%
#19595000000
1!
1%
#19600000000
0!
0%
#19605000000
1!
1%
#19610000000
0!
0%
#19615000000
1!
1%
#19620000000
0!
0%
#19625000000
1!
1%
#19630000000
0!
0%
#19635000000
1!
1%
#19640000000
0!
0%
#19645000000
1!
1%
#19650000000
0!
0%
#19655000000
1!
1%
#19660000000
0!
0%
#19665000000
1!
1%
#19670000000
0!
0%
#19675000000
1!
1%
#19680000000
0!
0%
#19685000000
1!
1%
#19690000000
0!
0%
#19695000000
1!
1%
#19700000000
0!
0%
#19705000000
1!
1%
#19710000000
0!
0%
#19715000000
1!
1%
#19720000000
0!
0%
#19725000000
1!
1%
#19730000000
0!
0%
#19735000000
1!
1%
#19740000000
0!
0%
#19745000000
1!
1%
#19750000000
0!
0%
#19755000000
1!
1%
#19760000000
0!
0%
#19765000000
1!
1%
#19770000000
0!
0%
#19775000000
1!
1%
#19780000000
0!
0%
#19785000000
1!
1%
#19790000000
0!
0%
#19795000000
1!
1%
#19800000000
0!
0%
#19805000000
1!
1%
#19810000000
0!
0%
#19815000000
1!
1%
#19820000000
0!
0%
#19825000000
1!
1%
#19830000000
0!
0%
#19835000000
1!
1%
#19840000000
0!
0%
#19845000000
1!
1%
#19850000000
0!
0%
#19855000000
1!
1%
#19860000000
0!
0%
#19865000000
1!
1%
#19870000000
0!
0%
#19875000000
1!
1%
#19880000000
0!
0%
#19885000000
1!
1%
#19890000000
0!
0%
#19895000000
1!
1%
#19900000000
0!
0%
#19905000000
1!
1%
#19910000000
0!
0%
#19915000000
1!
1%
#19920000000
0!
0%
#19925000000
1!
1%
#19930000000
0!
0%
#19935000000
1!
1%
#19940000000
0!
0%
#19945000000
1!
1%
#19950000000
0!
0%
#19955000000
1!
1%
#19960000000
0!
0%
#19965000000
1!
1%
#19970000000
0!
0%
#19975000000
1!
1%
#19980000000
0!
0%
#19985000000
1!
1%
#19990000000
0!
0%
#19995000000
1!
1%
#20000000000
0!
0%
#20005000000
1!
1%
#20010000000
0!
0%
#20015000000
1!
1%
#20020000000
0!
0%
#20025000000
1!
1%
#20030000000
0!
0%
#20035000000
1!
1%
#20040000000
0!
0%
#20045000000
1!
1%
#20050000000
0!
0%
#20055000000
1!
1%
#20060000000
0!
0%
#20065000000
1!
1%
#20070000000
0!
0%
#20075000000
1!
1%
#20080000000
0!
0%
#20085000000
1!
1%
#20090000000
0!
0%
#20095000000
1!
1%
#20100000000
0!
0%
#20105000000
1!
1%
#20110000000
0!
0%
#20115000000
1!
1%
#20120000000
0!
0%
#20125000000
1!
1%
#20130000000
0!
0%
#20135000000
1!
1%
#20140000000
0!
0%
#20145000000
1!
1%
#20150000000
0!
0%
#20155000000
1!
1%
#20160000000
0!
0%
#20165000000
1!
1%
#20170000000
0!
0%
#20175000000
1!
1%
#20180000000
0!
0%
#20185000000
1!
1%
#20190000000
0!
0%
#20195000000
1!
1%
#20200000000
0!
0%
#20205000000
1!
1%
#20210000000
0!
0%
#20215000000
1!
1%
#20220000000
0!
0%
#20225000000
1!
1%
#20230000000
0!
0%
#20235000000
1!
1%
#20240000000
0!
0%
#20245000000
1!
1%
#20250000000
0!
0%
#20255000000
1!
1%
#20260000000
0!
0%
#20265000000
1!
1%
#20270000000
0!
0%
#20275000000
1!
1%
#20280000000
0!
0%
#20285000000
1!
1%
#20290000000
0!
0%
#20295000000
1!
1%
#20300000000
0!
0%
#20305000000
1!
1%
#20310000000
0!
0%
#20315000000
1!
1%
#20320000000
0!
0%
#20325000000
1!
1%
#20330000000
0!
0%
#20335000000
1!
1%
#20340000000
0!
0%
#20345000000
1!
1%
#20350000000
0!
0%
#20355000000
1!
1%
#20360000000
0!
0%
#20365000000
1!
1%
#20370000000
0!
0%
#20375000000
1!
1%
#20380000000
0!
0%
#20385000000
1!
1%
#20390000000
0!
0%
#20395000000
1!
1%
#20400000000
0!
0%
#20405000000
1!
1%
#20410000000
0!
0%
#20415000000
1!
1%
#20420000000
0!
0%
#20425000000
1!
1%
#20430000000
0!
0%
#20435000000
1!
1%
#20440000000
0!
0%
#20445000000
1!
1%
#20450000000
0!
0%
#20455000000
1!
1%
#20460000000
0!
0%
#20465000000
1!
1%
#20470000000
0!
0%
#20475000000
1!
1%
#20480000000
0!
0%
#20485000000
1!
1%
#20490000000
0!
0%
#20495000000
1!
1%
#20500000000
0!
0%
#20505000000
1!
1%
#20510000000
0!
0%
#20515000000
1!
1%
#20520000000
0!
0%
#20525000000
1!
1%
#20530000000
0!
0%
#20535000000
1!
1%
#20540000000
0!
0%
#20545000000
1!
1%
#20550000000
0!
0%
#20555000000
1!
1%
#20560000000
0!
0%
#20565000000
1!
1%
#20570000000
0!
0%
#20575000000
1!
1%
#20580000000
0!
0%
#20585000000
1!
1%
#20590000000
0!
0%
#20595000000
1!
1%
#20600000000
0!
0%
#20605000000
1!
1%
#20610000000
0!
0%
#20615000000
1!
1%
#20620000000
0!
0%
#20625000000
1!
1%
#20630000000
0!
0%
#20635000000
1!
1%
#20640000000
0!
0%
#20645000000
1!
1%
#20650000000
0!
0%
#20655000000
1!
1%
#20660000000
0!
0%
#20665000000
1!
1%
#20670000000
0!
0%
#20675000000
1!
1%
#20680000000
0!
0%
#20685000000
1!
1%
#20690000000
0!
0%
#20695000000
1!
1%
#20700000000
0!
0%
#20705000000
1!
1%
#20710000000
0!
0%
#20715000000
1!
1%
#20720000000
0!
0%
#20725000000
1!
1%
#20730000000
0!
0%
#20735000000
1!
1%
#20740000000
0!
0%
#20745000000
1!
1%
#20750000000
0!
0%
#20755000000
1!
1%
#20760000000
0!
0%
#20765000000
1!
1%
#20770000000
0!
0%
#20775000000
1!
1%
#20780000000
0!
0%
#20785000000
1!
1%
#20790000000
0!
0%
#20795000000
1!
1%
#20800000000
0!
0%
#20805000000
1!
1%
#20810000000
0!
0%
#20815000000
1!
1%
#20820000000
0!
0%
#20825000000
1!
1%
#20830000000
0!
0%
#20835000000
1!
1%
#20840000000
0!
0%
#20845000000
1!
1%
#20850000000
0!
0%
#20855000000
1!
1%
#20860000000
0!
0%
#20865000000
1!
1%
#20870000000
0!
0%
#20875000000
1!
1%
#20880000000
0!
0%
#20885000000
1!
1%
#20890000000
0!
0%
#20895000000
1!
1%
#20900000000
0!
0%
#20905000000
1!
1%
#20910000000
0!
0%
#20915000000
1!
1%
#20920000000
0!
0%
#20925000000
1!
1%
#20930000000
0!
0%
#20935000000
1!
1%
#20940000000
0!
0%
#20945000000
1!
1%
#20950000000
0!
0%
#20955000000
1!
1%
#20960000000
0!
0%
#20965000000
1!
1%
#20970000000
0!
0%
#20975000000
1!
1%
#20980000000
0!
0%
#20985000000
1!
1%
#20990000000
0!
0%
#20995000000
1!
1%
#21000000000
0!
0%
#21005000000
1!
1%
#21010000000
0!
0%
#21015000000
1!
1%
#21020000000
0!
0%
#21025000000
1!
1%
#21030000000
0!
0%
#21035000000
1!
1%
#21040000000
0!
0%
#21045000000
1!
1%
#21050000000
0!
0%
#21055000000
1!
1%
#21060000000
0!
0%
#21065000000
1!
1%
#21070000000
0!
0%
#21075000000
1!
1%
#21080000000
0!
0%
#21085000000
1!
1%
#21090000000
0!
0%
#21095000000
1!
1%
#21100000000
0!
0%
#21105000000
1!
1%
#21110000000
0!
0%
#21115000000
1!
1%
#21120000000
0!
0%
#21125000000
1!
1%
#21130000000
0!
0%
#21135000000
1!
1%
#21140000000
0!
0%
#21145000000
1!
1%
#21150000000
0!
0%
#21155000000
1!
1%
#21160000000
0!
0%
#21165000000
1!
1%
#21170000000
0!
0%
#21175000000
1!
1%
#21180000000
0!
0%
#21185000000
1!
1%
#21190000000
0!
0%
#21195000000
1!
1%
#21200000000
0!
0%
#21205000000
1!
1%
#21210000000
0!
0%
#21215000000
1!
1%
#21220000000
0!
0%
#21225000000
1!
1%
#21230000000
0!
0%
#21235000000
1!
1%
#21240000000
0!
0%
#21245000000
1!
1%
#21250000000
0!
0%
#21255000000
1!
1%
#21260000000
0!
0%
#21265000000
1!
1%
#21270000000
0!
0%
#21275000000
1!
1%
#21280000000
0!
0%
#21285000000
1!
1%
#21290000000
0!
0%
#21295000000
1!
1%
#21300000000
0!
0%
#21305000000
1!
1%
#21310000000
0!
0%
#21315000000
1!
1%
#21320000000
0!
0%
#21325000000
1!
1%
#21330000000
0!
0%
#21335000000
1!
1%
#21340000000
0!
0%
#21345000000
1!
1%
#21350000000
0!
0%
#21355000000
1!
1%
#21360000000
0!
0%
#21365000000
1!
1%
#21370000000
0!
0%
#21375000000
1!
1%
#21380000000
0!
0%
#21385000000
1!
1%
#21390000000
0!
0%
#21395000000
1!
1%
#21400000000
0!
0%
#21405000000
1!
1%
#21410000000
0!
0%
#21415000000
1!
1%
#21420000000
0!
0%
#21425000000
1!
1%
#21430000000
0!
0%
#21435000000
1!
1%
#21440000000
0!
0%
#21445000000
1!
1%
#21450000000
0!
0%
#21455000000
1!
1%
#21460000000
0!
0%
#21465000000
1!
1%
#21470000000
0!
0%
#21475000000
1!
1%
#21480000000
0!
0%
#21485000000
1!
1%
#21490000000
0!
0%
#21495000000
1!
1%
#21500000000
0!
0%
#21505000000
1!
1%
#21510000000
0!
0%
#21515000000
1!
1%
#21520000000
0!
0%
#21525000000
1!
1%
#21530000000
0!
0%
#21535000000
1!
1%
#21540000000
0!
0%
#21545000000
1!
1%
#21550000000
0!
0%
#21555000000
1!
1%
#21560000000
0!
0%
#21565000000
1!
1%
#21570000000
0!
0%
#21575000000
1!
1%
#21580000000
0!
0%
#21585000000
1!
1%
#21590000000
0!
0%
#21595000000
1!
1%
#21600000000
0!
0%
#21605000000
1!
1%
#21610000000
0!
0%
#21615000000
1!
1%
#21620000000
0!
0%
#21625000000
1!
1%
#21630000000
0!
0%
#21635000000
1!
1%
#21640000000
0!
0%
#21645000000
1!
1%
#21650000000
0!
0%
#21655000000
1!
1%
#21660000000
0!
0%
#21665000000
1!
1%
#21670000000
0!
0%
#21675000000
1!
1%
#21680000000
0!
0%
#21685000000
1!
1%
#21690000000
0!
0%
#21695000000
1!
1%
#21700000000
0!
0%
#21705000000
1!
1%
#21710000000
0!
0%
#21715000000
1!
1%
#21720000000
0!
0%
#21725000000
1!
1%
#21730000000
0!
0%
#21735000000
1!
1%
#21740000000
0!
0%
#21745000000
1!
1%
#21750000000
0!
0%
#21755000000
1!
1%
#21760000000
0!
0%
#21765000000
1!
1%
#21770000000
0!
0%
#21775000000
1!
1%
#21780000000
0!
0%
#21785000000
1!
1%
#21790000000
0!
0%
#21795000000
1!
1%
#21800000000
0!
0%
#21805000000
1!
1%
#21810000000
0!
0%
#21815000000
1!
1%
#21820000000
0!
0%
#21825000000
1!
1%
#21830000000
0!
0%
#21835000000
1!
1%
#21840000000
0!
0%
#21845000000
1!
1%
#21850000000
0!
0%
#21855000000
1!
1%
#21860000000
0!
0%
#21865000000
1!
1%
#21870000000
0!
0%
#21875000000
1!
1%
#21880000000
0!
0%
#21885000000
1!
1%
#21890000000
0!
0%
#21895000000
1!
1%
#21900000000
0!
0%
#21905000000
1!
1%
#21910000000
0!
0%
#21915000000
1!
1%
#21920000000
0!
0%
#21925000000
1!
1%
#21930000000
0!
0%
#21935000000
1!
1%
#21940000000
0!
0%
#21945000000
1!
1%
#21950000000
0!
0%
#21955000000
1!
1%
#21960000000
0!
0%
#21965000000
1!
1%
#21970000000
0!
0%
#21975000000
1!
1%
#21980000000
0!
0%
#21985000000
1!
1%
#21990000000
0!
0%
#21995000000
1!
1%
#22000000000
0!
0%
#22005000000
1!
1%
#22010000000
0!
0%
#22015000000
1!
1%
#22020000000
0!
0%
#22025000000
1!
1%
#22030000000
0!
0%
#22035000000
1!
1%
#22040000000
0!
0%
#22045000000
1!
1%
#22050000000
0!
0%
#22055000000
1!
1%
#22060000000
0!
0%
#22065000000
1!
1%
#22070000000
0!
0%
#22075000000
1!
1%
#22080000000
0!
0%
#22085000000
1!
1%
#22090000000
0!
0%
#22095000000
1!
1%
#22100000000
0!
0%
#22105000000
1!
1%
#22110000000
0!
0%
#22115000000
1!
1%
#22120000000
0!
0%
#22125000000
1!
1%
#22130000000
0!
0%
#22135000000
1!
1%
#22140000000
0!
0%
#22145000000
1!
1%
#22150000000
0!
0%
#22155000000
1!
1%
#22160000000
0!
0%
#22165000000
1!
1%
#22170000000
0!
0%
#22175000000
1!
1%
#22180000000
0!
0%
#22185000000
1!
1%
#22190000000
0!
0%
#22195000000
1!
1%
#22200000000
0!
0%
#22205000000
1!
1%
#22210000000
0!
0%
#22215000000
1!
1%
#22220000000
0!
0%
#22225000000
1!
1%
#22230000000
0!
0%
#22235000000
1!
1%
#22240000000
0!
0%
#22245000000
1!
1%
#22250000000
0!
0%
#22255000000
1!
1%
#22260000000
0!
0%
#22265000000
1!
1%
#22270000000
0!
0%
#22275000000
1!
1%
#22280000000
0!
0%
#22285000000
1!
1%
#22290000000
0!
0%
#22295000000
1!
1%
#22300000000
0!
0%
#22305000000
1!
1%
#22310000000
0!
0%
#22315000000
1!
1%
#22320000000
0!
0%
#22325000000
1!
1%
#22330000000
0!
0%
#22335000000
1!
1%
#22340000000
0!
0%
#22345000000
1!
1%
#22350000000
0!
0%
#22355000000
1!
1%
#22360000000
0!
0%
#22365000000
1!
1%
#22370000000
0!
0%
#22375000000
1!
1%
#22380000000
0!
0%
#22385000000
1!
1%
#22390000000
0!
0%
#22395000000
1!
1%
#22400000000
0!
0%
#22405000000
1!
1%
#22410000000
0!
0%
#22415000000
1!
1%
#22420000000
0!
0%
#22425000000
1!
1%
#22430000000
0!
0%
#22435000000
1!
1%
#22440000000
0!
0%
#22445000000
1!
1%
#22450000000
0!
0%
#22455000000
1!
1%
#22460000000
0!
0%
#22465000000
1!
1%
#22470000000
0!
0%
#22475000000
1!
1%
#22480000000
0!
0%
#22485000000
1!
1%
#22490000000
0!
0%
#22495000000
1!
1%
#22500000000
0!
0%
#22505000000
1!
1%
#22510000000
0!
0%
#22515000000
1!
1%
#22520000000
0!
0%
#22525000000
1!
1%
#22530000000
0!
0%
#22535000000
1!
1%
#22540000000
0!
0%
#22545000000
1!
1%
#22550000000
0!
0%
#22555000000
1!
1%
#22560000000
0!
0%
#22565000000
1!
1%
#22570000000
0!
0%
#22575000000
1!
1%
#22580000000
0!
0%
#22585000000
1!
1%
#22590000000
0!
0%
#22595000000
1!
1%
#22600000000
0!
0%
#22605000000
1!
1%
#22610000000
0!
0%
#22615000000
1!
1%
#22620000000
0!
0%
#22625000000
1!
1%
#22630000000
0!
0%
#22635000000
1!
1%
#22640000000
0!
0%
#22645000000
1!
1%
#22650000000
0!
0%
#22655000000
1!
1%
#22660000000
0!
0%
#22665000000
1!
1%
#22670000000
0!
0%
#22675000000
1!
1%
#22680000000
0!
0%
#22685000000
1!
1%
#22690000000
0!
0%
#22695000000
1!
1%
#22700000000
0!
0%
#22705000000
1!
1%
#22710000000
0!
0%
#22715000000
1!
1%
#22720000000
0!
0%
#22725000000
1!
1%
#22730000000
0!
0%
#22735000000
1!
1%
#22740000000
0!
0%
#22745000000
1!
1%
#22750000000
0!
0%
#22755000000
1!
1%
#22760000000
0!
0%
#22765000000
1!
1%
#22770000000
0!
0%
#22775000000
1!
1%
#22780000000
0!
0%
#22785000000
1!
1%
#22790000000
0!
0%
#22795000000
1!
1%
#22800000000
0!
0%
#22805000000
1!
1%
#22810000000
0!
0%
#22815000000
1!
1%
#22820000000
0!
0%
#22825000000
1!
1%
#22830000000
0!
0%
#22835000000
1!
1%
#22840000000
0!
0%
#22845000000
1!
1%
#22850000000
0!
0%
#22855000000
1!
1%
#22860000000
0!
0%
#22865000000
1!
1%
#22870000000
0!
0%
#22875000000
1!
1%
#22880000000
0!
0%
#22885000000
1!
1%
#22890000000
0!
0%
#22895000000
1!
1%
#22900000000
0!
0%
#22905000000
1!
1%
#22910000000
0!
0%
#22915000000
1!
1%
#22920000000
0!
0%
#22925000000
1!
1%
#22930000000
0!
0%
#22935000000
1!
1%
#22940000000
0!
0%
#22945000000
1!
1%
#22950000000
0!
0%
#22955000000
1!
1%
#22960000000
0!
0%
#22965000000
1!
1%
#22970000000
0!
0%
#22975000000
1!
1%
#22980000000
0!
0%
#22985000000
1!
1%
#22990000000
0!
0%
#22995000000
1!
1%
#23000000000
0!
0%
#23005000000
1!
1%
#23010000000
0!
0%
#23015000000
1!
1%
#23020000000
0!
0%
#23025000000
1!
1%
#23030000000
0!
0%
#23035000000
1!
1%
#23040000000
0!
0%
#23045000000
1!
1%
#23050000000
0!
0%
#23055000000
1!
1%
#23060000000
0!
0%
#23065000000
1!
1%
#23070000000
0!
0%
#23075000000
1!
1%
#23080000000
0!
0%
#23085000000
1!
1%
#23090000000
0!
0%
#23095000000
1!
1%
#23100000000
0!
0%
#23105000000
1!
1%
#23110000000
0!
0%
#23115000000
1!
1%
#23120000000
0!
0%
#23125000000
1!
1%
#23130000000
0!
0%
#23135000000
1!
1%
#23140000000
0!
0%
#23145000000
1!
1%
#23150000000
0!
0%
#23155000000
1!
1%
#23160000000
0!
0%
#23165000000
1!
1%
#23170000000
0!
0%
#23175000000
1!
1%
#23180000000
0!
0%
#23185000000
1!
1%
#23190000000
0!
0%
#23195000000
1!
1%
#23200000000
0!
0%
#23205000000
1!
1%
#23210000000
0!
0%
#23215000000
1!
1%
#23220000000
0!
0%
#23225000000
1!
1%
#23230000000
0!
0%
#23235000000
1!
1%
#23240000000
0!
0%
#23245000000
1!
1%
#23250000000
0!
0%
#23255000000
1!
1%
#23260000000
0!
0%
#23265000000
1!
1%
#23270000000
0!
0%
#23275000000
1!
1%
#23280000000
0!
0%
#23285000000
1!
1%
#23290000000
0!
0%
#23295000000
1!
1%
#23300000000
0!
0%
#23305000000
1!
1%
#23310000000
0!
0%
#23315000000
1!
1%
#23320000000
0!
0%
#23325000000
1!
1%
#23330000000
0!
0%
#23335000000
1!
1%
#23340000000
0!
0%
#23345000000
1!
1%
#23350000000
0!
0%
#23355000000
1!
1%
#23360000000
0!
0%
#23365000000
1!
1%
#23370000000
0!
0%
#23375000000
1!
1%
#23380000000
0!
0%
#23385000000
1!
1%
#23390000000
0!
0%
#23395000000
1!
1%
#23400000000
0!
0%
#23405000000
1!
1%
#23410000000
0!
0%
#23415000000
1!
1%
#23420000000
0!
0%
#23425000000
1!
1%
#23430000000
0!
0%
#23435000000
1!
1%
#23440000000
0!
0%
#23445000000
1!
1%
#23450000000
0!
0%
#23455000000
1!
1%
#23460000000
0!
0%
#23465000000
1!
1%
#23470000000
0!
0%
#23475000000
1!
1%
#23480000000
0!
0%
#23485000000
1!
1%
#23490000000
0!
0%
#23495000000
1!
1%
#23500000000
0!
0%
#23505000000
1!
1%
#23510000000
0!
0%
#23515000000
1!
1%
#23520000000
0!
0%
#23525000000
1!
1%
#23530000000
0!
0%
#23535000000
1!
1%
#23540000000
0!
0%
#23545000000
1!
1%
#23550000000
0!
0%
#23555000000
1!
1%
#23560000000
0!
0%
#23565000000
1!
1%
#23570000000
0!
0%
#23575000000
1!
1%
#23580000000
0!
0%
#23585000000
1!
1%
#23590000000
0!
0%
#23595000000
1!
1%
#23600000000
0!
0%
#23605000000
1!
1%
#23610000000
0!
0%
#23615000000
1!
1%
#23620000000
0!
0%
#23625000000
1!
1%
#23630000000
0!
0%
#23635000000
1!
1%
#23640000000
0!
0%
#23645000000
1!
1%
#23650000000
0!
0%
#23655000000
1!
1%
#23660000000
0!
0%
#23665000000
1!
1%
#23670000000
0!
0%
#23675000000
1!
1%
#23680000000
0!
0%
#23685000000
1!
1%
#23690000000
0!
0%
#23695000000
1!
1%
#23700000000
0!
0%
#23705000000
1!
1%
#23710000000
0!
0%
#23715000000
1!
1%
#23720000000
0!
0%
#23725000000
1!
1%
#23730000000
0!
0%
#23735000000
1!
1%
#23740000000
0!
0%
#23745000000
1!
1%
#23750000000
0!
0%
#23755000000
1!
1%
#23760000000
0!
0%
#23765000000
1!
1%
#23770000000
0!
0%
#23775000000
1!
1%
#23780000000
0!
0%
#23785000000
1!
1%
#23790000000
0!
0%
#23795000000
1!
1%
#23800000000
0!
0%
#23805000000
1!
1%
#23810000000
0!
0%
#23815000000
1!
1%
#23820000000
0!
0%
#23825000000
1!
1%
#23830000000
0!
0%
#23835000000
1!
1%
#23840000000
0!
0%
#23845000000
1!
1%
#23850000000
0!
0%
#23855000000
1!
1%
#23860000000
0!
0%
#23865000000
1!
1%
#23870000000
0!
0%
#23875000000
1!
1%
#23880000000
0!
0%
#23885000000
1!
1%
#23890000000
0!
0%
#23895000000
1!
1%
#23900000000
0!
0%
#23905000000
1!
1%
#23910000000
0!
0%
#23915000000
1!
1%
#23920000000
0!
0%
#23925000000
1!
1%
#23930000000
0!
0%
#23935000000
1!
1%
#23940000000
0!
0%
#23945000000
1!
1%
#23950000000
0!
0%
#23955000000
1!
1%
#23960000000
0!
0%
#23965000000
1!
1%
#23970000000
0!
0%
#23975000000
1!
1%
#23980000000
0!
0%
#23985000000
1!
1%
#23990000000
0!
0%
#23995000000
1!
1%
#24000000000
0!
0%
#24005000000
1!
1%
#24010000000
0!
0%
#24015000000
1!
1%
#24020000000
0!
0%
#24025000000
1!
1%
#24030000000
0!
0%
#24035000000
1!
1%
#24040000000
0!
0%
#24045000000
1!
1%
#24050000000
0!
0%
#24055000000
1!
1%
#24060000000
0!
0%
#24065000000
1!
1%
#24070000000
0!
0%
#24075000000
1!
1%
#24080000000
0!
0%
#24085000000
1!
1%
#24090000000
0!
0%
#24095000000
1!
1%
#24100000000
0!
0%
#24105000000
1!
1%
#24110000000
0!
0%
#24115000000
1!
1%
#24120000000
0!
0%
#24125000000
1!
1%
#24130000000
0!
0%
#24135000000
1!
1%
#24140000000
0!
0%
#24145000000
1!
1%
#24150000000
0!
0%
#24155000000
1!
1%
#24160000000
0!
0%
#24165000000
1!
1%
#24170000000
0!
0%
#24175000000
1!
1%
#24180000000
0!
0%
#24185000000
1!
1%
#24190000000
0!
0%
#24195000000
1!
1%
#24200000000
0!
0%
#24205000000
1!
1%
#24210000000
0!
0%
#24215000000
1!
1%
#24220000000
0!
0%
#24225000000
1!
1%
#24230000000
0!
0%
#24235000000
1!
1%
#24240000000
0!
0%
#24245000000
1!
1%
#24250000000
0!
0%
#24255000000
1!
1%
#24260000000
0!
0%
#24265000000
1!
1%
#24270000000
0!
0%
#24275000000
1!
1%
#24280000000
0!
0%
#24285000000
1!
1%
#24290000000
0!
0%
#24295000000
1!
1%
#24300000000
0!
0%
#24305000000
1!
1%
#24310000000
0!
0%
#24315000000
1!
1%
#24320000000
0!
0%
#24325000000
1!
1%
#24330000000
0!
0%
#24335000000
1!
1%
#24340000000
0!
0%
#24345000000
1!
1%
#24350000000
0!
0%
#24355000000
1!
1%
#24360000000
0!
0%
#24365000000
1!
1%
#24370000000
0!
0%
#24375000000
1!
1%
#24380000000
0!
0%
#24385000000
1!
1%
#24390000000
0!
0%
#24395000000
1!
1%
#24400000000
0!
0%
#24405000000
1!
1%
#24410000000
0!
0%
#24415000000
1!
1%
#24420000000
0!
0%
#24425000000
1!
1%
#24430000000
0!
0%
#24435000000
1!
1%
#24440000000
0!
0%
#24445000000
1!
1%
#24450000000
0!
0%
#24455000000
1!
1%
#24460000000
0!
0%
#24465000000
1!
1%
#24470000000
0!
0%
#24475000000
1!
1%
#24480000000
0!
0%
#24485000000
1!
1%
#24490000000
0!
0%
#24495000000
1!
1%
#24500000000
0!
0%
#24505000000
1!
1%
#24510000000
0!
0%
#24515000000
1!
1%
#24520000000
0!
0%
#24525000000
1!
1%
#24530000000
0!
0%
#24535000000
1!
1%
#24540000000
0!
0%
#24545000000
1!
1%
#24550000000
0!
0%
#24555000000
1!
1%
#24560000000
0!
0%
#24565000000
1!
1%
#24570000000
0!
0%
#24575000000
1!
1%
#24580000000
0!
0%
#24585000000
1!
1%
#24590000000
0!
0%
#24595000000
1!
1%
#24600000000
0!
0%
#24605000000
1!
1%
#24610000000
0!
0%
#24615000000
1!
1%
#24620000000
0!
0%
#24625000000
1!
1%
#24630000000
0!
0%
#24635000000
1!
1%
#24640000000
0!
0%
#24645000000
1!
1%
#24650000000
0!
0%
#24655000000
1!
1%
#24660000000
0!
0%
#24665000000
1!
1%
#24670000000
0!
0%
#24675000000
1!
1%
#24680000000
0!
0%
#24685000000
1!
1%
#24690000000
0!
0%
#24695000000
1!
1%
#24700000000
0!
0%
#24705000000
1!
1%
#24710000000
0!
0%
#24715000000
1!
1%
#24720000000
0!
0%
#24725000000
1!
1%
#24730000000
0!
0%
#24735000000
1!
1%
#24740000000
0!
0%
#24745000000
1!
1%
#24750000000
0!
0%
#24755000000
1!
1%
#24760000000
0!
0%
#24765000000
1!
1%
#24770000000
0!
0%
#24775000000
1!
1%
#24780000000
0!
0%
#24785000000
1!
1%
#24790000000
0!
0%
#24795000000
1!
1%
#24800000000
0!
0%
#24805000000
1!
1%
#24810000000
0!
0%
#24815000000
1!
1%
#24820000000
0!
0%
#24825000000
1!
1%
#24830000000
0!
0%
#24835000000
1!
1%
#24840000000
0!
0%
#24845000000
1!
1%
#24850000000
0!
0%
#24855000000
1!
1%
#24860000000
0!
0%
#24865000000
1!
1%
#24870000000
0!
0%
#24875000000
1!
1%
#24880000000
0!
0%
#24885000000
1!
1%
#24890000000
0!
0%
#24895000000
1!
1%
#24900000000
0!
0%
#24905000000
1!
1%
#24910000000
0!
0%
#24915000000
1!
1%
#24920000000
0!
0%
#24925000000
1!
1%
#24930000000
0!
0%
#24935000000
1!
1%
#24940000000
0!
0%
#24945000000
1!
1%
#24950000000
0!
0%
#24955000000
1!
1%
#24960000000
0!
0%
#24965000000
1!
1%
#24970000000
0!
0%
#24975000000
1!
1%
#24980000000
0!
0%
#24985000000
1!
1%
#24990000000
0!
0%
#24995000000
1!
1%
#25000000000
0!
0%
#25005000000
1!
1%
#25010000000
0!
0%
#25015000000
1!
1%
#25020000000
0!
0%
#25025000000
1!
1%
#25030000000
0!
0%
#25035000000
1!
1%
#25040000000
0!
0%
#25045000000
1!
1%
#25050000000
0!
0%
#25055000000
1!
1%
#25060000000
0!
0%
#25065000000
1!
1%
#25070000000
0!
0%
#25075000000
1!
1%
#25080000000
0!
0%
#25085000000
1!
1%
#25090000000
0!
0%
#25095000000
1!
1%
#25100000000
0!
0%
#25105000000
1!
1%
#25110000000
0!
0%
#25115000000
1!
1%
#25120000000
0!
0%
#25125000000
1!
1%
#25130000000
0!
0%
#25135000000
1!
1%
#25140000000
0!
0%
#25145000000
1!
1%
#25150000000
0!
0%
#25155000000
1!
1%
#25160000000
0!
0%
#25165000000
1!
1%
#25170000000
0!
0%
#25175000000
1!
1%
#25180000000
0!
0%
#25185000000
1!
1%
#25190000000
0!
0%
#25195000000
1!
1%
#25200000000
0!
0%
#25205000000
1!
1%
#25210000000
0!
0%
#25215000000
1!
1%
#25220000000
0!
0%
#25225000000
1!
1%
#25230000000
0!
0%
#25235000000
1!
1%
#25240000000
0!
0%
#25245000000
1!
1%
#25250000000
0!
0%
#25255000000
1!
1%
#25260000000
0!
0%
#25265000000
1!
1%
#25270000000
0!
0%
#25275000000
1!
1%
#25280000000
0!
0%
#25285000000
1!
1%
#25290000000
0!
0%
#25295000000
1!
1%
#25300000000
0!
0%
#25305000000
1!
1%
#25310000000
0!
0%
#25315000000
1!
1%
#25320000000
0!
0%
#25325000000
1!
1%
#25330000000
0!
0%
#25335000000
1!
1%
#25340000000
0!
0%
#25345000000
1!
1%
#25350000000
0!
0%
#25355000000
1!
1%
#25360000000
0!
0%
#25365000000
1!
1%
#25370000000
0!
0%
#25375000000
1!
1%
#25380000000
0!
0%
#25385000000
1!
1%
#25390000000
0!
0%
#25395000000
1!
1%
#25400000000
0!
0%
#25405000000
1!
1%
#25410000000
0!
0%
#25415000000
1!
1%
#25420000000
0!
0%
#25425000000
1!
1%
#25430000000
0!
0%
#25435000000
1!
1%
#25440000000
0!
0%
#25445000000
1!
1%
#25450000000
0!
0%
#25455000000
1!
1%
#25460000000
0!
0%
#25465000000
1!
1%
#25470000000
0!
0%
#25475000000
1!
1%
#25480000000
0!
0%
#25485000000
1!
1%
#25490000000
0!
0%
#25495000000
1!
1%
#25500000000
0!
0%
#25505000000
1!
1%
#25510000000
0!
0%
#25515000000
1!
1%
#25520000000
0!
0%
#25525000000
1!
1%
#25530000000
0!
0%
#25535000000
1!
1%
#25540000000
0!
0%
#25545000000
1!
1%
#25550000000
0!
0%
#25555000000
1!
1%
#25560000000
0!
0%
#25565000000
1!
1%
#25570000000
0!
0%
#25575000000
1!
1%
#25580000000
0!
0%
#25585000000
1!
1%
#25590000000
0!
0%
#25595000000
1!
1%
#25600000000
0!
0%
#25605000000
1!
1%
#25610000000
0!
0%
#25615000000
1!
1%
#25620000000
0!
0%
#25625000000
1!
1%
#25630000000
0!
0%
#25635000000
1!
1%
#25640000000
0!
0%
#25645000000
1!
1%
#25650000000
0!
0%
#25655000000
1!
1%
#25660000000
0!
0%
#25665000000
1!
1%
#25670000000
0!
0%
#25675000000
1!
1%
#25680000000
0!
0%
#25685000000
1!
1%
#25690000000
0!
0%
#25695000000
1!
1%
#25700000000
0!
0%
#25705000000
1!
1%
#25710000000
0!
0%
#25715000000
1!
1%
#25720000000
0!
0%
#25725000000
1!
1%
#25730000000
0!
0%
#25735000000
1!
1%
#25740000000
0!
0%
#25745000000
1!
1%
#25750000000
0!
0%
#25755000000
1!
1%
#25760000000
0!
0%
#25765000000
1!
1%
#25770000000
0!
0%
#25775000000
1!
1%
#25780000000
0!
0%
#25785000000
1!
1%
#25790000000
0!
0%
#25795000000
1!
1%
#25800000000
0!
0%
#25805000000
1!
1%
#25810000000
0!
0%
#25815000000
1!
1%
#25820000000
0!
0%
#25825000000
1!
1%
#25830000000
0!
0%
#25835000000
1!
1%
#25840000000
0!
0%
#25845000000
1!
1%
#25850000000
0!
0%
#25855000000
1!
1%
#25860000000
0!
0%
#25865000000
1!
1%
#25870000000
0!
0%
#25875000000
1!
1%
#25880000000
0!
0%
#25885000000
1!
1%
#25890000000
0!
0%
#25895000000
1!
1%
#25900000000
0!
0%
#25905000000
1!
1%
#25910000000
0!
0%
#25915000000
1!
1%
#25920000000
0!
0%
#25925000000
1!
1%
#25930000000
0!
0%
#25935000000
1!
1%
#25940000000
0!
0%
#25945000000
1!
1%
#25950000000
0!
0%
#25955000000
1!
1%
#25960000000
0!
0%
#25965000000
1!
1%
#25970000000
0!
0%
#25975000000
1!
1%
#25980000000
0!
0%
#25985000000
1!
1%
#25990000000
0!
0%
#25995000000
1!
1%
#26000000000
0!
0%
#26005000000
1!
1%
#26010000000
0!
0%
#26015000000
1!
1%
#26020000000
0!
0%
#26025000000
1!
1%
#26030000000
0!
0%
#26035000000
1!
1%
#26040000000
0!
0%
#26045000000
1!
1%
#26050000000
0!
0%
#26055000000
1!
1%
#26060000000
0!
0%
#26065000000
1!
1%
#26070000000
0!
0%
#26075000000
1!
1%
#26080000000
0!
0%
#26085000000
1!
1%
#26090000000
0!
0%
#26095000000
1!
1%
#26100000000
0!
0%
#26105000000
1!
1%
#26110000000
0!
0%
#26115000000
1!
1%
#26120000000
0!
0%
#26125000000
1!
1%
#26130000000
0!
0%
#26135000000
1!
1%
#26140000000
0!
0%
#26145000000
1!
1%
#26150000000
0!
0%
#26155000000
1!
1%
#26160000000
0!
0%
#26165000000
1!
1%
#26170000000
0!
0%
#26175000000
1!
1%
#26180000000
0!
0%
#26185000000
1!
1%
#26190000000
0!
0%
#26195000000
1!
1%
#26200000000
0!
0%
#26205000000
1!
1%
#26210000000
0!
0%
#26215000000
1!
1%
#26220000000
0!
0%
#26225000000
1!
1%
#26230000000
0!
0%
#26235000000
1!
1%
#26240000000
0!
0%
#26245000000
1!
1%
#26250000000
0!
0%
#26255000000
1!
1%
#26260000000
0!
0%
#26265000000
1!
1%
#26270000000
0!
0%
#26275000000
1!
1%
#26280000000
0!
0%
#26285000000
1!
1%
#26290000000
0!
0%
#26295000000
1!
1%
#26300000000
0!
0%
#26305000000
1!
1%
#26310000000
0!
0%
#26315000000
1!
1%
#26320000000
0!
0%
#26325000000
1!
1%
#26330000000
0!
0%
#26335000000
1!
1%
#26340000000
0!
0%
#26345000000
1!
1%
#26350000000
0!
0%
#26355000000
1!
1%
#26360000000
0!
0%
#26365000000
1!
1%
#26370000000
0!
0%
#26375000000
1!
1%
#26380000000
0!
0%
#26385000000
1!
1%
#26390000000
0!
0%
#26395000000
1!
1%
#26400000000
0!
0%
#26405000000
1!
1%
#26410000000
0!
0%
#26415000000
1!
1%
#26420000000
0!
0%
#26425000000
1!
1%
#26430000000
0!
0%
#26435000000
1!
1%
#26440000000
0!
0%
#26445000000
1!
1%
#26450000000
0!
0%
#26455000000
1!
1%
#26460000000
0!
0%
#26465000000
1!
1%
#26470000000
0!
0%
#26475000000
1!
1%
#26480000000
0!
0%
#26485000000
1!
1%
#26490000000
0!
0%
#26495000000
1!
1%
#26500000000
0!
0%
#26505000000
1!
1%
#26510000000
0!
0%
#26515000000
1!
1%
#26520000000
0!
0%
#26525000000
1!
1%
#26530000000
0!
0%
#26535000000
1!
1%
#26540000000
0!
0%
#26545000000
1!
1%
#26550000000
0!
0%
#26555000000
1!
1%
#26560000000
0!
0%
#26565000000
1!
1%
#26570000000
0!
0%
#26575000000
1!
1%
#26580000000
0!
0%
#26585000000
1!
1%
#26590000000
0!
0%
#26595000000
1!
1%
#26600000000
0!
0%
#26605000000
1!
1%
#26610000000
0!
0%
#26615000000
1!
1%
#26620000000
0!
0%
#26625000000
1!
1%
#26630000000
0!
0%
#26635000000
1!
1%
#26640000000
0!
0%
#26645000000
1!
1%
#26650000000
0!
0%
#26655000000
1!
1%
#26660000000
0!
0%
#26665000000
1!
1%
#26670000000
0!
0%
#26675000000
1!
1%
#26680000000
0!
0%
#26685000000
1!
1%
#26690000000
0!
0%
#26695000000
1!
1%
#26700000000
0!
0%
#26705000000
1!
1%
#26710000000
0!
0%
#26715000000
1!
1%
#26720000000
0!
0%
#26725000000
1!
1%
#26730000000
0!
0%
#26735000000
1!
1%
#26740000000
0!
0%
#26745000000
1!
1%
#26750000000
0!
0%
#26755000000
1!
1%
#26760000000
0!
0%
#26765000000
1!
1%
#26770000000
0!
0%
#26775000000
1!
1%
#26780000000
0!
0%
#26785000000
1!
1%
#26790000000
0!
0%
#26795000000
1!
1%
#26800000000
0!
0%
#26805000000
1!
1%
#26810000000
0!
0%
#26815000000
1!
1%
#26820000000
0!
0%
#26825000000
1!
1%
#26830000000
0!
0%
#26835000000
1!
1%
#26840000000
0!
0%
#26845000000
1!
1%
#26850000000
0!
0%
#26855000000
1!
1%
#26860000000
0!
0%
#26865000000
1!
1%
#26870000000
0!
0%
#26875000000
1!
1%
#26880000000
0!
0%
#26885000000
1!
1%
#26890000000
0!
0%
#26895000000
1!
1%
#26900000000
0!
0%
#26905000000
1!
1%
#26910000000
0!
0%
#26915000000
1!
1%
#26920000000
0!
0%
#26925000000
1!
1%
#26930000000
0!
0%
#26935000000
1!
1%
#26940000000
0!
0%
#26945000000
1!
1%
#26950000000
0!
0%
#26955000000
1!
1%
#26960000000
0!
0%
#26965000000
1!
1%
#26970000000
0!
0%
#26975000000
1!
1%
#26980000000
0!
0%
#26985000000
1!
1%
#26990000000
0!
0%
#26995000000
1!
1%
#27000000000
0!
0%
#27005000000
1!
1%
#27010000000
0!
0%
#27015000000
1!
1%
#27020000000
0!
0%
#27025000000
1!
1%
#27030000000
0!
0%
#27035000000
1!
1%
#27040000000
0!
0%
#27045000000
1!
1%
#27050000000
0!
0%
#27055000000
1!
1%
#27060000000
0!
0%
#27065000000
1!
1%
#27070000000
0!
0%
#27075000000
1!
1%
#27080000000
0!
0%
#27085000000
1!
1%
#27090000000
0!
0%
#27095000000
1!
1%
#27100000000
0!
0%
#27105000000
1!
1%
#27110000000
0!
0%
#27115000000
1!
1%
#27120000000
0!
0%
#27125000000
1!
1%
#27130000000
0!
0%
#27135000000
1!
1%
#27140000000
0!
0%
#27145000000
1!
1%
#27150000000
0!
0%
#27155000000
1!
1%
#27160000000
0!
0%
#27165000000
1!
1%
#27170000000
0!
0%
#27175000000
1!
1%
#27180000000
0!
0%
#27185000000
1!
1%
#27190000000
0!
0%
#27195000000
1!
1%
#27200000000
0!
0%
#27205000000
1!
1%
#27210000000
0!
0%
#27215000000
1!
1%
#27220000000
0!
0%
#27225000000
1!
1%
#27230000000
0!
0%
#27235000000
1!
1%
#27240000000
0!
0%
#27245000000
1!
1%
#27250000000
0!
0%
#27255000000
1!
1%
#27260000000
0!
0%
#27265000000
1!
1%
#27270000000
0!
0%
#27275000000
1!
1%
#27280000000
0!
0%
#27285000000
1!
1%
#27290000000
0!
0%
#27295000000
1!
1%
#27300000000
0!
0%
#27305000000
1!
1%
#27310000000
0!
0%
#27315000000
1!
1%
#27320000000
0!
0%
#27325000000
1!
1%
#27330000000
0!
0%
#27335000000
1!
1%
#27340000000
0!
0%
#27345000000
1!
1%
#27350000000
0!
0%
#27355000000
1!
1%
#27360000000
0!
0%
#27365000000
1!
1%
#27370000000
0!
0%
#27375000000
1!
1%
#27380000000
0!
0%
#27385000000
1!
1%
#27390000000
0!
0%
#27395000000
1!
1%
#27400000000
0!
0%
#27405000000
1!
1%
#27410000000
0!
0%
#27415000000
1!
1%
#27420000000
0!
0%
#27425000000
1!
1%
#27430000000
0!
0%
#27435000000
1!
1%
#27440000000
0!
0%
#27445000000
1!
1%
#27450000000
0!
0%
#27455000000
1!
1%
#27460000000
0!
0%
#27465000000
1!
1%
#27470000000
0!
0%
#27475000000
1!
1%
#27480000000
0!
0%
#27485000000
1!
1%
#27490000000
0!
0%
#27495000000
1!
1%
#27500000000
0!
0%
#27505000000
1!
1%
#27510000000
0!
0%
#27515000000
1!
1%
#27520000000
0!
0%
#27525000000
1!
1%
#27530000000
0!
0%
#27535000000
1!
1%
#27540000000
0!
0%
#27545000000
1!
1%
#27550000000
0!
0%
#27555000000
1!
1%
#27560000000
0!
0%
#27565000000
1!
1%
#27570000000
0!
0%
#27575000000
1!
1%
#27580000000
0!
0%
#27585000000
1!
1%
#27590000000
0!
0%
#27595000000
1!
1%
#27600000000
0!
0%
#27605000000
1!
1%
#27610000000
0!
0%
#27615000000
1!
1%
#27620000000
0!
0%
#27625000000
1!
1%
#27630000000
0!
0%
#27635000000
1!
1%
#27640000000
0!
0%
#27645000000
1!
1%
#27650000000
0!
0%
#27655000000
1!
1%
#27660000000
0!
0%
#27665000000
1!
1%
#27670000000
0!
0%
#27675000000
1!
1%
#27680000000
0!
0%
#27685000000
1!
1%
#27690000000
0!
0%
#27695000000
1!
1%
#27700000000
0!
0%
#27705000000
1!
1%
#27710000000
0!
0%
#27715000000
1!
1%
#27720000000
0!
0%
#27725000000
1!
1%
#27730000000
0!
0%
#27735000000
1!
1%
#27740000000
0!
0%
#27745000000
1!
1%
#27750000000
0!
0%
#27755000000
1!
1%
#27760000000
0!
0%
#27765000000
1!
1%
#27770000000
0!
0%
#27775000000
1!
1%
#27780000000
0!
0%
#27785000000
1!
1%
#27790000000
0!
0%
#27795000000
1!
1%
#27800000000
0!
0%
#27805000000
1!
1%
#27810000000
0!
0%
#27815000000
1!
1%
#27820000000
0!
0%
#27825000000
1!
1%
#27830000000
0!
0%
#27835000000
1!
1%
#27840000000
0!
0%
#27845000000
1!
1%
#27850000000
0!
0%
#27855000000
1!
1%
#27860000000
0!
0%
#27865000000
1!
1%
#27870000000
0!
0%
#27875000000
1!
1%
#27880000000
0!
0%
#27885000000
1!
1%
#27890000000
0!
0%
#27895000000
1!
1%
#27900000000
0!
0%
#27905000000
1!
1%
#27910000000
0!
0%
#27915000000
1!
1%
#27920000000
0!
0%
#27925000000
1!
1%
#27930000000
0!
0%
#27935000000
1!
1%
#27940000000
0!
0%
#27945000000
1!
1%
#27950000000
0!
0%
#27955000000
1!
1%
#27960000000
0!
0%
#27965000000
1!
1%
#27970000000
0!
0%
#27975000000
1!
1%
#27980000000
0!
0%
#27985000000
1!
1%
#27990000000
0!
0%
#27995000000
1!
1%
#28000000000
0!
0%
#28005000000
1!
1%
#28010000000
0!
0%
#28015000000
1!
1%
#28020000000
0!
0%
#28025000000
1!
1%
#28030000000
0!
0%
#28035000000
1!
1%
#28040000000
0!
0%
#28045000000
1!
1%
#28050000000
0!
0%
#28055000000
1!
1%
#28060000000
0!
0%
#28065000000
1!
1%
#28070000000
0!
0%
#28075000000
1!
1%
#28080000000
0!
0%
#28085000000
1!
1%
#28090000000
0!
0%
#28095000000
1!
1%
#28100000000
0!
0%
#28105000000
1!
1%
#28110000000
0!
0%
#28115000000
1!
1%
#28120000000
0!
0%
#28125000000
1!
1%
#28130000000
0!
0%
#28135000000
1!
1%
#28140000000
0!
0%
#28145000000
1!
1%
#28150000000
0!
0%
#28155000000
1!
1%
#28160000000
0!
0%
#28165000000
1!
1%
#28170000000
0!
0%
#28175000000
1!
1%
#28180000000
0!
0%
#28185000000
1!
1%
#28190000000
0!
0%
#28195000000
1!
1%
#28200000000
0!
0%
#28205000000
1!
1%
#28210000000
0!
0%
#28215000000
1!
1%
#28220000000
0!
0%
#28225000000
1!
1%
#28230000000
0!
0%
#28235000000
1!
1%
#28240000000
0!
0%
#28245000000
1!
1%
#28250000000
0!
0%
#28255000000
1!
1%
#28260000000
0!
0%
#28265000000
1!
1%
#28270000000
0!
0%
#28275000000
1!
1%
#28280000000
0!
0%
#28285000000
1!
1%
#28290000000
0!
0%
#28295000000
1!
1%
#28300000000
0!
0%
#28305000000
1!
1%
#28310000000
0!
0%
#28315000000
1!
1%
#28320000000
0!
0%
#28325000000
1!
1%
#28330000000
0!
0%
#28335000000
1!
1%
#28340000000
0!
0%
#28345000000
1!
1%
#28350000000
0!
0%
#28355000000
1!
1%
#28360000000
0!
0%
#28365000000
1!
1%
#28370000000
0!
0%
#28375000000
1!
1%
#28380000000
0!
0%
#28385000000
1!
1%
#28390000000
0!
0%
#28395000000
1!
1%
#28400000000
0!
0%
#28405000000
1!
1%
#28410000000
0!
0%
#28415000000
1!
1%
#28420000000
0!
0%
#28425000000
1!
1%
#28430000000
0!
0%
#28435000000
1!
1%
#28440000000
0!
0%
#28445000000
1!
1%
#28450000000
0!
0%
#28455000000
1!
1%
#28460000000
0!
0%
#28465000000
1!
1%
#28470000000
0!
0%
#28475000000
1!
1%
#28480000000
0!
0%
#28485000000
1!
1%
#28490000000
0!
0%
#28495000000
1!
1%
#28500000000
0!
0%
#28505000000
1!
1%
#28510000000
0!
0%
#28515000000
1!
1%
#28520000000
0!
0%
#28525000000
1!
1%
#28530000000
0!
0%
#28535000000
1!
1%
#28540000000
0!
0%
#28545000000
1!
1%
#28550000000
0!
0%
#28555000000
1!
1%
#28560000000
0!
0%
#28565000000
1!
1%
#28570000000
0!
0%
#28575000000
1!
1%
#28580000000
0!
0%
#28585000000
1!
1%
#28590000000
0!
0%
#28595000000
1!
1%
#28600000000
0!
0%
#28605000000
1!
1%
#28610000000
0!
0%
#28615000000
1!
1%
#28620000000
0!
0%
#28625000000
1!
1%
#28630000000
0!
0%
#28635000000
1!
1%
#28640000000
0!
0%
#28645000000
1!
1%
#28650000000
0!
0%
#28655000000
1!
1%
#28660000000
0!
0%
#28665000000
1!
1%
#28670000000
0!
0%
#28675000000
1!
1%
#28680000000
0!
0%
#28685000000
1!
1%
#28690000000
0!
0%
#28695000000
1!
1%
#28700000000
0!
0%
#28705000000
1!
1%
#28710000000
0!
0%
#28715000000
1!
1%
#28720000000
0!
0%
#28725000000
1!
1%
#28730000000
0!
0%
#28735000000
1!
1%
#28740000000
0!
0%
#28745000000
1!
1%
#28750000000
0!
0%
#28755000000
1!
1%
#28760000000
0!
0%
#28765000000
1!
1%
#28770000000
0!
0%
#28775000000
1!
1%
#28780000000
0!
0%
#28785000000
1!
1%
#28790000000
0!
0%
#28795000000
1!
1%
#28800000000
0!
0%
#28805000000
1!
1%
#28810000000
0!
0%
#28815000000
1!
1%
#28820000000
0!
0%
#28825000000
1!
1%
#28830000000
0!
0%
#28835000000
1!
1%
#28840000000
0!
0%
#28845000000
1!
1%
#28850000000
0!
0%
#28855000000
1!
1%
#28860000000
0!
0%
#28865000000
1!
1%
#28870000000
0!
0%
#28875000000
1!
1%
#28880000000
0!
0%
#28885000000
1!
1%
#28890000000
0!
0%
#28895000000
1!
1%
#28900000000
0!
0%
#28905000000
1!
1%
#28910000000
0!
0%
#28915000000
1!
1%
#28920000000
0!
0%
#28925000000
1!
1%
#28930000000
0!
0%
#28935000000
1!
1%
#28940000000
0!
0%
#28945000000
1!
1%
#28950000000
0!
0%
#28955000000
1!
1%
#28960000000
0!
0%
#28965000000
1!
1%
#28970000000
0!
0%
#28975000000
1!
1%
#28980000000
0!
0%
#28985000000
1!
1%
#28990000000
0!
0%
#28995000000
1!
1%
#29000000000
0!
0%
#29005000000
1!
1%
#29010000000
0!
0%
#29015000000
1!
1%
#29020000000
0!
0%
#29025000000
1!
1%
#29030000000
0!
0%
#29035000000
1!
1%
#29040000000
0!
0%
#29045000000
1!
1%
#29050000000
0!
0%
#29055000000
1!
1%
#29060000000
0!
0%
#29065000000
1!
1%
#29070000000
0!
0%
#29075000000
1!
1%
#29080000000
0!
0%
#29085000000
1!
1%
#29090000000
0!
0%
#29095000000
1!
1%
#29100000000
0!
0%
#29105000000
1!
1%
#29110000000
0!
0%
#29115000000
1!
1%
#29120000000
0!
0%
#29125000000
1!
1%
#29130000000
0!
0%
#29135000000
1!
1%
#29140000000
0!
0%
#29145000000
1!
1%
#29150000000
0!
0%
#29155000000
1!
1%
#29160000000
0!
0%
#29165000000
1!
1%
#29170000000
0!
0%
#29175000000
1!
1%
#29180000000
0!
0%
#29185000000
1!
1%
#29190000000
0!
0%
#29195000000
1!
1%
#29200000000
0!
0%
#29205000000
1!
1%
#29210000000
0!
0%
#29215000000
1!
1%
#29220000000
0!
0%
#29225000000
1!
1%
#29230000000
0!
0%
#29235000000
1!
1%
#29240000000
0!
0%
#29245000000
1!
1%
#29250000000
0!
0%
#29255000000
1!
1%
#29260000000
0!
0%
#29265000000
1!
1%
#29270000000
0!
0%
#29275000000
1!
1%
#29280000000
0!
0%
#29285000000
1!
1%
#29290000000
0!
0%
#29295000000
1!
1%
#29300000000
0!
0%
#29305000000
1!
1%
#29310000000
0!
0%
#29315000000
1!
1%
#29320000000
0!
0%
#29325000000
1!
1%
#29330000000
0!
0%
#29335000000
1!
1%
#29340000000
0!
0%
#29345000000
1!
1%
#29350000000
0!
0%
#29355000000
1!
1%
#29360000000
0!
0%
#29365000000
1!
1%
#29370000000
0!
0%
#29375000000
1!
1%
#29380000000
0!
0%
#29385000000
1!
1%
#29390000000
0!
0%
#29395000000
1!
1%
#29400000000
0!
0%
#29405000000
1!
1%
#29410000000
0!
0%
#29415000000
1!
1%
#29420000000
0!
0%
#29425000000
1!
1%
#29430000000
0!
0%
#29435000000
1!
1%
#29440000000
0!
0%
#29445000000
1!
1%
#29450000000
0!
0%
#29455000000
1!
1%
#29460000000
0!
0%
#29465000000
1!
1%
#29470000000
0!
0%
#29475000000
1!
1%
#29480000000
0!
0%
#29485000000
1!
1%
#29490000000
0!
0%
#29495000000
1!
1%
#29500000000
0!
0%
#29505000000
1!
1%
#29510000000
0!
0%
#29515000000
1!
1%
#29520000000
0!
0%
#29525000000
1!
1%
#29530000000
0!
0%
#29535000000
1!
1%
#29540000000
0!
0%
#29545000000
1!
1%
#29550000000
0!
0%
#29555000000
1!
1%
#29560000000
0!
0%
#29565000000
1!
1%
#29570000000
0!
0%
#29575000000
1!
1%
#29580000000
0!
0%
#29585000000
1!
1%
#29590000000
0!
0%
#29595000000
1!
1%
#29600000000
0!
0%
#29605000000
1!
1%
#29610000000
0!
0%
#29615000000
1!
1%
#29620000000
0!
0%
#29625000000
1!
1%
#29630000000
0!
0%
#29635000000
1!
1%
#29640000000
0!
0%
#29645000000
1!
1%
#29650000000
0!
0%
#29655000000
1!
1%
#29660000000
0!
0%
#29665000000
1!
1%
#29670000000
0!
0%
#29675000000
1!
1%
#29680000000
0!
0%
#29685000000
1!
1%
#29690000000
0!
0%
#29695000000
1!
1%
#29700000000
0!
0%
#29705000000
1!
1%
#29710000000
0!
0%
#29715000000
1!
1%
#29720000000
0!
0%
#29725000000
1!
1%
#29730000000
0!
0%
#29735000000
1!
1%
#29740000000
0!
0%
#29745000000
1!
1%
#29750000000
0!
0%
#29755000000
1!
1%
#29760000000
0!
0%
#29765000000
1!
1%
#29770000000
0!
0%
#29775000000
1!
1%
#29780000000
0!
0%
#29785000000
1!
1%
#29790000000
0!
0%
#29795000000
1!
1%
#29800000000
0!
0%
#29805000000
1!
1%
#29810000000
0!
0%
#29815000000
1!
1%
#29820000000
0!
0%
#29825000000
1!
1%
#29830000000
0!
0%
#29835000000
1!
1%
#29840000000
0!
0%
#29845000000
1!
1%
#29850000000
0!
0%
#29855000000
1!
1%
#29860000000
0!
0%
#29865000000
1!
1%
#29870000000
0!
0%
#29875000000
1!
1%
#29880000000
0!
0%
#29885000000
1!
1%
#29890000000
0!
0%
#29895000000
1!
1%
#29900000000
0!
0%
#29905000000
1!
1%
#29910000000
0!
0%
#29915000000
1!
1%
#29920000000
0!
0%
#29925000000
1!
1%
#29930000000
0!
0%
#29935000000
1!
1%
#29940000000
0!
0%
#29945000000
1!
1%
#29950000000
0!
0%
#29955000000
1!
1%
#29960000000
0!
0%
#29965000000
1!
1%
#29970000000
0!
0%
#29975000000
1!
1%
#29980000000
0!
0%
#29985000000
1!
1%
#29990000000
0!
0%
#29995000000
1!
1%
#30000000000
0!
0%
#30005000000
1!
1%
#30010000000
0!
0%
#30015000000
1!
1%
#30020000000
0!
0%
#30025000000
1!
1%
#30030000000
0!
0%
#30035000000
1!
1%
#30040000000
0!
0%
#30045000000
1!
1%
#30050000000
0!
0%
#30055000000
1!
1%
#30060000000
0!
0%
#30065000000
1!
1%
#30070000000
0!
0%
#30075000000
1!
1%
#30080000000
0!
0%
#30085000000
1!
1%
#30090000000
0!
0%
#30095000000
1!
1%
#30100000000
0!
0%
#30105000000
1!
1%
#30110000000
0!
0%
#30115000000
1!
1%
#30120000000
0!
0%
#30125000000
1!
1%
#30130000000
0!
0%
#30135000000
1!
1%
#30140000000
0!
0%
#30145000000
1!
1%
#30150000000
0!
0%
#30155000000
1!
1%
#30160000000
0!
0%
#30165000000
1!
1%
#30170000000
0!
0%
#30175000000
1!
1%
#30180000000
0!
0%
#30185000000
1!
1%
#30190000000
0!
0%
#30195000000
1!
1%
#30200000000
0!
0%
#30205000000
1!
1%
#30210000000
0!
0%
#30215000000
1!
1%
#30220000000
0!
0%
#30225000000
1!
1%
#30230000000
0!
0%
#30235000000
1!
1%
#30240000000
0!
0%
#30245000000
1!
1%
#30250000000
0!
0%
#30255000000
1!
1%
#30260000000
0!
0%
#30265000000
1!
1%
#30270000000
0!
0%
#30275000000
1!
1%
#30280000000
0!
0%
#30285000000
1!
1%
#30290000000
0!
0%
#30295000000
1!
1%
#30300000000
0!
0%
#30305000000
1!
1%
#30310000000
0!
0%
#30315000000
1!
1%
#30320000000
0!
0%
#30325000000
1!
1%
#30330000000
0!
0%
#30335000000
1!
1%
#30340000000
0!
0%
#30345000000
1!
1%
#30350000000
0!
0%
#30355000000
1!
1%
#30360000000
0!
0%
#30365000000
1!
1%
#30370000000
0!
0%
#30375000000
1!
1%
#30380000000
0!
0%
#30385000000
1!
1%
#30390000000
0!
0%
#30395000000
1!
1%
#30400000000
0!
0%
#30405000000
1!
1%
#30410000000
0!
0%
#30415000000
1!
1%
#30420000000
0!
0%
#30425000000
1!
1%
#30430000000
0!
0%
#30435000000
1!
1%
#30440000000
0!
0%
#30445000000
1!
1%
#30450000000
0!
0%
#30455000000
1!
1%
#30460000000
0!
0%
#30465000000
1!
1%
#30470000000
0!
0%
#30475000000
1!
1%
#30480000000
0!
0%
#30485000000
1!
1%
#30490000000
0!
0%
#30495000000
1!
1%
#30500000000
0!
0%
#30505000000
1!
1%
#30510000000
0!
0%
#30515000000
1!
1%
#30520000000
0!
0%
#30525000000
1!
1%
#30530000000
0!
0%
#30535000000
1!
1%
#30540000000
0!
0%
#30545000000
1!
1%
#30550000000
0!
0%
#30555000000
1!
1%
#30560000000
0!
0%
#30565000000
1!
1%
#30570000000
0!
0%
#30575000000
1!
1%
#30580000000
0!
0%
#30585000000
1!
1%
#30590000000
0!
0%
#30595000000
1!
1%
#30600000000
0!
0%
#30605000000
1!
1%
#30610000000
0!
0%
#30615000000
1!
1%
#30620000000
0!
0%
#30625000000
1!
1%
#30630000000
0!
0%
#30635000000
1!
1%
#30640000000
0!
0%
#30645000000
1!
1%
#30650000000
0!
0%
#30655000000
1!
1%
#30660000000
0!
0%
#30665000000
1!
1%
#30670000000
0!
0%
#30675000000
1!
1%
#30680000000
0!
0%
#30685000000
1!
1%
#30690000000
0!
0%
#30695000000
1!
1%
#30700000000
0!
0%
#30705000000
1!
1%
#30710000000
0!
0%
#30715000000
1!
1%
#30720000000
0!
0%
#30725000000
1!
1%
#30730000000
0!
0%
#30735000000
1!
1%
#30740000000
0!
0%
#30745000000
1!
1%
#30750000000
0!
0%
#30755000000
1!
1%
#30760000000
0!
0%
#30765000000
1!
1%
#30770000000
0!
0%
#30775000000
1!
1%
#30780000000
0!
0%
#30785000000
1!
1%
#30790000000
0!
0%
#30795000000
1!
1%
#30800000000
0!
0%
#30805000000
1!
1%
#30810000000
0!
0%
#30815000000
1!
1%
#30820000000
0!
0%
#30825000000
1!
1%
#30830000000
0!
0%
#30835000000
1!
1%
#30840000000
0!
0%
#30845000000
1!
1%
#30850000000
0!
0%
#30855000000
1!
1%
#30860000000
0!
0%
#30865000000
1!
1%
#30870000000
0!
0%
#30875000000
1!
1%
#30880000000
0!
0%
#30885000000
1!
1%
#30890000000
0!
0%
#30895000000
1!
1%
#30900000000
0!
0%
#30905000000
1!
1%
#30910000000
0!
0%
#30915000000
1!
1%
#30920000000
0!
0%
#30925000000
1!
1%
#30930000000
0!
0%
#30935000000
1!
1%
#30940000000
0!
0%
#30945000000
1!
1%
#30950000000
0!
0%
#30955000000
1!
1%
#30960000000
0!
0%
#30965000000
1!
1%
#30970000000
0!
0%
#30975000000
1!
1%
#30980000000
0!
0%
#30985000000
1!
1%
#30990000000
0!
0%
#30995000000
1!
1%
#31000000000
0!
0%
#31005000000
1!
1%
#31010000000
0!
0%
#31015000000
1!
1%
#31020000000
0!
0%
#31025000000
1!
1%
#31030000000
0!
0%
#31035000000
1!
1%
#31040000000
0!
0%
#31045000000
1!
1%
#31050000000
0!
0%
#31055000000
1!
1%
#31060000000
0!
0%
#31065000000
1!
1%
#31070000000
0!
0%
#31075000000
1!
1%
#31080000000
0!
0%
#31085000000
1!
1%
#31090000000
0!
0%
#31095000000
1!
1%
#31100000000
0!
0%
#31105000000
1!
1%
#31110000000
0!
0%
#31115000000
1!
1%
#31120000000
0!
0%
#31125000000
1!
1%
#31130000000
0!
0%
#31135000000
1!
1%
#31140000000
0!
0%
#31145000000
1!
1%
#31150000000
0!
0%
#31155000000
1!
1%
#31160000000
0!
0%
#31165000000
1!
1%
#31170000000
0!
0%
#31175000000
1!
1%
#31180000000
0!
0%
#31185000000
1!
1%
#31190000000
0!
0%
#31195000000
1!
1%
#31200000000
0!
0%
#31205000000
1!
1%
#31210000000
0!
0%
#31215000000
1!
1%
#31220000000
0!
0%
#31225000000
1!
1%
#31230000000
0!
0%
#31235000000
1!
1%
#31240000000
0!
0%
#31245000000
1!
1%
#31250000000
0!
0%
#31255000000
1!
1%
#31260000000
0!
0%
#31265000000
1!
1%
#31270000000
0!
0%
#31275000000
1!
1%
#31280000000
0!
0%
#31285000000
1!
1%
#31290000000
0!
0%
#31295000000
1!
1%
#31300000000
0!
0%
#31305000000
1!
1%
#31310000000
0!
0%
#31315000000
1!
1%
#31320000000
0!
0%
#31325000000
1!
1%
#31330000000
0!
0%
#31335000000
1!
1%
#31340000000
0!
0%
#31345000000
1!
1%
#31350000000
0!
0%
#31355000000
1!
1%
#31360000000
0!
0%
#31365000000
1!
1%
#31370000000
0!
0%
#31375000000
1!
1%
#31380000000
0!
0%
#31385000000
1!
1%
#31390000000
0!
0%
#31395000000
1!
1%
#31400000000
0!
0%
#31405000000
1!
1%
#31410000000
0!
0%
#31415000000
1!
1%
#31420000000
0!
0%
#31425000000
1!
1%
#31430000000
0!
0%
#31435000000
1!
1%
#31440000000
0!
0%
#31445000000
1!
1%
#31450000000
0!
0%
#31455000000
1!
1%
#31460000000
0!
0%
#31465000000
1!
1%
#31470000000
0!
0%
#31475000000
1!
1%
#31480000000
0!
0%
#31485000000
1!
1%
#31490000000
0!
0%
#31495000000
1!
1%
#31500000000
0!
0%
#31505000000
1!
1%
#31510000000
0!
0%
#31515000000
1!
1%
#31520000000
0!
0%
#31525000000
1!
1%
#31530000000
0!
0%
#31535000000
1!
1%
#31540000000
0!
0%
#31545000000
1!
1%
#31550000000
0!
0%
#31555000000
1!
1%
#31560000000
0!
0%
#31565000000
1!
1%
#31570000000
0!
0%
#31575000000
1!
1%
#31580000000
0!
0%
#31585000000
1!
1%
#31590000000
0!
0%
#31595000000
1!
1%
#31600000000
0!
0%
#31605000000
1!
1%
#31610000000
0!
0%
#31615000000
1!
1%
#31620000000
0!
0%
#31625000000
1!
1%
#31630000000
0!
0%
#31635000000
1!
1%
#31640000000
0!
0%
#31645000000
1!
1%
#31650000000
0!
0%
#31655000000
1!
1%
#31660000000
0!
0%
#31665000000
1!
1%
#31670000000
0!
0%
#31675000000
1!
1%
#31680000000
0!
0%
#31685000000
1!
1%
#31690000000
0!
0%
#31695000000
1!
1%
#31700000000
0!
0%
#31705000000
1!
1%
#31710000000
0!
0%
#31715000000
1!
1%
#31720000000
0!
0%
#31725000000
1!
1%
#31730000000
0!
0%
#31735000000
1!
1%
#31740000000
0!
0%
#31745000000
1!
1%
#31750000000
0!
0%
#31755000000
1!
1%
#31760000000
0!
0%
#31765000000
1!
1%
#31770000000
0!
0%
#31775000000
1!
1%
#31780000000
0!
0%
#31785000000
1!
1%
#31790000000
0!
0%
#31795000000
1!
1%
#31800000000
0!
0%
#31805000000
1!
1%
#31810000000
0!
0%
#31815000000
1!
1%
#31820000000
0!
0%
#31825000000
1!
1%
#31830000000
0!
0%
#31835000000
1!
1%
#31840000000
0!
0%
#31845000000
1!
1%
#31850000000
0!
0%
#31855000000
1!
1%
#31860000000
0!
0%
#31865000000
1!
1%
#31870000000
0!
0%
#31875000000
1!
1%
#31880000000
0!
0%
#31885000000
1!
1%
#31890000000
0!
0%
#31895000000
1!
1%
#31900000000
0!
0%
#31905000000
1!
1%
#31910000000
0!
0%
#31915000000
1!
1%
#31920000000
0!
0%
#31925000000
1!
1%
#31930000000
0!
0%
#31935000000
1!
1%
#31940000000
0!
0%
#31945000000
1!
1%
#31950000000
0!
0%
#31955000000
1!
1%
#31960000000
0!
0%
#31965000000
1!
1%
#31970000000
0!
0%
#31975000000
1!
1%
#31980000000
0!
0%
#31985000000
1!
1%
#31990000000
0!
0%
#31995000000
1!
1%
#32000000000
0!
0%
#32005000000
1!
1%
#32010000000
0!
0%
#32015000000
1!
1%
#32020000000
0!
0%
#32025000000
1!
1%
#32030000000
0!
0%
#32035000000
1!
1%
#32040000000
0!
0%
#32045000000
1!
1%
#32050000000
0!
0%
#32055000000
1!
1%
#32060000000
0!
0%
#32065000000
1!
1%
#32070000000
0!
0%
#32075000000
1!
1%
#32080000000
0!
0%
#32085000000
1!
1%
#32090000000
0!
0%
#32095000000
1!
1%
#32100000000
0!
0%
#32105000000
1!
1%
#32110000000
0!
0%
#32115000000
1!
1%
#32120000000
0!
0%
#32125000000
1!
1%
#32130000000
0!
0%
#32135000000
1!
1%
#32140000000
0!
0%
#32145000000
1!
1%
#32150000000
0!
0%
#32155000000
1!
1%
#32160000000
0!
0%
#32165000000
1!
1%
#32170000000
0!
0%
#32175000000
1!
1%
#32180000000
0!
0%
#32185000000
1!
1%
#32190000000
0!
0%
#32195000000
1!
1%
#32200000000
0!
0%
#32205000000
1!
1%
#32210000000
0!
0%
#32215000000
1!
1%
#32220000000
0!
0%
#32225000000
1!
1%
#32230000000
0!
0%
#32235000000
1!
1%
#32240000000
0!
0%
#32245000000
1!
1%
#32250000000
0!
0%
#32255000000
1!
1%
#32260000000
0!
0%
#32265000000
1!
1%
#32270000000
0!
0%
#32275000000
1!
1%
#32280000000
0!
0%
#32285000000
1!
1%
#32290000000
0!
0%
#32295000000
1!
1%
#32300000000
0!
0%
#32305000000
1!
1%
#32310000000
0!
0%
#32315000000
1!
1%
#32320000000
0!
0%
#32325000000
1!
1%
#32330000000
0!
0%
#32335000000
1!
1%
#32340000000
0!
0%
#32345000000
1!
1%
#32350000000
0!
0%
#32355000000
1!
1%
#32360000000
0!
0%
#32365000000
1!
1%
#32370000000
0!
0%
#32375000000
1!
1%
#32380000000
0!
0%
#32385000000
1!
1%
#32390000000
0!
0%
#32395000000
1!
1%
#32400000000
0!
0%
#32405000000
1!
1%
#32410000000
0!
0%
#32415000000
1!
1%
#32420000000
0!
0%
#32425000000
1!
1%
#32430000000
0!
0%
#32435000000
1!
1%
#32440000000
0!
0%
#32445000000
1!
1%
#32450000000
0!
0%
#32455000000
1!
1%
#32460000000
0!
0%
#32465000000
1!
1%
#32470000000
0!
0%
#32475000000
1!
1%
#32480000000
0!
0%
#32485000000
1!
1%
#32490000000
0!
0%
#32495000000
1!
1%
#32500000000
0!
0%
#32505000000
1!
1%
#32510000000
0!
0%
#32515000000
1!
1%
#32520000000
0!
0%
#32525000000
1!
1%
#32530000000
0!
0%
#32535000000
1!
1%
#32540000000
0!
0%
#32545000000
1!
1%
#32550000000
0!
0%
#32555000000
1!
1%
#32560000000
0!
0%
#32565000000
1!
1%
#32570000000
0!
0%
#32575000000
1!
1%
#32580000000
0!
0%
#32585000000
1!
1%
#32590000000
0!
0%
#32595000000
1!
1%
#32600000000
0!
0%
#32605000000
1!
1%
#32610000000
0!
0%
#32615000000
1!
1%
#32620000000
0!
0%
#32625000000
1!
1%
#32630000000
0!
0%
#32635000000
1!
1%
#32640000000
0!
0%
#32645000000
1!
1%
#32650000000
0!
0%
#32655000000
1!
1%
#32660000000
0!
0%
#32665000000
1!
1%
#32670000000
0!
0%
#32675000000
1!
1%
#32680000000
0!
0%
#32685000000
1!
1%
#32690000000
0!
0%
#32695000000
1!
1%
#32700000000
0!
0%
#32705000000
1!
1%
#32710000000
0!
0%
#32715000000
1!
1%
#32720000000
0!
0%
#32725000000
1!
1%
#32730000000
0!
0%
#32735000000
1!
1%
#32740000000
0!
0%
#32745000000
1!
1%
#32750000000
0!
0%
#32755000000
1!
1%
#32760000000
0!
0%
#32765000000
1!
1%
#32770000000
0!
0%
#32775000000
1!
1%
#32780000000
0!
0%
#32785000000
1!
1%
#32790000000
0!
0%
#32795000000
1!
1%
#32800000000
0!
0%
#32805000000
1!
1%
#32810000000
0!
0%
#32815000000
1!
1%
#32820000000
0!
0%
#32825000000
1!
1%
#32830000000
0!
0%
#32835000000
1!
1%
#32840000000
0!
0%
#32845000000
1!
1%
#32850000000
0!
0%
#32855000000
1!
1%
#32860000000
0!
0%
#32865000000
1!
1%
#32870000000
0!
0%
#32875000000
1!
1%
#32880000000
0!
0%
#32885000000
1!
1%
#32890000000
0!
0%
#32895000000
1!
1%
#32900000000
0!
0%
#32905000000
1!
1%
#32910000000
0!
0%
#32915000000
1!
1%
#32920000000
0!
0%
#32925000000
1!
1%
#32930000000
0!
0%
#32935000000
1!
1%
#32940000000
0!
0%
#32945000000
1!
1%
#32950000000
0!
0%
#32955000000
1!
1%
#32960000000
0!
0%
#32965000000
1!
1%
#32970000000
0!
0%
#32975000000
1!
1%
#32980000000
0!
0%
#32985000000
1!
1%
#32990000000
0!
0%
#32995000000
1!
1%
#33000000000
0!
0%
#33005000000
1!
1%
#33010000000
0!
0%
#33015000000
1!
1%
#33020000000
0!
0%
#33025000000
1!
1%
#33030000000
0!
0%
#33035000000
1!
1%
#33040000000
0!
0%
#33045000000
1!
1%
#33050000000
0!
0%
#33055000000
1!
1%
#33060000000
0!
0%
#33065000000
1!
1%
#33070000000
0!
0%
#33075000000
1!
1%
#33080000000
0!
0%
#33085000000
1!
1%
#33090000000
0!
0%
#33095000000
1!
1%
#33100000000
0!
0%
#33105000000
1!
1%
#33110000000
0!
0%
#33115000000
1!
1%
#33120000000
0!
0%
#33125000000
1!
1%
#33130000000
0!
0%
#33135000000
1!
1%
#33140000000
0!
0%
#33145000000
1!
1%
#33150000000
0!
0%
#33155000000
1!
1%
#33160000000
0!
0%
#33165000000
1!
1%
#33170000000
0!
0%
#33175000000
1!
1%
#33180000000
0!
0%
#33185000000
1!
1%
#33190000000
0!
0%
#33195000000
1!
1%
#33200000000
0!
0%
#33205000000
1!
1%
#33210000000
0!
0%
#33215000000
1!
1%
#33220000000
0!
0%
#33225000000
1!
1%
#33230000000
0!
0%
#33235000000
1!
1%
#33240000000
0!
0%
#33245000000
1!
1%
#33250000000
0!
0%
#33255000000
1!
1%
#33260000000
0!
0%
#33265000000
1!
1%
#33270000000
0!
0%
#33275000000
1!
1%
#33280000000
0!
0%
#33285000000
1!
1%
#33290000000
0!
0%
#33295000000
1!
1%
#33300000000
0!
0%
#33305000000
1!
1%
#33310000000
0!
0%
#33315000000
1!
1%
#33320000000
0!
0%
#33325000000
1!
1%
#33330000000
0!
0%
#33335000000
1!
1%
#33340000000
0!
0%
#33345000000
1!
1%
#33350000000
0!
0%
#33355000000
1!
1%
#33360000000
0!
0%
#33365000000
1!
1%
#33370000000
0!
0%
#33375000000
1!
1%
#33380000000
0!
0%
#33385000000
1!
1%
#33390000000
0!
0%
#33395000000
1!
1%
#33400000000
0!
0%
#33405000000
1!
1%
#33410000000
0!
0%
#33415000000
1!
1%
#33420000000
0!
0%
#33425000000
1!
1%
#33430000000
0!
0%
#33435000000
1!
1%
#33440000000
0!
0%
#33445000000
1!
1%
#33450000000
0!
0%
#33455000000
1!
1%
#33460000000
0!
0%
#33465000000
1!
1%
#33470000000
0!
0%
#33475000000
1!
1%
#33480000000
0!
0%
#33485000000
1!
1%
#33490000000
0!
0%
#33495000000
1!
1%
#33500000000
0!
0%
#33505000000
1!
1%
#33510000000
0!
0%
#33515000000
1!
1%
#33520000000
0!
0%
#33525000000
1!
1%
#33530000000
0!
0%
#33535000000
1!
1%
#33540000000
0!
0%
#33545000000
1!
1%
#33550000000
0!
0%
#33555000000
1!
1%
#33560000000
0!
0%
#33565000000
1!
1%
#33570000000
0!
0%
#33575000000
1!
1%
#33580000000
0!
0%
#33585000000
1!
1%
#33590000000
0!
0%
#33595000000
1!
1%
#33600000000
0!
0%
#33605000000
1!
1%
#33610000000
0!
0%
#33615000000
1!
1%
#33620000000
0!
0%
#33625000000
1!
1%
#33630000000
0!
0%
#33635000000
1!
1%
#33640000000
0!
0%
#33645000000
1!
1%
#33650000000
0!
0%
#33655000000
1!
1%
#33660000000
0!
0%
#33665000000
1!
1%
#33670000000
0!
0%
#33675000000
1!
1%
#33680000000
0!
0%
#33685000000
1!
1%
#33690000000
0!
0%
#33695000000
1!
1%
#33700000000
0!
0%
#33705000000
1!
1%
#33710000000
0!
0%
#33715000000
1!
1%
#33720000000
0!
0%
#33725000000
1!
1%
#33730000000
0!
0%
#33735000000
1!
1%
#33740000000
0!
0%
#33745000000
1!
1%
#33750000000
0!
0%
#33755000000
1!
1%
#33760000000
0!
0%
#33765000000
1!
1%
#33770000000
0!
0%
#33775000000
1!
1%
#33780000000
0!
0%
#33785000000
1!
1%
#33790000000
0!
0%
#33795000000
1!
1%
#33800000000
0!
0%
#33805000000
1!
1%
#33810000000
0!
0%
#33815000000
1!
1%
#33820000000
0!
0%
#33825000000
1!
1%
#33830000000
0!
0%
#33835000000
1!
1%
#33840000000
0!
0%
#33845000000
1!
1%
#33850000000
0!
0%
#33855000000
1!
1%
#33860000000
0!
0%
#33865000000
1!
1%
#33870000000
0!
0%
#33875000000
1!
1%
#33880000000
0!
0%
#33885000000
1!
1%
#33890000000
0!
0%
#33895000000
1!
1%
#33900000000
0!
0%
#33905000000
1!
1%
#33910000000
0!
0%
#33915000000
1!
1%
#33920000000
0!
0%
#33925000000
1!
1%
#33930000000
0!
0%
#33935000000
1!
1%
#33940000000
0!
0%
#33945000000
1!
1%
#33950000000
0!
0%
#33955000000
1!
1%
#33960000000
0!
0%
#33965000000
1!
1%
#33970000000
0!
0%
#33975000000
1!
1%
#33980000000
0!
0%
#33985000000
1!
1%
#33990000000
0!
0%
#33995000000
1!
1%
#34000000000
0!
0%
#34005000000
1!
1%
#34010000000
0!
0%
#34015000000
1!
1%
#34020000000
0!
0%
#34025000000
1!
1%
#34030000000
0!
0%
#34035000000
1!
1%
#34040000000
0!
0%
#34045000000
1!
1%
#34050000000
0!
0%
#34055000000
1!
1%
#34060000000
0!
0%
#34065000000
1!
1%
#34070000000
0!
0%
#34075000000
1!
1%
#34080000000
0!
0%
#34085000000
1!
1%
#34090000000
0!
0%
#34095000000
1!
1%
#34100000000
0!
0%
#34105000000
1!
1%
#34110000000
0!
0%
#34115000000
1!
1%
#34120000000
0!
0%
#34125000000
1!
1%
#34130000000
0!
0%
#34135000000
1!
1%
#34140000000
0!
0%
#34145000000
1!
1%
#34150000000
0!
0%
#34155000000
1!
1%
#34160000000
0!
0%
#34165000000
1!
1%
#34170000000
0!
0%
#34175000000
1!
1%
#34180000000
0!
0%
#34185000000
1!
1%
#34190000000
0!
0%
#34195000000
1!
1%
#34200000000
0!
0%
#34205000000
1!
1%
#34210000000
0!
0%
#34215000000
1!
1%
#34220000000
0!
0%
#34225000000
1!
1%
#34230000000
0!
0%
#34235000000
1!
1%
#34240000000
0!
0%
#34245000000
1!
1%
#34250000000
0!
0%
#34255000000
1!
1%
#34260000000
0!
0%
#34265000000
1!
1%
#34270000000
0!
0%
#34275000000
1!
1%
#34280000000
0!
0%
#34285000000
1!
1%
#34290000000
0!
0%
#34295000000
1!
1%
#34300000000
0!
0%
#34305000000
1!
1%
#34310000000
0!
0%
#34315000000
1!
1%
#34320000000
0!
0%
#34325000000
1!
1%
#34330000000
0!
0%
#34335000000
1!
1%
#34340000000
0!
0%
#34345000000
1!
1%
#34350000000
0!
0%
#34355000000
1!
1%
#34360000000
0!
0%
#34365000000
1!
1%
#34370000000
0!
0%
#34375000000
1!
1%
#34380000000
0!
0%
#34385000000
1!
1%
#34390000000
0!
0%
#34395000000
1!
1%
#34400000000
0!
0%
#34405000000
1!
1%
#34410000000
0!
0%
#34415000000
1!
1%
#34420000000
0!
0%
#34425000000
1!
1%
#34430000000
0!
0%
#34435000000
1!
1%
#34440000000
0!
0%
#34445000000
1!
1%
#34450000000
0!
0%
#34455000000
1!
1%
#34460000000
0!
0%
#34465000000
1!
1%
#34470000000
0!
0%
#34475000000
1!
1%
#34480000000
0!
0%
#34485000000
1!
1%
#34490000000
0!
0%
#34495000000
1!
1%
#34500000000
0!
0%
#34505000000
1!
1%
#34510000000
0!
0%
#34515000000
1!
1%
#34520000000
0!
0%
#34525000000
1!
1%
#34530000000
0!
0%
#34535000000
1!
1%
#34540000000
0!
0%
#34545000000
1!
1%
#34550000000
0!
0%
#34555000000
1!
1%
#34560000000
0!
0%
#34565000000
1!
1%
#34570000000
0!
0%
#34575000000
1!
1%
#34580000000
0!
0%
#34585000000
1!
1%
#34590000000
0!
0%
#34595000000
1!
1%
#34600000000
0!
0%
#34605000000
1!
1%
#34610000000
0!
0%
#34615000000
1!
1%
#34620000000
0!
0%
#34625000000
1!
1%
#34630000000
0!
0%
#34635000000
1!
1%
#34640000000
0!
0%
#34645000000
1!
1%
#34650000000
0!
0%
#34655000000
1!
1%
#34660000000
0!
0%
#34665000000
1!
1%
#34670000000
0!
0%
#34675000000
1!
1%
#34680000000
0!
0%
#34685000000
1!
1%
#34690000000
0!
0%
#34695000000
1!
1%
#34700000000
0!
0%
#34705000000
1!
1%
#34710000000
0!
0%
#34715000000
1!
1%
#34720000000
0!
0%
#34725000000
1!
1%
#34730000000
0!
0%
#34735000000
1!
1%
#34740000000
0!
0%
#34745000000
1!
1%
#34750000000
0!
0%
#34755000000
1!
1%
#34760000000
0!
0%
#34765000000
1!
1%
#34770000000
0!
0%
#34775000000
1!
1%
#34780000000
0!
0%
#34785000000
1!
1%
#34790000000
0!
0%
#34795000000
1!
1%
#34800000000
0!
0%
#34805000000
1!
1%
#34810000000
0!
0%
#34815000000
1!
1%
#34820000000
0!
0%
#34825000000
1!
1%
#34830000000
0!
0%
#34835000000
1!
1%
#34840000000
0!
0%
#34845000000
1!
1%
#34850000000
0!
0%
#34855000000
1!
1%
#34860000000
0!
0%
#34865000000
1!
1%
#34870000000
0!
0%
#34875000000
1!
1%
#34880000000
0!
0%
#34885000000
1!
1%
#34890000000
0!
0%
#34895000000
1!
1%
#34900000000
0!
0%
#34905000000
1!
1%
#34910000000
0!
0%
#34915000000
1!
1%
#34920000000
0!
0%
#34925000000
1!
1%
#34930000000
0!
0%
#34935000000
1!
1%
#34940000000
0!
0%
#34945000000
1!
1%
#34950000000
0!
0%
#34955000000
1!
1%
#34960000000
0!
0%
#34965000000
1!
1%
#34970000000
0!
0%
#34975000000
1!
1%
#34980000000
0!
0%
#34985000000
1!
1%
#34990000000
0!
0%
#34995000000
1!
1%
#35000000000
0!
0%
#35005000000
1!
1%
#35010000000
0!
0%
#35015000000
1!
1%
#35020000000
0!
0%
#35025000000
1!
1%
#35030000000
0!
0%
#35035000000
1!
1%
#35040000000
0!
0%
#35045000000
1!
1%
#35050000000
0!
0%
#35055000000
1!
1%
#35060000000
0!
0%
#35065000000
1!
1%
#35070000000
0!
0%
#35075000000
1!
1%
#35080000000
0!
0%
#35085000000
1!
1%
#35090000000
0!
0%
#35095000000
1!
1%
#35100000000
0!
0%
#35105000000
1!
1%
#35110000000
0!
0%
#35115000000
1!
1%
#35120000000
0!
0%
#35125000000
1!
1%
#35130000000
0!
0%
#35135000000
1!
1%
#35140000000
0!
0%
#35145000000
1!
1%
#35150000000
0!
0%
#35155000000
1!
1%
#35160000000
0!
0%
#35165000000
1!
1%
#35170000000
0!
0%
#35175000000
1!
1%
#35180000000
0!
0%
#35185000000
1!
1%
#35190000000
0!
0%
#35195000000
1!
1%
#35200000000
0!
0%
#35205000000
1!
1%
#35210000000
0!
0%
#35215000000
1!
1%
#35220000000
0!
0%
#35225000000
1!
1%
#35230000000
0!
0%
#35235000000
1!
1%
#35240000000
0!
0%
#35245000000
1!
1%
#35250000000
0!
0%
#35255000000
1!
1%
#35260000000
0!
0%
#35265000000
1!
1%
#35270000000
0!
0%
#35275000000
1!
1%
#35280000000
0!
0%
#35285000000
1!
1%
#35290000000
0!
0%
#35295000000
1!
1%
#35300000000
0!
0%
#35305000000
1!
1%
#35310000000
0!
0%
#35315000000
1!
1%
#35320000000
0!
0%
#35325000000
1!
1%
#35330000000
0!
0%
#35335000000
1!
1%
#35340000000
0!
0%
#35345000000
1!
1%
#35350000000
0!
0%
#35355000000
1!
1%
#35360000000
0!
0%
#35365000000
1!
1%
#35370000000
0!
0%
#35375000000
1!
1%
#35380000000
0!
0%
#35385000000
1!
1%
#35390000000
0!
0%
#35395000000
1!
1%
#35400000000
0!
0%
#35405000000
1!
1%
#35410000000
0!
0%
#35415000000
1!
1%
#35420000000
0!
0%
#35425000000
1!
1%
#35430000000
0!
0%
#35435000000
1!
1%
#35440000000
0!
0%
#35445000000
1!
1%
#35450000000
0!
0%
#35455000000
1!
1%
#35460000000
0!
0%
#35465000000
1!
1%
#35470000000
0!
0%
#35475000000
1!
1%
#35480000000
0!
0%
#35485000000
1!
1%
#35490000000
0!
0%
#35495000000
1!
1%
#35500000000
0!
0%
#35505000000
1!
1%
#35510000000
0!
0%
#35515000000
1!
1%
#35520000000
0!
0%
#35525000000
1!
1%
#35530000000
0!
0%
#35535000000
1!
1%
#35540000000
0!
0%
#35545000000
1!
1%
#35550000000
0!
0%
#35555000000
1!
1%
#35560000000
0!
0%
#35565000000
1!
1%
#35570000000
0!
0%
#35575000000
1!
1%
#35580000000
0!
0%
#35585000000
1!
1%
#35590000000
0!
0%
#35595000000
1!
1%
#35600000000
0!
0%
#35605000000
1!
1%
#35610000000
0!
0%
#35615000000
1!
1%
#35620000000
0!
0%
#35625000000
1!
1%
#35630000000
0!
0%
#35635000000
1!
1%
#35640000000
0!
0%
#35645000000
1!
1%
#35650000000
0!
0%
#35655000000
1!
1%
#35660000000
0!
0%
#35665000000
1!
1%
#35670000000
0!
0%
#35675000000
1!
1%
#35680000000
0!
0%
#35685000000
1!
1%
#35690000000
0!
0%
#35695000000
1!
1%
#35700000000
0!
0%
#35705000000
1!
1%
#35710000000
0!
0%
#35715000000
1!
1%
#35720000000
0!
0%
#35725000000
1!
1%
#35730000000
0!
0%
#35735000000
1!
1%
#35740000000
0!
0%
#35745000000
1!
1%
#35750000000
0!
0%
#35755000000
1!
1%
#35760000000
0!
0%
#35765000000
1!
1%
#35770000000
0!
0%
#35775000000
1!
1%
#35780000000
0!
0%
#35785000000
1!
1%
#35790000000
0!
0%
#35795000000
1!
1%
#35800000000
0!
0%
#35805000000
1!
1%
#35810000000
0!
0%
#35815000000
1!
1%
#35820000000
0!
0%
#35825000000
1!
1%
#35830000000
0!
0%
#35835000000
1!
1%
#35840000000
0!
0%
#35845000000
1!
1%
#35850000000
0!
0%
#35855000000
1!
1%
#35860000000
0!
0%
#35865000000
1!
1%
#35870000000
0!
0%
#35875000000
1!
1%
#35880000000
0!
0%
#35885000000
1!
1%
#35890000000
0!
0%
#35895000000
1!
1%
#35900000000
0!
0%
#35905000000
1!
1%
#35910000000
0!
0%
#35915000000
1!
1%
#35920000000
0!
0%
#35925000000
1!
1%
#35930000000
0!
0%
#35935000000
1!
1%
#35940000000
0!
0%
#35945000000
1!
1%
#35950000000
0!
0%
#35955000000
1!
1%
#35960000000
0!
0%
#35965000000
1!
1%
#35970000000
0!
0%
#35975000000
1!
1%
#35980000000
0!
0%
#35985000000
1!
1%
#35990000000
0!
0%
#35995000000
1!
1%
#36000000000
0!
0%
#36005000000
1!
1%
#36010000000
0!
0%
#36015000000
1!
1%
#36020000000
0!
0%
#36025000000
1!
1%
#36030000000
0!
0%
#36035000000
1!
1%
#36040000000
0!
0%
#36045000000
1!
1%
#36050000000
0!
0%
#36055000000
1!
1%
#36060000000
0!
0%
#36065000000
1!
1%
#36070000000
0!
0%
#36075000000
1!
1%
#36080000000
0!
0%
#36085000000
1!
1%
#36090000000
0!
0%
#36095000000
1!
1%
#36100000000
0!
0%
#36105000000
1!
1%
#36110000000
0!
0%
#36115000000
1!
1%
#36120000000
0!
0%
#36125000000
1!
1%
#36130000000
0!
0%
#36135000000
1!
1%
#36140000000
0!
0%
#36145000000
1!
1%
#36150000000
0!
0%
#36155000000
1!
1%
#36160000000
0!
0%
#36165000000
1!
1%
#36170000000
0!
0%
#36175000000
1!
1%
#36180000000
0!
0%
#36185000000
1!
1%
#36190000000
0!
0%
#36195000000
1!
1%
#36200000000
0!
0%
#36205000000
1!
1%
#36210000000
0!
0%
#36215000000
1!
1%
#36220000000
0!
0%
#36225000000
1!
1%
#36230000000
0!
0%
#36235000000
1!
1%
#36240000000
0!
0%
#36245000000
1!
1%
#36250000000
0!
0%
#36255000000
1!
1%
#36260000000
0!
0%
#36265000000
1!
1%
#36270000000
0!
0%
#36275000000
1!
1%
#36280000000
0!
0%
#36285000000
1!
1%
#36290000000
0!
0%
#36295000000
1!
1%
#36300000000
0!
0%
#36305000000
1!
1%
#36310000000
0!
0%
#36315000000
1!
1%
#36320000000
0!
0%
#36325000000
1!
1%
#36330000000
0!
0%
#36335000000
1!
1%
#36340000000
0!
0%
#36345000000
1!
1%
#36350000000
0!
0%
#36355000000
1!
1%
#36360000000
0!
0%
#36365000000
1!
1%
#36370000000
0!
0%
#36375000000
1!
1%
#36380000000
0!
0%
#36385000000
1!
1%
#36390000000
0!
0%
#36395000000
1!
1%
#36400000000
0!
0%
#36405000000
1!
1%
#36410000000
0!
0%
#36415000000
1!
1%
#36420000000
0!
0%
#36425000000
1!
1%
#36430000000
0!
0%
#36435000000
1!
1%
#36440000000
0!
0%
#36445000000
1!
1%
#36450000000
0!
0%
#36455000000
1!
1%
#36460000000
0!
0%
#36465000000
1!
1%
#36470000000
0!
0%
#36475000000
1!
1%
#36480000000
0!
0%
#36485000000
1!
1%
#36490000000
0!
0%
#36495000000
1!
1%
#36500000000
0!
0%
#36505000000
1!
1%
#36510000000
0!
0%
#36515000000
1!
1%
#36520000000
0!
0%
#36525000000
1!
1%
#36530000000
0!
0%
#36535000000
1!
1%
#36540000000
0!
0%
#36545000000
1!
1%
#36550000000
0!
0%
#36555000000
1!
1%
#36560000000
0!
0%
#36565000000
1!
1%
#36570000000
0!
0%
#36575000000
1!
1%
#36580000000
0!
0%
#36585000000
1!
1%
#36590000000
0!
0%
#36595000000
1!
1%
#36600000000
0!
0%
#36605000000
1!
1%
#36610000000
0!
0%
#36615000000
1!
1%
#36620000000
0!
0%
#36625000000
1!
1%
#36630000000
0!
0%
#36635000000
1!
1%
#36640000000
0!
0%
#36645000000
1!
1%
#36650000000
0!
0%
#36655000000
1!
1%
#36660000000
0!
0%
#36665000000
1!
1%
#36670000000
0!
0%
#36675000000
1!
1%
#36680000000
0!
0%
#36685000000
1!
1%
#36690000000
0!
0%
#36695000000
1!
1%
#36700000000
0!
0%
#36705000000
1!
1%
#36710000000
0!
0%
#36715000000
1!
1%
#36720000000
0!
0%
#36725000000
1!
1%
#36730000000
0!
0%
#36735000000
1!
1%
#36740000000
0!
0%
#36745000000
1!
1%
#36750000000
0!
0%
#36755000000
1!
1%
#36760000000
0!
0%
#36765000000
1!
1%
#36770000000
0!
0%
#36775000000
1!
1%
#36780000000
0!
0%
#36785000000
1!
1%
#36790000000
0!
0%
#36795000000
1!
1%
#36800000000
0!
0%
#36805000000
1!
1%
#36810000000
0!
0%
#36815000000
1!
1%
#36820000000
0!
0%
#36825000000
1!
1%
#36830000000
0!
0%
#36835000000
1!
1%
#36840000000
0!
0%
#36845000000
1!
1%
#36850000000
0!
0%
#36855000000
1!
1%
#36860000000
0!
0%
#36865000000
1!
1%
#36870000000
0!
0%
#36875000000
1!
1%
#36880000000
0!
0%
#36885000000
1!
1%
#36890000000
0!
0%
#36895000000
1!
1%
#36900000000
0!
0%
#36905000000
1!
1%
#36910000000
0!
0%
#36915000000
1!
1%
#36920000000
0!
0%
#36925000000
1!
1%
#36930000000
0!
0%
#36935000000
1!
1%
#36940000000
0!
0%
#36945000000
1!
1%
#36950000000
0!
0%
#36955000000
1!
1%
#36960000000
0!
0%
#36965000000
1!
1%
#36970000000
0!
0%
#36975000000
1!
1%
#36980000000
0!
0%
#36985000000
1!
1%
#36990000000
0!
0%
#36995000000
1!
1%
#37000000000
0!
0%
#37005000000
1!
1%
#37010000000
0!
0%
#37015000000
1!
1%
#37020000000
0!
0%
#37025000000
1!
1%
#37030000000
0!
0%
#37035000000
1!
1%
#37040000000
0!
0%
#37045000000
1!
1%
#37050000000
0!
0%
#37055000000
1!
1%
#37060000000
0!
0%
#37065000000
1!
1%
#37070000000
0!
0%
#37075000000
1!
1%
#37080000000
0!
0%
#37085000000
1!
1%
#37090000000
0!
0%
#37095000000
1!
1%
#37100000000
0!
0%
#37105000000
1!
1%
#37110000000
0!
0%
#37115000000
1!
1%
#37120000000
0!
0%
#37125000000
1!
1%
#37130000000
0!
0%
#37135000000
1!
1%
#37140000000
0!
0%
#37145000000
1!
1%
#37150000000
0!
0%
#37155000000
1!
1%
#37160000000
0!
0%
#37165000000
1!
1%
#37170000000
0!
0%
#37175000000
1!
1%
#37180000000
0!
0%
#37185000000
1!
1%
#37190000000
0!
0%
#37195000000
1!
1%
#37200000000
0!
0%
#37205000000
1!
1%
#37210000000
0!
0%
#37215000000
1!
1%
#37220000000
0!
0%
#37225000000
1!
1%
#37230000000
0!
0%
#37235000000
1!
1%
#37240000000
0!
0%
#37245000000
1!
1%
#37250000000
0!
0%
#37255000000
1!
1%
#37260000000
0!
0%
#37265000000
1!
1%
#37270000000
0!
0%
#37275000000
1!
1%
#37280000000
0!
0%
#37285000000
1!
1%
#37290000000
0!
0%
#37295000000
1!
1%
#37300000000
0!
0%
#37305000000
1!
1%
#37310000000
0!
0%
#37315000000
1!
1%
#37320000000
0!
0%
#37325000000
1!
1%
#37330000000
0!
0%
#37335000000
1!
1%
#37340000000
0!
0%
#37345000000
1!
1%
#37350000000
0!
0%
#37355000000
1!
1%
#37360000000
0!
0%
#37365000000
1!
1%
#37370000000
0!
0%
#37375000000
1!
1%
#37380000000
0!
0%
#37385000000
1!
1%
#37390000000
0!
0%
#37395000000
1!
1%
#37400000000
0!
0%
#37405000000
1!
1%
#37410000000
0!
0%
#37415000000
1!
1%
#37420000000
0!
0%
#37425000000
1!
1%
#37430000000
0!
0%
#37435000000
1!
1%
#37440000000
0!
0%
#37445000000
1!
1%
#37450000000
0!
0%
#37455000000
1!
1%
#37460000000
0!
0%
#37465000000
1!
1%
#37470000000
0!
0%
#37475000000
1!
1%
#37480000000
0!
0%
#37485000000
1!
1%
#37490000000
0!
0%
#37495000000
1!
1%
#37500000000
0!
0%
#37505000000
1!
1%
#37510000000
0!
0%
#37515000000
1!
1%
#37520000000
0!
0%
#37525000000
1!
1%
#37530000000
0!
0%
#37535000000
1!
1%
#37540000000
0!
0%
#37545000000
1!
1%
#37550000000
0!
0%
#37555000000
1!
1%
#37560000000
0!
0%
#37565000000
1!
1%
#37570000000
0!
0%
#37575000000
1!
1%
#37580000000
0!
0%
#37585000000
1!
1%
#37590000000
0!
0%
#37595000000
1!
1%
#37600000000
0!
0%
#37605000000
1!
1%
#37610000000
0!
0%
#37615000000
1!
1%
#37620000000
0!
0%
#37625000000
1!
1%
#37630000000
0!
0%
#37635000000
1!
1%
#37640000000
0!
0%
#37645000000
1!
1%
#37650000000
0!
0%
#37655000000
1!
1%
#37660000000
0!
0%
#37665000000
1!
1%
#37670000000
0!
0%
#37675000000
1!
1%
#37680000000
0!
0%
#37685000000
1!
1%
#37690000000
0!
0%
#37695000000
1!
1%
#37700000000
0!
0%
#37705000000
1!
1%
#37710000000
0!
0%
#37715000000
1!
1%
#37720000000
0!
0%
#37725000000
1!
1%
#37730000000
0!
0%
#37735000000
1!
1%
#37740000000
0!
0%
#37745000000
1!
1%
#37750000000
0!
0%
#37755000000
1!
1%
#37760000000
0!
0%
#37765000000
1!
1%
#37770000000
0!
0%
#37775000000
1!
1%
#37780000000
0!
0%
#37785000000
1!
1%
#37790000000
0!
0%
#37795000000
1!
1%
#37800000000
0!
0%
#37805000000
1!
1%
#37810000000
0!
0%
#37815000000
1!
1%
#37820000000
0!
0%
#37825000000
1!
1%
#37830000000
0!
0%
#37835000000
1!
1%
#37840000000
0!
0%
#37845000000
1!
1%
#37850000000
0!
0%
#37855000000
1!
1%
#37860000000
0!
0%
#37865000000
1!
1%
#37870000000
0!
0%
#37875000000
1!
1%
#37880000000
0!
0%
#37885000000
1!
1%
#37890000000
0!
0%
#37895000000
1!
1%
#37900000000
0!
0%
#37905000000
1!
1%
#37910000000
0!
0%
#37915000000
1!
1%
#37920000000
0!
0%
#37925000000
1!
1%
#37930000000
0!
0%
#37935000000
1!
1%
#37940000000
0!
0%
#37945000000
1!
1%
#37950000000
0!
0%
#37955000000
1!
1%
#37960000000
0!
0%
#37965000000
1!
1%
#37970000000
0!
0%
#37975000000
1!
1%
#37980000000
0!
0%
#37985000000
1!
1%
#37990000000
0!
0%
#37995000000
1!
1%
#38000000000
0!
0%
#38005000000
1!
1%
#38010000000
0!
0%
#38015000000
1!
1%
#38020000000
0!
0%
#38025000000
1!
1%
#38030000000
0!
0%
#38035000000
1!
1%
#38040000000
0!
0%
#38045000000
1!
1%
#38050000000
0!
0%
#38055000000
1!
1%
#38060000000
0!
0%
#38065000000
1!
1%
#38070000000
0!
0%
#38075000000
1!
1%
#38080000000
0!
0%
#38085000000
1!
1%
#38090000000
0!
0%
#38095000000
1!
1%
#38100000000
0!
0%
#38105000000
1!
1%
#38110000000
0!
0%
#38115000000
1!
1%
#38120000000
0!
0%
#38125000000
1!
1%
#38130000000
0!
0%
#38135000000
1!
1%
#38140000000
0!
0%
#38145000000
1!
1%
#38150000000
0!
0%
#38155000000
1!
1%
#38160000000
0!
0%
#38165000000
1!
1%
#38170000000
0!
0%
#38175000000
1!
1%
#38180000000
0!
0%
#38185000000
1!
1%
#38190000000
0!
0%
#38195000000
1!
1%
#38200000000
0!
0%
#38205000000
1!
1%
#38210000000
0!
0%
#38215000000
1!
1%
#38220000000
0!
0%
#38225000000
1!
1%
#38230000000
0!
0%
#38235000000
1!
1%
#38240000000
0!
0%
#38245000000
1!
1%
#38250000000
0!
0%
#38255000000
1!
1%
#38260000000
0!
0%
#38265000000
1!
1%
#38270000000
0!
0%
#38275000000
1!
1%
#38280000000
0!
0%
#38285000000
1!
1%
#38290000000
0!
0%
#38295000000
1!
1%
#38300000000
0!
0%
#38305000000
1!
1%
#38310000000
0!
0%
#38315000000
1!
1%
#38320000000
0!
0%
#38325000000
1!
1%
#38330000000
0!
0%
#38335000000
1!
1%
#38340000000
0!
0%
#38345000000
1!
1%
#38350000000
0!
0%
#38355000000
1!
1%
#38360000000
0!
0%
#38365000000
1!
1%
#38370000000
0!
0%
#38375000000
1!
1%
#38380000000
0!
0%
#38385000000
1!
1%
#38390000000
0!
0%
#38395000000
1!
1%
#38400000000
0!
0%
#38405000000
1!
1%
#38410000000
0!
0%
#38415000000
1!
1%
#38420000000
0!
0%
#38425000000
1!
1%
#38430000000
0!
0%
#38435000000
1!
1%
#38440000000
0!
0%
#38445000000
1!
1%
#38450000000
0!
0%
#38455000000
1!
1%
#38460000000
0!
0%
#38465000000
1!
1%
#38470000000
0!
0%
#38475000000
1!
1%
#38480000000
0!
0%
#38485000000
1!
1%
#38490000000
0!
0%
#38495000000
1!
1%
#38500000000
0!
0%
#38505000000
1!
1%
#38510000000
0!
0%
#38515000000
1!
1%
#38520000000
0!
0%
#38525000000
1!
1%
#38530000000
0!
0%
#38535000000
1!
1%
#38540000000
0!
0%
#38545000000
1!
1%
#38550000000
0!
0%
#38555000000
1!
1%
#38560000000
0!
0%
#38565000000
1!
1%
#38570000000
0!
0%
#38575000000
1!
1%
#38580000000
0!
0%
#38585000000
1!
1%
#38590000000
0!
0%
#38595000000
1!
1%
#38600000000
0!
0%
#38605000000
1!
1%
#38610000000
0!
0%
#38615000000
1!
1%
#38620000000
0!
0%
#38625000000
1!
1%
#38630000000
0!
0%
#38635000000
1!
1%
#38640000000
0!
0%
#38645000000
1!
1%
#38650000000
0!
0%
#38655000000
1!
1%
#38660000000
0!
0%
#38665000000
1!
1%
#38670000000
0!
0%
#38675000000
1!
1%
#38680000000
0!
0%
#38685000000
1!
1%
#38690000000
0!
0%
#38695000000
1!
1%
#38700000000
0!
0%
#38705000000
1!
1%
#38710000000
0!
0%
#38715000000
1!
1%
#38720000000
0!
0%
#38725000000
1!
1%
#38730000000
0!
0%
#38735000000
1!
1%
#38740000000
0!
0%
#38745000000
1!
1%
#38750000000
0!
0%
#38755000000
1!
1%
#38760000000
0!
0%
#38765000000
1!
1%
#38770000000
0!
0%
#38775000000
1!
1%
#38780000000
0!
0%
#38785000000
1!
1%
#38790000000
0!
0%
#38795000000
1!
1%
#38800000000
0!
0%
#38805000000
1!
1%
#38810000000
0!
0%
#38815000000
1!
1%
#38820000000
0!
0%
#38825000000
1!
1%
#38830000000
0!
0%
#38835000000
1!
1%
#38840000000
0!
0%
#38845000000
1!
1%
#38850000000
0!
0%
#38855000000
1!
1%
#38860000000
0!
0%
#38865000000
1!
1%
#38870000000
0!
0%
#38875000000
1!
1%
#38880000000
0!
0%
#38885000000
1!
1%
#38890000000
0!
0%
#38895000000
1!
1%
#38900000000
0!
0%
#38905000000
1!
1%
#38910000000
0!
0%
#38915000000
1!
1%
#38920000000
0!
0%
#38925000000
1!
1%
#38930000000
0!
0%
#38935000000
1!
1%
#38940000000
0!
0%
#38945000000
1!
1%
#38950000000
0!
0%
#38955000000
1!
1%
#38960000000
0!
0%
#38965000000
1!
1%
#38970000000
0!
0%
#38975000000
1!
1%
#38980000000
0!
0%
#38985000000
1!
1%
#38990000000
0!
0%
#38995000000
1!
1%
#39000000000
0!
0%
#39005000000
1!
1%
#39010000000
0!
0%
#39015000000
1!
1%
#39020000000
0!
0%
#39025000000
1!
1%
#39030000000
0!
0%
#39035000000
1!
1%
#39040000000
0!
0%
#39045000000
1!
1%
#39050000000
0!
0%
#39055000000
1!
1%
#39060000000
0!
0%
#39065000000
1!
1%
#39070000000
0!
0%
#39075000000
1!
1%
#39080000000
0!
0%
#39085000000
1!
1%
#39090000000
0!
0%
#39095000000
1!
1%
#39100000000
0!
0%
#39105000000
1!
1%
#39110000000
0!
0%
#39115000000
1!
1%
#39120000000
0!
0%
#39125000000
1!
1%
#39130000000
0!
0%
#39135000000
1!
1%
#39140000000
0!
0%
#39145000000
1!
1%
#39150000000
0!
0%
#39155000000
1!
1%
#39160000000
0!
0%
#39165000000
1!
1%
#39170000000
0!
0%
#39175000000
1!
1%
#39180000000
0!
0%
#39185000000
1!
1%
#39190000000
0!
0%
#39195000000
1!
1%
#39200000000
0!
0%
#39205000000
1!
1%
#39210000000
0!
0%
#39215000000
1!
1%
#39220000000
0!
0%
#39225000000
1!
1%
#39230000000
0!
0%
#39235000000
1!
1%
#39240000000
0!
0%
#39245000000
1!
1%
#39250000000
0!
0%
#39255000000
1!
1%
#39260000000
0!
0%
#39265000000
1!
1%
#39270000000
0!
0%
#39275000000
1!
1%
#39280000000
0!
0%
#39285000000
1!
1%
#39290000000
0!
0%
#39295000000
1!
1%
#39300000000
0!
0%
#39305000000
1!
1%
#39310000000
0!
0%
#39315000000
1!
1%
#39320000000
0!
0%
#39325000000
1!
1%
#39330000000
0!
0%
#39335000000
1!
1%
#39340000000
0!
0%
#39345000000
1!
1%
#39350000000
0!
0%
#39355000000
1!
1%
#39360000000
0!
0%
#39365000000
1!
1%
#39370000000
0!
0%
#39375000000
1!
1%
#39380000000
0!
0%
#39385000000
1!
1%
#39390000000
0!
0%
#39395000000
1!
1%
#39400000000
0!
0%
#39405000000
1!
1%
#39410000000
0!
0%
#39415000000
1!
1%
#39420000000
0!
0%
#39425000000
1!
1%
#39430000000
0!
0%
#39435000000
1!
1%
#39440000000
0!
0%
#39445000000
1!
1%
#39450000000
0!
0%
#39455000000
1!
1%
#39460000000
0!
0%
#39465000000
1!
1%
#39470000000
0!
0%
#39475000000
1!
1%
#39480000000
0!
0%
#39485000000
1!
1%
#39490000000
0!
0%
#39495000000
1!
1%
#39500000000
0!
0%
#39505000000
1!
1%
#39510000000
0!
0%
#39515000000
1!
1%
#39520000000
0!
0%
#39525000000
1!
1%
#39530000000
0!
0%
#39535000000
1!
1%
#39540000000
0!
0%
#39545000000
1!
1%
#39550000000
0!
0%
#39555000000
1!
1%
#39560000000
0!
0%
#39565000000
1!
1%
#39570000000
0!
0%
#39575000000
1!
1%
#39580000000
0!
0%
#39585000000
1!
1%
#39590000000
0!
0%
#39595000000
1!
1%
#39600000000
0!
0%
#39605000000
1!
1%
#39610000000
0!
0%
#39615000000
1!
1%
#39620000000
0!
0%
#39625000000
1!
1%
#39630000000
0!
0%
#39635000000
1!
1%
#39640000000
0!
0%
#39645000000
1!
1%
#39650000000
0!
0%
#39655000000
1!
1%
#39660000000
0!
0%
#39665000000
1!
1%
#39670000000
0!
0%
#39675000000
1!
1%
#39680000000
0!
0%
#39685000000
1!
1%
#39690000000
0!
0%
#39695000000
1!
1%
#39700000000
0!
0%
#39705000000
1!
1%
#39710000000
0!
0%
#39715000000
1!
1%
#39720000000
0!
0%
#39725000000
1!
1%
#39730000000
0!
0%
#39735000000
1!
1%
#39740000000
0!
0%
#39745000000
1!
1%
#39750000000
0!
0%
#39755000000
1!
1%
#39760000000
0!
0%
#39765000000
1!
1%
#39770000000
0!
0%
#39775000000
1!
1%
#39780000000
0!
0%
#39785000000
1!
1%
#39790000000
0!
0%
#39795000000
1!
1%
#39800000000
0!
0%
#39805000000
1!
1%
#39810000000
0!
0%
#39815000000
1!
1%
#39820000000
0!
0%
#39825000000
1!
1%
#39830000000
0!
0%
#39835000000
1!
1%
#39840000000
0!
0%
#39845000000
1!
1%
#39850000000
0!
0%
#39855000000
1!
1%
#39860000000
0!
0%
#39865000000
1!
1%
#39870000000
0!
0%
#39875000000
1!
1%
#39880000000
0!
0%
#39885000000
1!
1%
#39890000000
0!
0%
#39895000000
1!
1%
#39900000000
0!
0%
#39905000000
1!
1%
#39910000000
0!
0%
#39915000000
1!
1%
#39920000000
0!
0%
#39925000000
1!
1%
#39930000000
0!
0%
#39935000000
1!
1%
#39940000000
0!
0%
#39945000000
1!
1%
#39950000000
0!
0%
#39955000000
1!
1%
#39960000000
0!
0%
#39965000000
1!
1%
#39970000000
0!
0%
#39975000000
1!
1%
#39980000000
0!
0%
#39985000000
1!
1%
#39990000000
0!
0%
#39995000000
1!
1%
#40000000000
0!
0%
#40005000000
1!
1%
#40010000000
0!
0%
#40015000000
1!
1%
#40020000000
0!
0%
#40025000000
1!
1%
#40030000000
0!
0%
#40035000000
1!
1%
#40040000000
0!
0%
#40045000000
1!
1%
#40050000000
0!
0%
#40055000000
1!
1%
#40060000000
0!
0%
#40065000000
1!
1%
#40070000000
0!
0%
#40075000000
1!
1%
#40080000000
0!
0%
#40085000000
1!
1%
#40090000000
0!
0%
#40095000000
1!
1%
#40100000000
0!
0%
#40105000000
1!
1%
#40110000000
0!
0%
#40115000000
1!
1%
#40120000000
0!
0%
#40125000000
1!
1%
#40130000000
0!
0%
#40135000000
1!
1%
#40140000000
0!
0%
#40145000000
1!
1%
#40150000000
0!
0%
#40155000000
1!
1%
#40160000000
0!
0%
#40165000000
1!
1%
#40170000000
0!
0%
#40175000000
1!
1%
#40180000000
0!
0%
#40185000000
1!
1%
#40190000000
0!
0%
#40195000000
1!
1%
#40200000000
0!
0%
#40205000000
1!
1%
#40210000000
0!
0%
#40215000000
1!
1%
#40220000000
0!
0%
#40225000000
1!
1%
#40230000000
0!
0%
#40235000000
1!
1%
#40240000000
0!
0%
#40245000000
1!
1%
#40250000000
0!
0%
#40255000000
1!
1%
#40260000000
0!
0%
#40265000000
1!
1%
#40270000000
0!
0%
#40275000000
1!
1%
#40280000000
0!
0%
#40285000000
1!
1%
#40290000000
0!
0%
#40295000000
1!
1%
#40300000000
0!
0%
#40305000000
1!
1%
#40310000000
0!
0%
#40315000000
1!
1%
#40320000000
0!
0%
#40325000000
1!
1%
#40330000000
0!
0%
#40335000000
1!
1%
#40340000000
0!
0%
#40345000000
1!
1%
#40350000000
0!
0%
#40355000000
1!
1%
#40360000000
0!
0%
#40365000000
1!
1%
#40370000000
0!
0%
#40375000000
1!
1%
#40380000000
0!
0%
#40385000000
1!
1%
#40390000000
0!
0%
#40395000000
1!
1%
#40400000000
0!
0%
#40405000000
1!
1%
#40410000000
0!
0%
#40415000000
1!
1%
#40420000000
0!
0%
#40425000000
1!
1%
#40430000000
0!
0%
#40435000000
1!
1%
#40440000000
0!
0%
#40445000000
1!
1%
#40450000000
0!
0%
#40455000000
1!
1%
#40460000000
0!
0%
#40465000000
1!
1%
#40470000000
0!
0%
#40475000000
1!
1%
#40480000000
0!
0%
#40485000000
1!
1%
#40490000000
0!
0%
#40495000000
1!
1%
#40500000000
0!
0%
#40505000000
1!
1%
#40510000000
0!
0%
#40515000000
1!
1%
#40520000000
0!
0%
#40525000000
1!
1%
#40530000000
0!
0%
#40535000000
1!
1%
#40540000000
0!
0%
#40545000000
1!
1%
#40550000000
0!
0%
#40555000000
1!
1%
#40560000000
0!
0%
#40565000000
1!
1%
#40570000000
0!
0%
#40575000000
1!
1%
#40580000000
0!
0%
#40585000000
1!
1%
#40590000000
0!
0%
#40595000000
1!
1%
#40600000000
0!
0%
#40605000000
1!
1%
#40610000000
0!
0%
#40615000000
1!
1%
#40620000000
0!
0%
#40625000000
1!
1%
#40630000000
0!
0%
#40635000000
1!
1%
#40640000000
0!
0%
#40645000000
1!
1%
#40650000000
0!
0%
#40655000000
1!
1%
#40660000000
0!
0%
#40665000000
1!
1%
#40670000000
0!
0%
#40675000000
1!
1%
#40680000000
0!
0%
#40685000000
1!
1%
#40690000000
0!
0%
#40695000000
1!
1%
#40700000000
0!
0%
#40705000000
1!
1%
#40710000000
0!
0%
#40715000000
1!
1%
#40720000000
0!
0%
#40725000000
1!
1%
#40730000000
0!
0%
#40735000000
1!
1%
#40740000000
0!
0%
#40745000000
1!
1%
#40750000000
0!
0%
#40755000000
1!
1%
#40760000000
0!
0%
#40765000000
1!
1%
#40770000000
0!
0%
#40775000000
1!
1%
#40780000000
0!
0%
#40785000000
1!
1%
#40790000000
0!
0%
#40795000000
1!
1%
#40800000000
0!
0%
#40805000000
1!
1%
#40810000000
0!
0%
#40815000000
1!
1%
#40820000000
0!
0%
#40825000000
1!
1%
#40830000000
0!
0%
#40835000000
1!
1%
#40840000000
0!
0%
#40845000000
1!
1%
#40850000000
0!
0%
#40855000000
1!
1%
#40860000000
0!
0%
#40865000000
1!
1%
#40870000000
0!
0%
#40875000000
1!
1%
#40880000000
0!
0%
#40885000000
1!
1%
#40890000000
0!
0%
#40895000000
1!
1%
#40900000000
0!
0%
#40905000000
1!
1%
#40910000000
0!
0%
#40915000000
1!
1%
#40920000000
0!
0%
#40925000000
1!
1%
#40930000000
0!
0%
#40935000000
1!
1%
#40940000000
0!
0%
#40945000000
1!
1%
#40950000000
0!
0%
#40955000000
1!
1%
#40960000000
0!
0%
#40965000000
1!
1%
#40970000000
0!
0%
#40975000000
1!
1%
#40980000000
0!
0%
#40985000000
1!
1%
#40990000000
0!
0%
#40995000000
1!
1%
#41000000000
0!
0%
#41005000000
1!
1%
#41010000000
0!
0%
#41015000000
1!
1%
#41020000000
0!
0%
#41025000000
1!
1%
#41030000000
0!
0%
#41035000000
1!
1%
#41040000000
0!
0%
#41045000000
1!
1%
#41050000000
0!
0%
#41055000000
1!
1%
#41060000000
0!
0%
#41065000000
1!
1%
#41070000000
0!
0%
#41075000000
1!
1%
#41080000000
0!
0%
#41085000000
1!
1%
#41090000000
0!
0%
#41095000000
1!
1%
#41100000000
0!
0%
#41105000000
1!
1%
#41110000000
0!
0%
#41115000000
1!
1%
#41120000000
0!
0%
#41125000000
1!
1%
#41130000000
0!
0%
#41135000000
1!
1%
#41140000000
0!
0%
#41145000000
1!
1%
#41150000000
0!
0%
#41155000000
1!
1%
#41160000000
0!
0%
#41165000000
1!
1%
#41170000000
0!
0%
#41175000000
1!
1%
#41180000000
0!
0%
#41185000000
1!
1%
#41190000000
0!
0%
#41195000000
1!
1%
#41200000000
0!
0%
#41205000000
1!
1%
#41210000000
0!
0%
#41215000000
1!
1%
#41220000000
0!
0%
#41225000000
1!
1%
#41230000000
0!
0%
#41235000000
1!
1%
#41240000000
0!
0%
#41245000000
1!
1%
#41250000000
0!
0%
#41255000000
1!
1%
#41260000000
0!
0%
#41265000000
1!
1%
#41270000000
0!
0%
#41275000000
1!
1%
#41280000000
0!
0%
#41285000000
1!
1%
#41290000000
0!
0%
#41295000000
1!
1%
#41300000000
0!
0%
#41305000000
1!
1%
#41310000000
0!
0%
#41315000000
1!
1%
#41320000000
0!
0%
#41325000000
1!
1%
#41330000000
0!
0%
#41335000000
1!
1%
#41340000000
0!
0%
#41345000000
1!
1%
#41350000000
0!
0%
#41355000000
1!
1%
#41360000000
0!
0%
#41365000000
1!
1%
#41370000000
0!
0%
#41375000000
1!
1%
#41380000000
0!
0%
#41385000000
1!
1%
#41390000000
0!
0%
#41395000000
1!
1%
#41400000000
0!
0%
#41405000000
1!
1%
#41410000000
0!
0%
#41415000000
1!
1%
#41420000000
0!
0%
#41425000000
1!
1%
#41430000000
0!
0%
#41435000000
1!
1%
#41440000000
0!
0%
#41445000000
1!
1%
#41450000000
0!
0%
#41455000000
1!
1%
#41460000000
0!
0%
#41465000000
1!
1%
#41470000000
0!
0%
#41475000000
1!
1%
#41480000000
0!
0%
#41485000000
1!
1%
#41490000000
0!
0%
#41495000000
1!
1%
#41500000000
0!
0%
#41505000000
1!
1%
#41510000000
0!
0%
#41515000000
1!
1%
#41520000000
0!
0%
#41525000000
1!
1%
#41530000000
0!
0%
#41535000000
1!
1%
#41540000000
0!
0%
#41545000000
1!
1%
#41550000000
0!
0%
#41555000000
1!
1%
#41560000000
0!
0%
#41565000000
1!
1%
#41570000000
0!
0%
#41575000000
1!
1%
#41580000000
0!
0%
#41585000000
1!
1%
#41590000000
0!
0%
#41595000000
1!
1%
#41600000000
0!
0%
#41605000000
1!
1%
#41610000000
0!
0%
#41615000000
1!
1%
#41620000000
0!
0%
#41625000000
1!
1%
#41630000000
0!
0%
#41635000000
1!
1%
#41640000000
0!
0%
#41645000000
1!
1%
#41650000000
0!
0%
#41655000000
1!
1%
#41660000000
0!
0%
#41665000000
1!
1%
#41670000000
0!
0%
#41675000000
1!
1%
#41680000000
0!
0%
#41685000000
1!
1%
#41690000000
0!
0%
#41695000000
1!
1%
#41700000000
0!
0%
#41705000000
1!
1%
#41710000000
0!
0%
#41715000000
1!
1%
#41720000000
0!
0%
#41725000000
1!
1%
#41730000000
0!
0%
#41735000000
1!
1%
#41740000000
0!
0%
#41745000000
1!
1%
#41750000000
0!
0%
#41755000000
1!
1%
#41760000000
0!
0%
#41765000000
1!
1%
#41770000000
0!
0%
#41775000000
1!
1%
#41780000000
0!
0%
#41785000000
1!
1%
#41790000000
0!
0%
#41795000000
1!
1%
#41800000000
0!
0%
#41805000000
1!
1%
#41810000000
0!
0%
#41815000000
1!
1%
#41820000000
0!
0%
#41825000000
1!
1%
#41830000000
0!
0%
#41835000000
1!
1%
#41840000000
0!
0%
#41845000000
1!
1%
#41850000000
0!
0%
#41855000000
1!
1%
#41860000000
0!
0%
#41865000000
1!
1%
#41870000000
0!
0%
#41875000000
1!
1%
#41880000000
0!
0%
#41885000000
1!
1%
#41890000000
0!
0%
#41895000000
1!
1%
#41900000000
0!
0%
#41905000000
1!
1%
#41910000000
0!
0%
#41915000000
1!
1%
#41920000000
0!
0%
#41925000000
1!
1%
#41930000000
0!
0%
#41935000000
1!
1%
#41940000000
0!
0%
#41945000000
1!
1%
#41950000000
0!
0%
#41955000000
1!
1%
#41960000000
0!
0%
#41965000000
1!
1%
#41970000000
0!
0%
#41975000000
1!
1%
#41980000000
0!
0%
#41985000000
1!
1%
#41990000000
0!
0%
#41995000000
1!
1%
#42000000000
0!
0%
#42005000000
1!
1%
#42010000000
0!
0%
#42015000000
1!
1%
#42020000000
0!
0%
#42025000000
1!
1%
#42030000000
0!
0%
#42035000000
1!
1%
#42040000000
0!
0%
#42045000000
1!
1%
#42050000000
0!
0%
#42055000000
1!
1%
#42060000000
0!
0%
#42065000000
1!
1%
#42070000000
0!
0%
#42075000000
1!
1%
#42080000000
0!
0%
#42085000000
1!
1%
#42090000000
0!
0%
#42095000000
1!
1%
#42100000000
0!
0%
#42105000000
1!
1%
#42110000000
0!
0%
#42115000000
1!
1%
#42120000000
0!
0%
#42125000000
1!
1%
#42130000000
0!
0%
#42135000000
1!
1%
#42140000000
0!
0%
#42145000000
1!
1%
#42150000000
0!
0%
#42155000000
1!
1%
#42160000000
0!
0%
#42165000000
1!
1%
#42170000000
0!
0%
#42175000000
1!
1%
#42180000000
0!
0%
#42185000000
1!
1%
#42190000000
0!
0%
#42195000000
1!
1%
#42200000000
0!
0%
#42205000000
1!
1%
#42210000000
0!
0%
#42215000000
1!
1%
#42220000000
0!
0%
#42225000000
1!
1%
#42230000000
0!
0%
#42235000000
1!
1%
#42240000000
0!
0%
#42245000000
1!
1%
#42250000000
0!
0%
#42255000000
1!
1%
#42260000000
0!
0%
#42265000000
1!
1%
#42270000000
0!
0%
#42275000000
1!
1%
#42280000000
0!
0%
#42285000000
1!
1%
#42290000000
0!
0%
#42295000000
1!
1%
#42300000000
0!
0%
#42305000000
1!
1%
#42310000000
0!
0%
#42315000000
1!
1%
#42320000000
0!
0%
#42325000000
1!
1%
#42330000000
0!
0%
#42335000000
1!
1%
#42340000000
0!
0%
#42345000000
1!
1%
#42350000000
0!
0%
#42355000000
1!
1%
#42360000000
0!
0%
#42365000000
1!
1%
#42370000000
0!
0%
#42375000000
1!
1%
#42380000000
0!
0%
#42385000000
1!
1%
#42390000000
0!
0%
#42395000000
1!
1%
#42400000000
0!
0%
#42405000000
1!
1%
#42410000000
0!
0%
#42415000000
1!
1%
#42420000000
0!
0%
#42425000000
1!
1%
#42430000000
0!
0%
#42435000000
1!
1%
#42440000000
0!
0%
#42445000000
1!
1%
#42450000000
0!
0%
#42455000000
1!
1%
#42460000000
0!
0%
#42465000000
1!
1%
#42470000000
0!
0%
#42475000000
1!
1%
#42480000000
0!
0%
#42485000000
1!
1%
#42490000000
0!
0%
#42495000000
1!
1%
#42500000000
0!
0%
#42505000000
1!
1%
#42510000000
0!
0%
#42515000000
1!
1%
#42520000000
0!
0%
#42525000000
1!
1%
#42530000000
0!
0%
#42535000000
1!
1%
#42540000000
0!
0%
#42545000000
1!
1%
#42550000000
0!
0%
#42555000000
1!
1%
#42560000000
0!
0%
#42565000000
1!
1%
#42570000000
0!
0%
#42575000000
1!
1%
#42580000000
0!
0%
#42585000000
1!
1%
#42590000000
0!
0%
#42595000000
1!
1%
#42600000000
0!
0%
#42605000000
1!
1%
#42610000000
0!
0%
#42615000000
1!
1%
#42620000000
0!
0%
#42625000000
1!
1%
#42630000000
0!
0%
#42635000000
1!
1%
#42640000000
0!
0%
#42645000000
1!
1%
#42650000000
0!
0%
#42655000000
1!
1%
#42660000000
0!
0%
#42665000000
1!
1%
#42670000000
0!
0%
#42675000000
1!
1%
#42680000000
0!
0%
#42685000000
1!
1%
#42690000000
0!
0%
#42695000000
1!
1%
#42700000000
0!
0%
#42705000000
1!
1%
#42710000000
0!
0%
#42715000000
1!
1%
#42720000000
0!
0%
#42725000000
1!
1%
#42730000000
0!
0%
#42735000000
1!
1%
#42740000000
0!
0%
#42745000000
1!
1%
#42750000000
0!
0%
#42755000000
1!
1%
#42760000000
0!
0%
#42765000000
1!
1%
#42770000000
0!
0%
#42775000000
1!
1%
#42780000000
0!
0%
#42785000000
1!
1%
#42790000000
0!
0%
#42795000000
1!
1%
#42800000000
0!
0%
#42805000000
1!
1%
#42810000000
0!
0%
#42815000000
1!
1%
#42820000000
0!
0%
#42825000000
1!
1%
#42830000000
0!
0%
#42835000000
1!
1%
#42840000000
0!
0%
#42845000000
1!
1%
#42850000000
0!
0%
#42855000000
1!
1%
#42860000000
0!
0%
#42865000000
1!
1%
#42870000000
0!
0%
#42875000000
1!
1%
#42880000000
0!
0%
#42885000000
1!
1%
#42890000000
0!
0%
#42895000000
1!
1%
#42900000000
0!
0%
#42905000000
1!
1%
#42910000000
0!
0%
#42915000000
1!
1%
#42920000000
0!
0%
#42925000000
1!
1%
#42930000000
0!
0%
#42935000000
1!
1%
#42940000000
0!
0%
#42945000000
1!
1%
#42950000000
0!
0%
#42955000000
1!
1%
#42960000000
0!
0%
#42965000000
1!
1%
#42970000000
0!
0%
#42975000000
1!
1%
#42980000000
0!
0%
#42985000000
1!
1%
#42990000000
0!
0%
#42995000000
1!
1%
#43000000000
0!
0%
#43005000000
1!
1%
#43010000000
0!
0%
#43015000000
1!
1%
#43020000000
0!
0%
#43025000000
1!
1%
#43030000000
0!
0%
#43035000000
1!
1%
#43040000000
0!
0%
#43045000000
1!
1%
#43050000000
0!
0%
#43055000000
1!
1%
#43060000000
0!
0%
#43065000000
1!
1%
#43070000000
0!
0%
#43075000000
1!
1%
#43080000000
0!
0%
#43085000000
1!
1%
#43090000000
0!
0%
#43095000000
1!
1%
#43100000000
0!
0%
#43105000000
1!
1%
#43110000000
0!
0%
#43115000000
1!
1%
#43120000000
0!
0%
#43125000000
1!
1%
#43130000000
0!
0%
#43135000000
1!
1%
#43140000000
0!
0%
#43145000000
1!
1%
#43150000000
0!
0%
#43155000000
1!
1%
#43160000000
0!
0%
#43165000000
1!
1%
#43170000000
0!
0%
#43175000000
1!
1%
#43180000000
0!
0%
#43185000000
1!
1%
#43190000000
0!
0%
#43195000000
1!
1%
#43200000000
0!
0%
#43205000000
1!
1%
#43210000000
0!
0%
#43215000000
1!
1%
#43220000000
0!
0%
#43225000000
1!
1%
#43230000000
0!
0%
#43235000000
1!
1%
#43240000000
0!
0%
#43245000000
1!
1%
#43250000000
0!
0%
#43255000000
1!
1%
#43260000000
0!
0%
#43265000000
1!
1%
#43270000000
0!
0%
#43275000000
1!
1%
#43280000000
0!
0%
#43285000000
1!
1%
#43290000000
0!
0%
#43295000000
1!
1%
#43300000000
0!
0%
#43305000000
1!
1%
#43310000000
0!
0%
#43315000000
1!
1%
#43320000000
0!
0%
#43325000000
1!
1%
#43330000000
0!
0%
#43335000000
1!
1%
#43340000000
0!
0%
#43345000000
1!
1%
#43350000000
0!
0%
#43355000000
1!
1%
#43360000000
0!
0%
#43365000000
1!
1%
#43370000000
0!
0%
#43375000000
1!
1%
#43380000000
0!
0%
#43385000000
1!
1%
#43390000000
0!
0%
#43395000000
1!
1%
#43400000000
0!
0%
#43405000000
1!
1%
#43410000000
0!
0%
#43415000000
1!
1%
#43420000000
0!
0%
#43425000000
1!
1%
#43430000000
0!
0%
#43435000000
1!
1%
#43440000000
0!
0%
#43445000000
1!
1%
#43450000000
0!
0%
#43455000000
1!
1%
#43460000000
0!
0%
#43465000000
1!
1%
#43470000000
0!
0%
#43475000000
1!
1%
#43480000000
0!
0%
#43485000000
1!
1%
#43490000000
0!
0%
#43495000000
1!
1%
#43500000000
0!
0%
#43505000000
1!
1%
#43510000000
0!
0%
#43515000000
1!
1%
#43520000000
0!
0%
#43525000000
1!
1%
#43530000000
0!
0%
#43535000000
1!
1%
#43540000000
0!
0%
#43545000000
1!
1%
#43550000000
0!
0%
#43555000000
1!
1%
#43560000000
0!
0%
#43565000000
1!
1%
#43570000000
0!
0%
#43575000000
1!
1%
#43580000000
0!
0%
#43585000000
1!
1%
#43590000000
0!
0%
#43595000000
1!
1%
#43600000000
0!
0%
#43605000000
1!
1%
#43610000000
0!
0%
#43615000000
1!
1%
#43620000000
0!
0%
#43625000000
1!
1%
#43630000000
0!
0%
#43635000000
1!
1%
#43640000000
0!
0%
#43645000000
1!
1%
#43650000000
0!
0%
#43655000000
1!
1%
#43660000000
0!
0%
#43665000000
1!
1%
#43670000000
0!
0%
#43675000000
1!
1%
#43680000000
0!
0%
#43685000000
1!
1%
#43690000000
0!
0%
#43695000000
1!
1%
#43700000000
0!
0%
#43705000000
1!
1%
#43710000000
0!
0%
#43715000000
1!
1%
#43720000000
0!
0%
#43725000000
1!
1%
#43730000000
0!
0%
#43735000000
1!
1%
#43740000000
0!
0%
#43745000000
1!
1%
#43750000000
0!
0%
#43755000000
1!
1%
#43760000000
0!
0%
#43765000000
1!
1%
#43770000000
0!
0%
#43775000000
1!
1%
#43780000000
0!
0%
#43785000000
1!
1%
#43790000000
0!
0%
#43795000000
1!
1%
#43800000000
0!
0%
#43805000000
1!
1%
#43810000000
0!
0%
#43815000000
1!
1%
#43820000000
0!
0%
#43825000000
1!
1%
#43830000000
0!
0%
#43835000000
1!
1%
#43840000000
0!
0%
#43845000000
1!
1%
#43850000000
0!
0%
#43855000000
1!
1%
#43860000000
0!
0%
#43865000000
1!
1%
#43870000000
0!
0%
#43875000000
1!
1%
#43880000000
0!
0%
#43885000000
1!
1%
#43890000000
0!
0%
#43895000000
1!
1%
#43900000000
0!
0%
#43905000000
1!
1%
#43910000000
0!
0%
#43915000000
1!
1%
#43920000000
0!
0%
#43925000000
1!
1%
#43930000000
0!
0%
#43935000000
1!
1%
#43940000000
0!
0%
#43945000000
1!
1%
#43950000000
0!
0%
#43955000000
1!
1%
#43960000000
0!
0%
#43965000000
1!
1%
#43970000000
0!
0%
#43975000000
1!
1%
#43980000000
0!
0%
#43985000000
1!
1%
#43990000000
0!
0%
#43995000000
1!
1%
#44000000000
0!
0%
#44005000000
1!
1%
#44010000000
0!
0%
#44015000000
1!
1%
#44020000000
0!
0%
#44025000000
1!
1%
#44030000000
0!
0%
#44035000000
1!
1%
#44040000000
0!
0%
#44045000000
1!
1%
#44050000000
0!
0%
#44055000000
1!
1%
#44060000000
0!
0%
#44065000000
1!
1%
#44070000000
0!
0%
#44075000000
1!
1%
#44080000000
0!
0%
#44085000000
1!
1%
#44090000000
0!
0%
#44095000000
1!
1%
#44100000000
0!
0%
#44105000000
1!
1%
#44110000000
0!
0%
#44115000000
1!
1%
#44120000000
0!
0%
#44125000000
1!
1%
#44130000000
0!
0%
#44135000000
1!
1%
#44140000000
0!
0%
#44145000000
1!
1%
#44150000000
0!
0%
#44155000000
1!
1%
#44160000000
0!
0%
#44165000000
1!
1%
#44170000000
0!
0%
#44175000000
1!
1%
#44180000000
0!
0%
#44185000000
1!
1%
#44190000000
0!
0%
#44195000000
1!
1%
#44200000000
0!
0%
#44205000000
1!
1%
#44210000000
0!
0%
#44215000000
1!
1%
#44220000000
0!
0%
#44225000000
1!
1%
#44230000000
0!
0%
#44235000000
1!
1%
#44240000000
0!
0%
#44245000000
1!
1%
#44250000000
0!
0%
#44255000000
1!
1%
#44260000000
0!
0%
#44265000000
1!
1%
#44270000000
0!
0%
#44275000000
1!
1%
#44280000000
0!
0%
#44285000000
1!
1%
#44290000000
0!
0%
#44295000000
1!
1%
#44300000000
0!
0%
#44305000000
1!
1%
#44310000000
0!
0%
#44315000000
1!
1%
#44320000000
0!
0%
#44325000000
1!
1%
#44330000000
0!
0%
#44335000000
1!
1%
#44340000000
0!
0%
#44345000000
1!
1%
#44350000000
0!
0%
#44355000000
1!
1%
#44360000000
0!
0%
#44365000000
1!
1%
#44370000000
0!
0%
#44375000000
1!
1%
#44380000000
0!
0%
#44385000000
1!
1%
#44390000000
0!
0%
#44395000000
1!
1%
#44400000000
0!
0%
#44405000000
1!
1%
#44410000000
0!
0%
#44415000000
1!
1%
#44420000000
0!
0%
#44425000000
1!
1%
#44430000000
0!
0%
#44435000000
1!
1%
#44440000000
0!
0%
#44445000000
1!
1%
#44450000000
0!
0%
#44455000000
1!
1%
#44460000000
0!
0%
#44465000000
1!
1%
#44470000000
0!
0%
#44475000000
1!
1%
#44480000000
0!
0%
#44485000000
1!
1%
#44490000000
0!
0%
#44495000000
1!
1%
#44500000000
0!
0%
#44505000000
1!
1%
#44510000000
0!
0%
#44515000000
1!
1%
#44520000000
0!
0%
#44525000000
1!
1%
#44530000000
0!
0%
#44535000000
1!
1%
#44540000000
0!
0%
#44545000000
1!
1%
#44550000000
0!
0%
#44555000000
1!
1%
#44560000000
0!
0%
#44565000000
1!
1%
#44570000000
0!
0%
#44575000000
1!
1%
#44580000000
0!
0%
#44585000000
1!
1%
#44590000000
0!
0%
#44595000000
1!
1%
#44600000000
0!
0%
#44605000000
1!
1%
#44610000000
0!
0%
#44615000000
1!
1%
#44620000000
0!
0%
#44625000000
1!
1%
#44630000000
0!
0%
#44635000000
1!
1%
#44640000000
0!
0%
#44645000000
1!
1%
#44650000000
0!
0%
#44655000000
1!
1%
#44660000000
0!
0%
#44665000000
1!
1%
#44670000000
0!
0%
#44675000000
1!
1%
#44680000000
0!
0%
#44685000000
1!
1%
#44690000000
0!
0%
#44695000000
1!
1%
#44700000000
0!
0%
#44705000000
1!
1%
#44710000000
0!
0%
#44715000000
1!
1%
#44720000000
0!
0%
#44725000000
1!
1%
#44730000000
0!
0%
#44735000000
1!
1%
#44740000000
0!
0%
#44745000000
1!
1%
#44750000000
0!
0%
#44755000000
1!
1%
#44760000000
0!
0%
#44765000000
1!
1%
#44770000000
0!
0%
#44775000000
1!
1%
#44780000000
0!
0%
#44785000000
1!
1%
#44790000000
0!
0%
#44795000000
1!
1%
#44800000000
0!
0%
#44805000000
1!
1%
#44810000000
0!
0%
#44815000000
1!
1%
#44820000000
0!
0%
#44825000000
1!
1%
#44830000000
0!
0%
#44835000000
1!
1%
#44840000000
0!
0%
#44845000000
1!
1%
#44850000000
0!
0%
#44855000000
1!
1%
#44860000000
0!
0%
#44865000000
1!
1%
#44870000000
0!
0%
#44875000000
1!
1%
#44880000000
0!
0%
#44885000000
1!
1%
#44890000000
0!
0%
#44895000000
1!
1%
#44900000000
0!
0%
#44905000000
1!
1%
#44910000000
0!
0%
#44915000000
1!
1%
#44920000000
0!
0%
#44925000000
1!
1%
#44930000000
0!
0%
#44935000000
1!
1%
#44940000000
0!
0%
#44945000000
1!
1%
#44950000000
0!
0%
#44955000000
1!
1%
#44960000000
0!
0%
#44965000000
1!
1%
#44970000000
0!
0%
#44975000000
1!
1%
#44980000000
0!
0%
#44985000000
1!
1%
#44990000000
0!
0%
#44995000000
1!
1%
#45000000000
0!
0%
#45005000000
1!
1%
#45010000000
0!
0%
#45015000000
1!
1%
#45020000000
0!
0%
#45025000000
1!
1%
#45030000000
0!
0%
#45035000000
1!
1%
#45040000000
0!
0%
#45045000000
1!
1%
#45050000000
0!
0%
#45055000000
1!
1%
#45060000000
0!
0%
#45065000000
1!
1%
#45070000000
0!
0%
#45075000000
1!
1%
#45080000000
0!
0%
#45085000000
1!
1%
#45090000000
0!
0%
#45095000000
1!
1%
#45100000000
0!
0%
#45105000000
1!
1%
#45110000000
0!
0%
#45115000000
1!
1%
#45120000000
0!
0%
#45125000000
1!
1%
#45130000000
0!
0%
#45135000000
1!
1%
#45140000000
0!
0%
#45145000000
1!
1%
#45150000000
0!
0%
#45155000000
1!
1%
#45160000000
0!
0%
#45165000000
1!
1%
#45170000000
0!
0%
#45175000000
1!
1%
#45180000000
0!
0%
#45185000000
1!
1%
#45190000000
0!
0%
#45195000000
1!
1%
#45200000000
0!
0%
#45205000000
1!
1%
#45210000000
0!
0%
#45215000000
1!
1%
#45220000000
0!
0%
#45225000000
1!
1%
#45230000000
0!
0%
#45235000000
1!
1%
#45240000000
0!
0%
#45245000000
1!
1%
#45250000000
0!
0%
#45255000000
1!
1%
#45260000000
0!
0%
#45265000000
1!
1%
#45270000000
0!
0%
#45275000000
1!
1%
#45280000000
0!
0%
#45285000000
1!
1%
#45290000000
0!
0%
#45295000000
1!
1%
#45300000000
0!
0%
#45305000000
1!
1%
#45310000000
0!
0%
#45315000000
1!
1%
#45320000000
0!
0%
#45325000000
1!
1%
#45330000000
0!
0%
#45335000000
1!
1%
#45340000000
0!
0%
#45345000000
1!
1%
#45350000000
0!
0%
#45355000000
1!
1%
#45360000000
0!
0%
#45365000000
1!
1%
#45370000000
0!
0%
#45375000000
1!
1%
#45380000000
0!
0%
#45385000000
1!
1%
#45390000000
0!
0%
#45395000000
1!
1%
#45400000000
0!
0%
#45405000000
1!
1%
#45410000000
0!
0%
#45415000000
1!
1%
#45420000000
0!
0%
#45425000000
1!
1%
#45430000000
0!
0%
#45435000000
1!
1%
#45440000000
0!
0%
#45445000000
1!
1%
#45450000000
0!
0%
#45455000000
1!
1%
#45460000000
0!
0%
#45465000000
1!
1%
#45470000000
0!
0%
#45475000000
1!
1%
#45480000000
0!
0%
#45485000000
1!
1%
#45490000000
0!
0%
#45495000000
1!
1%
#45500000000
0!
0%
#45505000000
1!
1%
#45510000000
0!
0%
#45515000000
1!
1%
#45520000000
0!
0%
#45525000000
1!
1%
#45530000000
0!
0%
#45535000000
1!
1%
#45540000000
0!
0%
#45545000000
1!
1%
#45550000000
0!
0%
#45555000000
1!
1%
#45560000000
0!
0%
#45565000000
1!
1%
#45570000000
0!
0%
#45575000000
1!
1%
#45580000000
0!
0%
#45585000000
1!
1%
#45590000000
0!
0%
#45595000000
1!
1%
#45600000000
0!
0%
#45605000000
1!
1%
#45610000000
0!
0%
#45615000000
1!
1%
#45620000000
0!
0%
#45625000000
1!
1%
#45630000000
0!
0%
#45635000000
1!
1%
#45640000000
0!
0%
#45645000000
1!
1%
#45650000000
0!
0%
#45655000000
1!
1%
#45660000000
0!
0%
#45665000000
1!
1%
#45670000000
0!
0%
#45675000000
1!
1%
#45680000000
0!
0%
#45685000000
1!
1%
#45690000000
0!
0%
#45695000000
1!
1%
#45700000000
0!
0%
#45705000000
1!
1%
#45710000000
0!
0%
#45715000000
1!
1%
#45720000000
0!
0%
#45725000000
1!
1%
#45730000000
0!
0%
#45735000000
1!
1%
#45740000000
0!
0%
#45745000000
1!
1%
#45750000000
0!
0%
#45755000000
1!
1%
#45760000000
0!
0%
#45765000000
1!
1%
#45770000000
0!
0%
#45775000000
1!
1%
#45780000000
0!
0%
#45785000000
1!
1%
#45790000000
0!
0%
#45795000000
1!
1%
#45800000000
0!
0%
#45805000000
1!
1%
#45810000000
0!
0%
#45815000000
1!
1%
#45820000000
0!
0%
#45825000000
1!
1%
#45830000000
0!
0%
#45835000000
1!
1%
#45840000000
0!
0%
#45845000000
1!
1%
#45850000000
0!
0%
#45855000000
1!
1%
#45860000000
0!
0%
#45865000000
1!
1%
#45870000000
0!
0%
#45875000000
1!
1%
#45880000000
0!
0%
#45885000000
1!
1%
#45890000000
0!
0%
#45895000000
1!
1%
#45900000000
0!
0%
#45905000000
1!
1%
#45910000000
0!
0%
#45915000000
1!
1%
#45920000000
0!
0%
#45925000000
1!
1%
#45930000000
0!
0%
#45935000000
1!
1%
#45940000000
0!
0%
#45945000000
1!
1%
#45950000000
0!
0%
#45955000000
1!
1%
#45960000000
0!
0%
#45965000000
1!
1%
#45970000000
0!
0%
#45975000000
1!
1%
#45980000000
0!
0%
#45985000000
1!
1%
#45990000000
0!
0%
#45995000000
1!
1%
#46000000000
0!
0%
#46005000000
1!
1%
#46010000000
0!
0%
#46015000000
1!
1%
#46020000000
0!
0%
#46025000000
1!
1%
#46030000000
0!
0%
#46035000000
1!
1%
#46040000000
0!
0%
#46045000000
1!
1%
#46050000000
0!
0%
#46055000000
1!
1%
#46060000000
0!
0%
#46065000000
1!
1%
#46070000000
0!
0%
#46075000000
1!
1%
#46080000000
0!
0%
#46085000000
1!
1%
#46090000000
0!
0%
#46095000000
1!
1%
#46100000000
0!
0%
#46105000000
1!
1%
#46110000000
0!
0%
#46115000000
1!
1%
#46120000000
0!
0%
#46125000000
1!
1%
#46130000000
0!
0%
#46135000000
1!
1%
#46140000000
0!
0%
#46145000000
1!
1%
#46150000000
0!
0%
#46155000000
1!
1%
#46160000000
0!
0%
#46165000000
1!
1%
#46170000000
0!
0%
#46175000000
1!
1%
#46180000000
0!
0%
#46185000000
1!
1%
#46190000000
0!
0%
#46195000000
1!
1%
#46200000000
0!
0%
#46205000000
1!
1%
#46210000000
0!
0%
#46215000000
1!
1%
#46220000000
0!
0%
#46225000000
1!
1%
#46230000000
0!
0%
#46235000000
1!
1%
#46240000000
0!
0%
#46245000000
1!
1%
#46250000000
0!
0%
#46255000000
1!
1%
#46260000000
0!
0%
#46265000000
1!
1%
#46270000000
0!
0%
#46275000000
1!
1%
#46280000000
0!
0%
#46285000000
1!
1%
#46290000000
0!
0%
#46295000000
1!
1%
#46300000000
0!
0%
#46305000000
1!
1%
#46310000000
0!
0%
#46315000000
1!
1%
#46320000000
0!
0%
#46325000000
1!
1%
#46330000000
0!
0%
#46335000000
1!
1%
#46340000000
0!
0%
#46345000000
1!
1%
#46350000000
0!
0%
#46355000000
1!
1%
#46360000000
0!
0%
#46365000000
1!
1%
#46370000000
0!
0%
#46375000000
1!
1%
#46380000000
0!
0%
#46385000000
1!
1%
#46390000000
0!
0%
#46395000000
1!
1%
#46400000000
0!
0%
#46405000000
1!
1%
#46410000000
0!
0%
#46415000000
1!
1%
#46420000000
0!
0%
#46425000000
1!
1%
#46430000000
0!
0%
#46435000000
1!
1%
#46440000000
0!
0%
#46445000000
1!
1%
#46450000000
0!
0%
#46455000000
1!
1%
#46460000000
0!
0%
#46465000000
1!
1%
#46470000000
0!
0%
#46475000000
1!
1%
#46480000000
0!
0%
#46485000000
1!
1%
#46490000000
0!
0%
#46495000000
1!
1%
#46500000000
0!
0%
#46505000000
1!
1%
#46510000000
0!
0%
#46515000000
1!
1%
#46520000000
0!
0%
#46525000000
1!
1%
#46530000000
0!
0%
#46535000000
1!
1%
#46540000000
0!
0%
#46545000000
1!
1%
#46550000000
0!
0%
#46555000000
1!
1%
#46560000000
0!
0%
#46565000000
1!
1%
#46570000000
0!
0%
#46575000000
1!
1%
#46580000000
0!
0%
#46585000000
1!
1%
#46590000000
0!
0%
#46595000000
1!
1%
#46600000000
0!
0%
#46605000000
1!
1%
#46610000000
0!
0%
#46615000000
1!
1%
#46620000000
0!
0%
#46625000000
1!
1%
#46630000000
0!
0%
#46635000000
1!
1%
#46640000000
0!
0%
#46645000000
1!
1%
#46650000000
0!
0%
#46655000000
1!
1%
#46660000000
0!
0%
#46665000000
1!
1%
#46670000000
0!
0%
#46675000000
1!
1%
#46680000000
0!
0%
#46685000000
1!
1%
#46690000000
0!
0%
#46695000000
1!
1%
#46700000000
0!
0%
#46705000000
1!
1%
#46710000000
0!
0%
#46715000000
1!
1%
#46720000000
0!
0%
#46725000000
1!
1%
#46730000000
0!
0%
#46735000000
1!
1%
#46740000000
0!
0%
#46745000000
1!
1%
#46750000000
0!
0%
#46755000000
1!
1%
#46760000000
0!
0%
#46765000000
1!
1%
#46770000000
0!
0%
#46775000000
1!
1%
#46780000000
0!
0%
#46785000000
1!
1%
#46790000000
0!
0%
#46795000000
1!
1%
#46800000000
0!
0%
#46805000000
1!
1%
#46810000000
0!
0%
#46815000000
1!
1%
#46820000000
0!
0%
#46825000000
1!
1%
#46830000000
0!
0%
#46835000000
1!
1%
#46840000000
0!
0%
#46845000000
1!
1%
#46850000000
0!
0%
#46855000000
1!
1%
#46860000000
0!
0%
#46865000000
1!
1%
#46870000000
0!
0%
#46875000000
1!
1%
#46880000000
0!
0%
#46885000000
1!
1%
#46890000000
0!
0%
#46895000000
1!
1%
#46900000000
0!
0%
#46905000000
1!
1%
#46910000000
0!
0%
#46915000000
1!
1%
#46920000000
0!
0%
#46925000000
1!
1%
#46930000000
0!
0%
#46935000000
1!
1%
#46940000000
0!
0%
#46945000000
1!
1%
#46950000000
0!
0%
#46955000000
1!
1%
#46960000000
0!
0%
#46965000000
1!
1%
#46970000000
0!
0%
#46975000000
1!
1%
#46980000000
0!
0%
#46985000000
1!
1%
#46990000000
0!
0%
#46995000000
1!
1%
#47000000000
0!
0%
#47005000000
1!
1%
#47010000000
0!
0%
#47015000000
1!
1%
#47020000000
0!
0%
#47025000000
1!
1%
#47030000000
0!
0%
#47035000000
1!
1%
#47040000000
0!
0%
#47045000000
1!
1%
#47050000000
0!
0%
#47055000000
1!
1%
#47060000000
0!
0%
#47065000000
1!
1%
#47070000000
0!
0%
#47075000000
1!
1%
#47080000000
0!
0%
#47085000000
1!
1%
#47090000000
0!
0%
#47095000000
1!
1%
#47100000000
0!
0%
#47105000000
1!
1%
#47110000000
0!
0%
#47115000000
1!
1%
#47120000000
0!
0%
#47125000000
1!
1%
#47130000000
0!
0%
#47135000000
1!
1%
#47140000000
0!
0%
#47145000000
1!
1%
#47150000000
0!
0%
#47155000000
1!
1%
#47160000000
0!
0%
#47165000000
1!
1%
#47170000000
0!
0%
#47175000000
1!
1%
#47180000000
0!
0%
#47185000000
1!
1%
#47190000000
0!
0%
#47195000000
1!
1%
#47200000000
0!
0%
#47205000000
1!
1%
#47210000000
0!
0%
#47215000000
1!
1%
#47220000000
0!
0%
#47225000000
1!
1%
#47230000000
0!
0%
#47235000000
1!
1%
#47240000000
0!
0%
#47245000000
1!
1%
#47250000000
0!
0%
#47255000000
1!
1%
#47260000000
0!
0%
#47265000000
1!
1%
#47270000000
0!
0%
#47275000000
1!
1%
#47280000000
0!
0%
#47285000000
1!
1%
#47290000000
0!
0%
#47295000000
1!
1%
#47300000000
0!
0%
#47305000000
1!
1%
#47310000000
0!
0%
#47315000000
1!
1%
#47320000000
0!
0%
#47325000000
1!
1%
#47330000000
0!
0%
#47335000000
1!
1%
#47340000000
0!
0%
#47345000000
1!
1%
#47350000000
0!
0%
#47355000000
1!
1%
#47360000000
0!
0%
#47365000000
1!
1%
#47370000000
0!
0%
#47375000000
1!
1%
#47380000000
0!
0%
#47385000000
1!
1%
#47390000000
0!
0%
#47395000000
1!
1%
#47400000000
0!
0%
#47405000000
1!
1%
#47410000000
0!
0%
#47415000000
1!
1%
#47420000000
0!
0%
#47425000000
1!
1%
#47430000000
0!
0%
#47435000000
1!
1%
#47440000000
0!
0%
#47445000000
1!
1%
#47450000000
0!
0%
#47455000000
1!
1%
#47460000000
0!
0%
#47465000000
1!
1%
#47470000000
0!
0%
#47475000000
1!
1%
#47480000000
0!
0%
#47485000000
1!
1%
#47490000000
0!
0%
#47495000000
1!
1%
#47500000000
0!
0%
#47505000000
1!
1%
#47510000000
0!
0%
#47515000000
1!
1%
#47520000000
0!
0%
#47525000000
1!
1%
#47530000000
0!
0%
#47535000000
1!
1%
#47540000000
0!
0%
#47545000000
1!
1%
#47550000000
0!
0%
#47555000000
1!
1%
#47560000000
0!
0%
#47565000000
1!
1%
#47570000000
0!
0%
#47575000000
1!
1%
#47580000000
0!
0%
#47585000000
1!
1%
#47590000000
0!
0%
#47595000000
1!
1%
#47600000000
0!
0%
#47605000000
1!
1%
#47610000000
0!
0%
#47615000000
1!
1%
#47620000000
0!
0%
#47625000000
1!
1%
#47630000000
0!
0%
#47635000000
1!
1%
#47640000000
0!
0%
#47645000000
1!
1%
#47650000000
0!
0%
#47655000000
1!
1%
#47660000000
0!
0%
#47665000000
1!
1%
#47670000000
0!
0%
#47675000000
1!
1%
#47680000000
0!
0%
#47685000000
1!
1%
#47690000000
0!
0%
#47695000000
1!
1%
#47700000000
0!
0%
#47705000000
1!
1%
#47710000000
0!
0%
#47715000000
1!
1%
#47720000000
0!
0%
#47725000000
1!
1%
#47730000000
0!
0%
#47735000000
1!
1%
#47740000000
0!
0%
#47745000000
1!
1%
#47750000000
0!
0%
#47755000000
1!
1%
#47760000000
0!
0%
#47765000000
1!
1%
#47770000000
0!
0%
#47775000000
1!
1%
#47780000000
0!
0%
#47785000000
1!
1%
#47790000000
0!
0%
#47795000000
1!
1%
#47800000000
0!
0%
#47805000000
1!
1%
#47810000000
0!
0%
#47815000000
1!
1%
#47820000000
0!
0%
#47825000000
1!
1%
#47830000000
0!
0%
#47835000000
1!
1%
#47840000000
0!
0%
#47845000000
1!
1%
#47850000000
0!
0%
#47855000000
1!
1%
#47860000000
0!
0%
#47865000000
1!
1%
#47870000000
0!
0%
#47875000000
1!
1%
#47880000000
0!
0%
#47885000000
1!
1%
#47890000000
0!
0%
#47895000000
1!
1%
#47900000000
0!
0%
#47905000000
1!
1%
#47910000000
0!
0%
#47915000000
1!
1%
#47920000000
0!
0%
#47925000000
1!
1%
#47930000000
0!
0%
#47935000000
1!
1%
#47940000000
0!
0%
#47945000000
1!
1%
#47950000000
0!
0%
#47955000000
1!
1%
#47960000000
0!
0%
#47965000000
1!
1%
#47970000000
0!
0%
#47975000000
1!
1%
#47980000000
0!
0%
#47985000000
1!
1%
#47990000000
0!
0%
#47995000000
1!
1%
#48000000000
0!
0%
#48005000000
1!
1%
#48010000000
0!
0%
#48015000000
1!
1%
#48020000000
0!
0%
#48025000000
1!
1%
#48030000000
0!
0%
#48035000000
1!
1%
#48040000000
0!
0%
#48045000000
1!
1%
#48050000000
0!
0%
#48055000000
1!
1%
#48060000000
0!
0%
#48065000000
1!
1%
#48070000000
0!
0%
#48075000000
1!
1%
#48080000000
0!
0%
#48085000000
1!
1%
#48090000000
0!
0%
#48095000000
1!
1%
#48100000000
0!
0%
#48105000000
1!
1%
#48110000000
0!
0%
#48115000000
1!
1%
#48120000000
0!
0%
#48125000000
1!
1%
#48130000000
0!
0%
#48135000000
1!
1%
#48140000000
0!
0%
#48145000000
1!
1%
#48150000000
0!
0%
#48155000000
1!
1%
#48160000000
0!
0%
#48165000000
1!
1%
#48170000000
0!
0%
#48175000000
1!
1%
#48180000000
0!
0%
#48185000000
1!
1%
#48190000000
0!
0%
#48195000000
1!
1%
#48200000000
0!
0%
#48205000000
1!
1%
#48210000000
0!
0%
#48215000000
1!
1%
#48220000000
0!
0%
#48225000000
1!
1%
#48230000000
0!
0%
#48235000000
1!
1%
#48240000000
0!
0%
#48245000000
1!
1%
#48250000000
0!
0%
#48255000000
1!
1%
#48260000000
0!
0%
#48265000000
1!
1%
#48270000000
0!
0%
#48275000000
1!
1%
#48280000000
0!
0%
#48285000000
1!
1%
#48290000000
0!
0%
#48295000000
1!
1%
#48300000000
0!
0%
#48305000000
1!
1%
#48310000000
0!
0%
#48315000000
1!
1%
#48320000000
0!
0%
#48325000000
1!
1%
#48330000000
0!
0%
#48335000000
1!
1%
#48340000000
0!
0%
#48345000000
1!
1%
#48350000000
0!
0%
#48355000000
1!
1%
#48360000000
0!
0%
#48365000000
1!
1%
#48370000000
0!
0%
#48375000000
1!
1%
#48380000000
0!
0%
#48385000000
1!
1%
#48390000000
0!
0%
#48395000000
1!
1%
#48400000000
0!
0%
#48405000000
1!
1%
#48410000000
0!
0%
#48415000000
1!
1%
#48420000000
0!
0%
#48425000000
1!
1%
#48430000000
0!
0%
#48435000000
1!
1%
#48440000000
0!
0%
#48445000000
1!
1%
#48450000000
0!
0%
#48455000000
1!
1%
#48460000000
0!
0%
#48465000000
1!
1%
#48470000000
0!
0%
#48475000000
1!
1%
#48480000000
0!
0%
#48485000000
1!
1%
#48490000000
0!
0%
#48495000000
1!
1%
#48500000000
0!
0%
#48505000000
1!
1%
#48510000000
0!
0%
#48515000000
1!
1%
#48520000000
0!
0%
#48525000000
1!
1%
#48530000000
0!
0%
#48535000000
1!
1%
#48540000000
0!
0%
#48545000000
1!
1%
#48550000000
0!
0%
#48555000000
1!
1%
#48560000000
0!
0%
#48565000000
1!
1%
#48570000000
0!
0%
#48575000000
1!
1%
#48580000000
0!
0%
#48585000000
1!
1%
#48590000000
0!
0%
#48595000000
1!
1%
#48600000000
0!
0%
#48605000000
1!
1%
#48610000000
0!
0%
#48615000000
1!
1%
#48620000000
0!
0%
#48625000000
1!
1%
#48630000000
0!
0%
#48635000000
1!
1%
#48640000000
0!
0%
#48645000000
1!
1%
#48650000000
0!
0%
#48655000000
1!
1%
#48660000000
0!
0%
#48665000000
1!
1%
#48670000000
0!
0%
#48675000000
1!
1%
#48680000000
0!
0%
#48685000000
1!
1%
#48690000000
0!
0%
#48695000000
1!
1%
#48700000000
0!
0%
#48705000000
1!
1%
#48710000000
0!
0%
#48715000000
1!
1%
#48720000000
0!
0%
#48725000000
1!
1%
#48730000000
0!
0%
#48735000000
1!
1%
#48740000000
0!
0%
#48745000000
1!
1%
#48750000000
0!
0%
#48755000000
1!
1%
#48760000000
0!
0%
#48765000000
1!
1%
#48770000000
0!
0%
#48775000000
1!
1%
#48780000000
0!
0%
#48785000000
1!
1%
#48790000000
0!
0%
#48795000000
1!
1%
#48800000000
0!
0%
#48805000000
1!
1%
#48810000000
0!
0%
#48815000000
1!
1%
#48820000000
0!
0%
#48825000000
1!
1%
#48830000000
0!
0%
#48835000000
1!
1%
#48840000000
0!
0%
#48845000000
1!
1%
#48850000000
0!
0%
#48855000000
1!
1%
#48860000000
0!
0%
#48865000000
1!
1%
#48870000000
0!
0%
#48875000000
1!
1%
#48880000000
0!
0%
#48885000000
1!
1%
#48890000000
0!
0%
#48895000000
1!
1%
#48900000000
0!
0%
#48905000000
1!
1%
#48910000000
0!
0%
#48915000000
1!
1%
#48920000000
0!
0%
#48925000000
1!
1%
#48930000000
0!
0%
#48935000000
1!
1%
#48940000000
0!
0%
#48945000000
1!
1%
#48950000000
0!
0%
#48955000000
1!
1%
#48960000000
0!
0%
#48965000000
1!
1%
#48970000000
0!
0%
#48975000000
1!
1%
#48980000000
0!
0%
#48985000000
1!
1%
#48990000000
0!
0%
#48995000000
1!
1%
#49000000000
0!
0%
#49005000000
1!
1%
#49010000000
0!
0%
#49015000000
1!
1%
#49020000000
0!
0%
#49025000000
1!
1%
#49030000000
0!
0%
#49035000000
1!
1%
#49040000000
0!
0%
#49045000000
1!
1%
#49050000000
0!
0%
#49055000000
1!
1%
#49060000000
0!
0%
#49065000000
1!
1%
#49070000000
0!
0%
#49075000000
1!
1%
#49080000000
0!
0%
#49085000000
1!
1%
#49090000000
0!
0%
#49095000000
1!
1%
#49100000000
0!
0%
#49105000000
1!
1%
#49110000000
0!
0%
#49115000000
1!
1%
#49120000000
0!
0%
#49125000000
1!
1%
#49130000000
0!
0%
#49135000000
1!
1%
#49140000000
0!
0%
#49145000000
1!
1%
#49150000000
0!
0%
#49155000000
1!
1%
#49160000000
0!
0%
#49165000000
1!
1%
#49170000000
0!
0%
#49175000000
1!
1%
#49180000000
0!
0%
#49185000000
1!
1%
#49190000000
0!
0%
#49195000000
1!
1%
#49200000000
0!
0%
#49205000000
1!
1%
#49210000000
0!
0%
#49215000000
1!
1%
#49220000000
0!
0%
#49225000000
1!
1%
#49230000000
0!
0%
#49235000000
1!
1%
#49240000000
0!
0%
#49245000000
1!
1%
#49250000000
0!
0%
#49255000000
1!
1%
#49260000000
0!
0%
#49265000000
1!
1%
#49270000000
0!
0%
#49275000000
1!
1%
#49280000000
0!
0%
#49285000000
1!
1%
#49290000000
0!
0%
#49295000000
1!
1%
#49300000000
0!
0%
#49305000000
1!
1%
#49310000000
0!
0%
#49315000000
1!
1%
#49320000000
0!
0%
#49325000000
1!
1%
#49330000000
0!
0%
#49335000000
1!
1%
#49340000000
0!
0%
#49345000000
1!
1%
#49350000000
0!
0%
#49355000000
1!
1%
#49360000000
0!
0%
#49365000000
1!
1%
#49370000000
0!
0%
#49375000000
1!
1%
#49380000000
0!
0%
#49385000000
1!
1%
#49390000000
0!
0%
#49395000000
1!
1%
#49400000000
0!
0%
#49405000000
1!
1%
#49410000000
0!
0%
#49415000000
1!
1%
#49420000000
0!
0%
#49425000000
1!
1%
#49430000000
0!
0%
#49435000000
1!
1%
#49440000000
0!
0%
#49445000000
1!
1%
#49450000000
0!
0%
#49455000000
1!
1%
#49460000000
0!
0%
#49465000000
1!
1%
#49470000000
0!
0%
#49475000000
1!
1%
#49480000000
0!
0%
#49485000000
1!
1%
#49490000000
0!
0%
#49495000000
1!
1%
#49500000000
0!
0%
#49505000000
1!
1%
#49510000000
0!
0%
#49515000000
1!
1%
#49520000000
0!
0%
#49525000000
1!
1%
#49530000000
0!
0%
#49535000000
1!
1%
#49540000000
0!
0%
#49545000000
1!
1%
#49550000000
0!
0%
#49555000000
1!
1%
#49560000000
0!
0%
#49565000000
1!
1%
#49570000000
0!
0%
#49575000000
1!
1%
#49580000000
0!
0%
#49585000000
1!
1%
#49590000000
0!
0%
#49595000000
1!
1%
#49600000000
0!
0%
#49605000000
1!
1%
#49610000000
0!
0%
#49615000000
1!
1%
#49620000000
0!
0%
#49625000000
1!
1%
#49630000000
0!
0%
#49635000000
1!
1%
#49640000000
0!
0%
#49645000000
1!
1%
#49650000000
0!
0%
#49655000000
1!
1%
#49660000000
0!
0%
#49665000000
1!
1%
#49670000000
0!
0%
#49675000000
1!
1%
#49680000000
0!
0%
#49685000000
1!
1%
#49690000000
0!
0%
#49695000000
1!
1%
#49700000000
0!
0%
#49705000000
1!
1%
#49710000000
0!
0%
#49715000000
1!
1%
#49720000000
0!
0%
#49725000000
1!
1%
#49730000000
0!
0%
#49735000000
1!
1%
#49740000000
0!
0%
#49745000000
1!
1%
#49750000000
0!
0%
#49755000000
1!
1%
#49760000000
0!
0%
#49765000000
1!
1%
#49770000000
0!
0%
#49775000000
1!
1%
#49780000000
0!
0%
#49785000000
1!
1%
#49790000000
0!
0%
#49795000000
1!
1%
#49800000000
0!
0%
#49805000000
1!
1%
#49810000000
0!
0%
#49815000000
1!
1%
#49820000000
0!
0%
#49825000000
1!
1%
#49830000000
0!
0%
#49835000000
1!
1%
#49840000000
0!
0%
#49845000000
1!
1%
#49850000000
0!
0%
#49855000000
1!
1%
#49860000000
0!
0%
#49865000000
1!
1%
#49870000000
0!
0%
#49875000000
1!
1%
#49880000000
0!
0%
#49885000000
1!
1%
#49890000000
0!
0%
#49895000000
1!
1%
#49900000000
0!
0%
#49905000000
1!
1%
#49910000000
0!
0%
#49915000000
1!
1%
#49920000000
0!
0%
#49925000000
1!
1%
#49930000000
0!
0%
#49935000000
1!
1%
#49940000000
0!
0%
#49945000000
1!
1%
#49950000000
0!
0%
#49955000000
1!
1%
#49960000000
0!
0%
#49965000000
1!
1%
#49970000000
0!
0%
#49975000000
1!
1%
#49980000000
0!
0%
#49985000000
1!
1%
#49990000000
0!
0%
#49995000000
1!
1%
#50000000000
0!
0%
#50005000000
1!
1%
#50010000000
0!
0%
#50015000000
1!
1%
#50020000000
0!
0%
#50025000000
1!
1%
#50030000000
0!
0%
#50035000000
1!
1%
#50040000000
0!
0%
#50045000000
1!
1%
#50050000000
0!
0%
#50055000000
1!
1%
#50060000000
0!
0%
#50065000000
1!
1%
#50070000000
0!
0%
#50075000000
1!
1%
#50080000000
0!
0%
#50085000000
1!
1%
#50090000000
0!
0%
#50095000000
1!
1%
#50100000000
0!
0%
#50105000000
1!
1%
#50110000000
0!
0%
#50115000000
1!
1%
#50120000000
0!
0%
#50125000000
1!
1%
#50130000000
0!
0%
#50135000000
1!
1%
#50140000000
0!
0%
#50145000000
1!
1%
#50150000000
0!
0%
#50155000000
1!
1%
#50160000000
0!
0%
#50165000000
1!
1%
#50170000000
0!
0%
#50175000000
1!
1%
#50180000000
0!
0%
#50185000000
1!
1%
#50190000000
0!
0%
#50195000000
1!
1%
#50200000000
0!
0%
#50205000000
1!
1%
#50210000000
0!
0%
#50215000000
1!
1%
#50220000000
0!
0%
#50225000000
1!
1%
#50230000000
0!
0%
#50235000000
1!
1%
#50240000000
0!
0%
#50245000000
1!
1%
#50250000000
0!
0%
#50255000000
1!
1%
#50260000000
0!
0%
#50265000000
1!
1%
#50270000000
0!
0%
#50275000000
1!
1%
#50280000000
0!
0%
#50285000000
1!
1%
#50290000000
0!
0%
#50295000000
1!
1%
#50300000000
0!
0%
#50305000000
1!
1%
#50310000000
0!
0%
#50315000000
1!
1%
#50320000000
0!
0%
#50325000000
1!
1%
#50330000000
0!
0%
#50335000000
1!
1%
#50340000000
0!
0%
#50345000000
1!
1%
#50350000000
0!
0%
#50355000000
1!
1%
#50360000000
0!
0%
#50365000000
1!
1%
#50370000000
0!
0%
#50375000000
1!
1%
#50380000000
0!
0%
#50385000000
1!
1%
#50390000000
0!
0%
#50395000000
1!
1%
#50400000000
0!
0%
#50405000000
1!
1%
#50410000000
0!
0%
#50415000000
1!
1%
#50420000000
0!
0%
#50425000000
1!
1%
#50430000000
0!
0%
#50435000000
1!
1%
#50440000000
0!
0%
#50445000000
1!
1%
#50450000000
0!
0%
#50455000000
1!
1%
#50460000000
0!
0%
#50465000000
1!
1%
#50470000000
0!
0%
#50475000000
1!
1%
#50480000000
0!
0%
#50485000000
1!
1%
#50490000000
0!
0%
#50495000000
1!
1%
#50500000000
0!
0%
#50505000000
1!
1%
#50510000000
0!
0%
#50515000000
1!
1%
#50520000000
0!
0%
#50525000000
1!
1%
#50530000000
0!
0%
#50535000000
1!
1%
#50540000000
0!
0%
#50545000000
1!
1%
#50550000000
0!
0%
#50555000000
1!
1%
#50560000000
0!
0%
#50565000000
1!
1%
#50570000000
0!
0%
#50575000000
1!
1%
#50580000000
0!
0%
#50585000000
1!
1%
#50590000000
0!
0%
#50595000000
1!
1%
#50600000000
0!
0%
#50605000000
1!
1%
#50610000000
0!
0%
#50615000000
1!
1%
#50620000000
0!
0%
#50625000000
1!
1%
#50630000000
0!
0%
#50635000000
1!
1%
#50640000000
0!
0%
#50645000000
1!
1%
#50650000000
0!
0%
#50655000000
1!
1%
#50660000000
0!
0%
#50665000000
1!
1%
#50670000000
0!
0%
#50675000000
1!
1%
#50680000000
0!
0%
#50685000000
1!
1%
#50690000000
0!
0%
#50695000000
1!
1%
#50700000000
0!
0%
#50705000000
1!
1%
#50710000000
0!
0%
#50715000000
1!
1%
#50720000000
0!
0%
#50725000000
1!
1%
#50730000000
0!
0%
#50735000000
1!
1%
#50740000000
0!
0%
#50745000000
1!
1%
#50750000000
0!
0%
#50755000000
1!
1%
#50760000000
0!
0%
#50765000000
1!
1%
#50770000000
0!
0%
#50775000000
1!
1%
#50780000000
0!
0%
#50785000000
1!
1%
#50790000000
0!
0%
#50795000000
1!
1%
#50800000000
0!
0%
#50805000000
1!
1%
#50810000000
0!
0%
#50815000000
1!
1%
#50820000000
0!
0%
#50825000000
1!
1%
#50830000000
0!
0%
#50835000000
1!
1%
#50840000000
0!
0%
#50845000000
1!
1%
#50850000000
0!
0%
#50855000000
1!
1%
#50860000000
0!
0%
#50865000000
1!
1%
#50870000000
0!
0%
#50875000000
1!
1%
#50880000000
0!
0%
#50885000000
1!
1%
#50890000000
0!
0%
#50895000000
1!
1%
#50900000000
0!
0%
#50905000000
1!
1%
#50910000000
0!
0%
#50915000000
1!
1%
#50920000000
0!
0%
#50925000000
1!
1%
#50930000000
0!
0%
#50935000000
1!
1%
#50940000000
0!
0%
#50945000000
1!
1%
#50950000000
0!
0%
#50955000000
1!
1%
#50960000000
0!
0%
#50965000000
1!
1%
#50970000000
0!
0%
#50975000000
1!
1%
#50980000000
0!
0%
#50985000000
1!
1%
#50990000000
0!
0%
#50995000000
1!
1%
#51000000000
0!
0%
#51005000000
1!
1%
#51010000000
0!
0%
#51015000000
1!
1%
#51020000000
0!
0%
#51025000000
1!
1%
#51030000000
0!
0%
#51035000000
1!
1%
#51040000000
0!
0%
#51045000000
1!
1%
#51050000000
0!
0%
#51055000000
1!
1%
#51060000000
0!
0%
#51065000000
1!
1%
#51070000000
0!
0%
#51075000000
1!
1%
#51080000000
0!
0%
#51085000000
1!
1%
#51090000000
0!
0%
#51095000000
1!
1%
#51100000000
0!
0%
#51105000000
1!
1%
#51110000000
0!
0%
#51115000000
1!
1%
#51120000000
0!
0%
#51125000000
1!
1%
#51130000000
0!
0%
#51135000000
1!
1%
#51140000000
0!
0%
#51145000000
1!
1%
#51150000000
0!
0%
#51155000000
1!
1%
#51160000000
0!
0%
#51165000000
1!
1%
#51170000000
0!
0%
#51175000000
1!
1%
#51180000000
0!
0%
#51185000000
1!
1%
#51190000000
0!
0%
#51195000000
1!
1%
#51200000000
0!
0%
#51205000000
1!
1%
#51210000000
0!
0%
#51215000000
1!
1%
#51220000000
0!
0%
#51225000000
1!
1%
#51230000000
0!
0%
#51235000000
1!
1%
#51240000000
0!
0%
#51245000000
1!
1%
#51250000000
0!
0%
#51255000000
1!
1%
#51260000000
0!
0%
#51265000000
1!
1%
#51270000000
0!
0%
#51275000000
1!
1%
#51280000000
0!
0%
#51285000000
1!
1%
#51290000000
0!
0%
#51295000000
1!
1%
#51300000000
0!
0%
#51305000000
1!
1%
#51310000000
0!
0%
#51315000000
1!
1%
#51320000000
0!
0%
#51325000000
1!
1%
#51330000000
0!
0%
#51335000000
1!
1%
#51340000000
0!
0%
#51345000000
1!
1%
#51350000000
0!
0%
#51355000000
1!
1%
#51360000000
0!
0%
#51365000000
1!
1%
#51370000000
0!
0%
#51375000000
1!
1%
#51380000000
0!
0%
#51385000000
1!
1%
#51390000000
0!
0%
#51395000000
1!
1%
#51400000000
0!
0%
#51405000000
1!
1%
#51410000000
0!
0%
#51415000000
1!
1%
#51420000000
0!
0%
#51425000000
1!
1%
#51430000000
0!
0%
#51435000000
1!
1%
#51440000000
0!
0%
#51445000000
1!
1%
#51450000000
0!
0%
#51455000000
1!
1%
#51460000000
0!
0%
#51465000000
1!
1%
#51470000000
0!
0%
#51475000000
1!
1%
#51480000000
0!
0%
#51485000000
1!
1%
#51490000000
0!
0%
#51495000000
1!
1%
#51500000000
0!
0%
#51505000000
1!
1%
#51510000000
0!
0%
#51515000000
1!
1%
#51520000000
0!
0%
#51525000000
1!
1%
#51530000000
0!
0%
#51535000000
1!
1%
#51540000000
0!
0%
#51545000000
1!
1%
#51550000000
0!
0%
#51555000000
1!
1%
#51560000000
0!
0%
#51565000000
1!
1%
#51570000000
0!
0%
#51575000000
1!
1%
#51580000000
0!
0%
#51585000000
1!
1%
#51590000000
0!
0%
#51595000000
1!
1%
#51600000000
0!
0%
#51605000000
1!
1%
#51610000000
0!
0%
#51615000000
1!
1%
#51620000000
0!
0%
#51625000000
1!
1%
#51630000000
0!
0%
#51635000000
1!
1%
#51640000000
0!
0%
#51645000000
1!
1%
#51650000000
0!
0%
#51655000000
1!
1%
#51660000000
0!
0%
#51665000000
1!
1%
#51670000000
0!
0%
#51675000000
1!
1%
#51680000000
0!
0%
#51685000000
1!
1%
#51690000000
0!
0%
#51695000000
1!
1%
#51700000000
0!
0%
#51705000000
1!
1%
#51710000000
0!
0%
#51715000000
1!
1%
#51720000000
0!
0%
#51725000000
1!
1%
#51730000000
0!
0%
#51735000000
1!
1%
#51740000000
0!
0%
#51745000000
1!
1%
#51750000000
0!
0%
#51755000000
1!
1%
#51760000000
0!
0%
#51765000000
1!
1%
#51770000000
0!
0%
#51775000000
1!
1%
#51780000000
0!
0%
#51785000000
1!
1%
#51790000000
0!
0%
#51795000000
1!
1%
#51800000000
0!
0%
#51805000000
1!
1%
#51810000000
0!
0%
#51815000000
1!
1%
#51820000000
0!
0%
#51825000000
1!
1%
#51830000000
0!
0%
#51835000000
1!
1%
#51840000000
0!
0%
#51845000000
1!
1%
#51850000000
0!
0%
#51855000000
1!
1%
#51860000000
0!
0%
#51865000000
1!
1%
#51870000000
0!
0%
#51875000000
1!
1%
#51880000000
0!
0%
#51885000000
1!
1%
#51890000000
0!
0%
#51895000000
1!
1%
#51900000000
0!
0%
#51905000000
1!
1%
#51910000000
0!
0%
#51915000000
1!
1%
#51920000000
0!
0%
#51925000000
1!
1%
#51930000000
0!
0%
#51935000000
1!
1%
#51940000000
0!
0%
#51945000000
1!
1%
#51950000000
0!
0%
#51955000000
1!
1%
#51960000000
0!
0%
#51965000000
1!
1%
#51970000000
0!
0%
#51975000000
1!
1%
#51980000000
0!
0%
#51985000000
1!
1%
#51990000000
0!
0%
#51995000000
1!
1%
#52000000000
0!
0%
#52005000000
1!
1%
#52010000000
0!
0%
#52015000000
1!
1%
#52020000000
0!
0%
#52025000000
1!
1%
#52030000000
0!
0%
#52035000000
1!
1%
#52040000000
0!
0%
#52045000000
1!
1%
#52050000000
0!
0%
#52055000000
1!
1%
#52060000000
0!
0%
#52065000000
1!
1%
#52070000000
0!
0%
#52075000000
1!
1%
#52080000000
0!
0%
#52085000000
1!
1%
#52090000000
0!
0%
#52095000000
1!
1%
#52100000000
0!
0%
#52105000000
1!
1%
#52110000000
0!
0%
#52115000000
1!
1%
#52120000000
0!
0%
#52125000000
1!
1%
#52130000000
0!
0%
#52135000000
1!
1%
#52140000000
0!
0%
#52145000000
1!
1%
#52150000000
0!
0%
#52155000000
1!
1%
#52160000000
0!
0%
#52165000000
1!
1%
#52170000000
0!
0%
#52175000000
1!
1%
#52180000000
0!
0%
#52185000000
1!
1%
#52190000000
0!
0%
#52195000000
1!
1%
#52200000000
0!
0%
#52205000000
1!
1%
#52210000000
0!
0%
#52215000000
1!
1%
#52220000000
0!
0%
#52225000000
1!
1%
#52230000000
0!
0%
#52235000000
1!
1%
#52240000000
0!
0%
#52245000000
1!
1%
#52250000000
0!
0%
#52255000000
1!
1%
#52260000000
0!
0%
#52265000000
1!
1%
#52270000000
0!
0%
#52275000000
1!
1%
#52280000000
0!
0%
#52285000000
1!
1%
#52290000000
0!
0%
#52295000000
1!
1%
#52300000000
0!
0%
#52305000000
1!
1%
#52310000000
0!
0%
#52315000000
1!
1%
#52320000000
0!
0%
#52325000000
1!
1%
#52330000000
0!
0%
#52335000000
1!
1%
#52340000000
0!
0%
#52345000000
1!
1%
#52350000000
0!
0%
#52355000000
1!
1%
#52360000000
0!
0%
#52365000000
1!
1%
#52370000000
0!
0%
#52375000000
1!
1%
#52380000000
0!
0%
#52385000000
1!
1%
#52390000000
0!
0%
#52395000000
1!
1%
#52400000000
0!
0%
#52405000000
1!
1%
#52410000000
0!
0%
#52415000000
1!
1%
#52420000000
0!
0%
#52425000000
1!
1%
#52430000000
0!
0%
#52435000000
1!
1%
#52440000000
0!
0%
#52445000000
1!
1%
#52450000000
0!
0%
#52455000000
1!
1%
#52460000000
0!
0%
#52465000000
1!
1%
#52470000000
0!
0%
#52475000000
1!
1%
#52480000000
0!
0%
#52485000000
1!
1%
#52490000000
0!
0%
#52495000000
1!
1%
#52500000000
0!
0%
#52505000000
1!
1%
#52510000000
0!
0%
#52515000000
1!
1%
#52520000000
0!
0%
#52525000000
1!
1%
#52530000000
0!
0%
#52535000000
1!
1%
#52540000000
0!
0%
#52545000000
1!
1%
#52550000000
0!
0%
#52555000000
1!
1%
#52560000000
0!
0%
#52565000000
1!
1%
#52570000000
0!
0%
#52575000000
1!
1%
#52580000000
0!
0%
#52585000000
1!
1%
#52590000000
0!
0%
#52595000000
1!
1%
#52600000000
0!
0%
#52605000000
1!
1%
#52610000000
0!
0%
#52615000000
1!
1%
#52620000000
0!
0%
#52625000000
1!
1%
#52630000000
0!
0%
#52635000000
1!
1%
#52640000000
0!
0%
#52645000000
1!
1%
#52650000000
0!
0%
#52655000000
1!
1%
#52660000000
0!
0%
#52665000000
1!
1%
#52670000000
0!
0%
#52675000000
1!
1%
#52680000000
0!
0%
#52685000000
1!
1%
#52690000000
0!
0%
#52695000000
1!
1%
#52700000000
0!
0%
#52705000000
1!
1%
#52710000000
0!
0%
#52715000000
1!
1%
#52720000000
0!
0%
#52725000000
1!
1%
#52730000000
0!
0%
#52735000000
1!
1%
#52740000000
0!
0%
#52745000000
1!
1%
#52750000000
0!
0%
#52755000000
1!
1%
#52760000000
0!
0%
#52765000000
1!
1%
#52770000000
0!
0%
#52775000000
1!
1%
#52780000000
0!
0%
#52785000000
1!
1%
#52790000000
0!
0%
#52795000000
1!
1%
#52800000000
0!
0%
#52805000000
1!
1%
#52810000000
0!
0%
#52815000000
1!
1%
#52820000000
0!
0%
#52825000000
1!
1%
#52830000000
0!
0%
#52835000000
1!
1%
#52840000000
0!
0%
#52845000000
1!
1%
#52850000000
0!
0%
#52855000000
1!
1%
#52860000000
0!
0%
#52865000000
1!
1%
#52870000000
0!
0%
#52875000000
1!
1%
#52880000000
0!
0%
#52885000000
1!
1%
#52890000000
0!
0%
#52895000000
1!
1%
#52900000000
0!
0%
#52905000000
1!
1%
#52910000000
0!
0%
#52915000000
1!
1%
#52920000000
0!
0%
#52925000000
1!
1%
#52930000000
0!
0%
#52935000000
1!
1%
#52940000000
0!
0%
#52945000000
1!
1%
#52950000000
0!
0%
#52955000000
1!
1%
#52960000000
0!
0%
#52965000000
1!
1%
#52970000000
0!
0%
#52975000000
1!
1%
#52980000000
0!
0%
#52985000000
1!
1%
#52990000000
0!
0%
#52995000000
1!
1%
#53000000000
0!
0%
#53005000000
1!
1%
#53010000000
0!
0%
#53015000000
1!
1%
#53020000000
0!
0%
#53025000000
1!
1%
#53030000000
0!
0%
#53035000000
1!
1%
#53040000000
0!
0%
#53045000000
1!
1%
#53050000000
0!
0%
#53055000000
1!
1%
#53060000000
0!
0%
#53065000000
1!
1%
#53070000000
0!
0%
#53075000000
1!
1%
#53080000000
0!
0%
#53085000000
1!
1%
#53090000000
0!
0%
#53095000000
1!
1%
#53100000000
0!
0%
#53105000000
1!
1%
#53110000000
0!
0%
#53115000000
1!
1%
#53120000000
0!
0%
#53125000000
1!
1%
#53130000000
0!
0%
#53135000000
1!
1%
#53140000000
0!
0%
#53145000000
1!
1%
#53150000000
0!
0%
#53155000000
1!
1%
#53160000000
0!
0%
#53165000000
1!
1%
#53170000000
0!
0%
#53175000000
1!
1%
#53180000000
0!
0%
#53185000000
1!
1%
#53190000000
0!
0%
#53195000000
1!
1%
#53200000000
0!
0%
#53205000000
1!
1%
#53210000000
0!
0%
#53215000000
1!
1%
#53220000000
0!
0%
#53225000000
1!
1%
#53230000000
0!
0%
#53235000000
1!
1%
#53240000000
0!
0%
#53245000000
1!
1%
#53250000000
0!
0%
#53255000000
1!
1%
#53260000000
0!
0%
#53265000000
1!
1%
#53270000000
0!
0%
#53275000000
1!
1%
#53280000000
0!
0%
#53285000000
1!
1%
#53290000000
0!
0%
#53295000000
1!
1%
#53300000000
0!
0%
#53305000000
1!
1%
#53310000000
0!
0%
#53315000000
1!
1%
#53320000000
0!
0%
#53325000000
1!
1%
#53330000000
0!
0%
#53335000000
1!
1%
#53340000000
0!
0%
#53345000000
1!
1%
#53350000000
0!
0%
#53355000000
1!
1%
#53360000000
0!
0%
#53365000000
1!
1%
#53370000000
0!
0%
#53375000000
1!
1%
#53380000000
0!
0%
#53385000000
1!
1%
#53390000000
0!
0%
#53395000000
1!
1%
#53400000000
0!
0%
#53405000000
1!
1%
#53410000000
0!
0%
#53415000000
1!
1%
#53420000000
0!
0%
#53425000000
1!
1%
#53430000000
0!
0%
#53435000000
1!
1%
#53440000000
0!
0%
#53445000000
1!
1%
#53450000000
0!
0%
#53455000000
1!
1%
#53460000000
0!
0%
#53465000000
1!
1%
#53470000000
0!
0%
#53475000000
1!
1%
#53480000000
0!
0%
#53485000000
1!
1%
#53490000000
0!
0%
#53495000000
1!
1%
#53500000000
0!
0%
#53505000000
1!
1%
#53510000000
0!
0%
#53515000000
1!
1%
#53520000000
0!
0%
#53525000000
1!
1%
#53530000000
0!
0%
#53535000000
1!
1%
#53540000000
0!
0%
#53545000000
1!
1%
#53550000000
0!
0%
#53555000000
1!
1%
#53560000000
0!
0%
#53565000000
1!
1%
#53570000000
0!
0%
#53575000000
1!
1%
#53580000000
0!
0%
#53585000000
1!
1%
#53590000000
0!
0%
#53595000000
1!
1%
#53600000000
0!
0%
#53605000000
1!
1%
#53610000000
0!
0%
#53615000000
1!
1%
#53620000000
0!
0%
#53625000000
1!
1%
#53630000000
0!
0%
#53635000000
1!
1%
#53640000000
0!
0%
#53645000000
1!
1%
#53650000000
0!
0%
#53655000000
1!
1%
#53660000000
0!
0%
#53665000000
1!
1%
#53670000000
0!
0%
#53675000000
1!
1%
#53680000000
0!
0%
#53685000000
1!
1%
#53690000000
0!
0%
#53695000000
1!
1%
#53700000000
0!
0%
#53705000000
1!
1%
#53710000000
0!
0%
#53715000000
1!
1%
#53720000000
0!
0%
#53725000000
1!
1%
#53730000000
0!
0%
#53735000000
1!
1%
#53740000000
0!
0%
#53745000000
1!
1%
#53750000000
0!
0%
#53755000000
1!
1%
#53760000000
0!
0%
#53765000000
1!
1%
#53770000000
0!
0%
#53775000000
1!
1%
#53780000000
0!
0%
#53785000000
1!
1%
#53790000000
0!
0%
#53795000000
1!
1%
#53800000000
0!
0%
#53805000000
1!
1%
#53810000000
0!
0%
#53815000000
1!
1%
#53820000000
0!
0%
#53825000000
1!
1%
#53830000000
0!
0%
#53835000000
1!
1%
#53840000000
0!
0%
#53845000000
1!
1%
#53850000000
0!
0%
#53855000000
1!
1%
#53860000000
0!
0%
#53865000000
1!
1%
#53870000000
0!
0%
#53875000000
1!
1%
#53880000000
0!
0%
#53885000000
1!
1%
#53890000000
0!
0%
#53895000000
1!
1%
#53900000000
0!
0%
#53905000000
1!
1%
#53910000000
0!
0%
#53915000000
1!
1%
#53920000000
0!
0%
#53925000000
1!
1%
#53930000000
0!
0%
#53935000000
1!
1%
#53940000000
0!
0%
#53945000000
1!
1%
#53950000000
0!
0%
#53955000000
1!
1%
#53960000000
0!
0%
#53965000000
1!
1%
#53970000000
0!
0%
#53975000000
1!
1%
#53980000000
0!
0%
#53985000000
1!
1%
#53990000000
0!
0%
#53995000000
1!
1%
#54000000000
0!
0%
#54005000000
1!
1%
#54010000000
0!
0%
#54015000000
1!
1%
#54020000000
0!
0%
#54025000000
1!
1%
#54030000000
0!
0%
#54035000000
1!
1%
#54040000000
0!
0%
#54045000000
1!
1%
#54050000000
0!
0%
#54055000000
1!
1%
#54060000000
0!
0%
#54065000000
1!
1%
#54070000000
0!
0%
#54075000000
1!
1%
#54080000000
0!
0%
#54085000000
1!
1%
#54090000000
0!
0%
#54095000000
1!
1%
#54100000000
0!
0%
#54105000000
1!
1%
#54110000000
0!
0%
#54115000000
1!
1%
#54120000000
0!
0%
#54125000000
1!
1%
#54130000000
0!
0%
#54135000000
1!
1%
#54140000000
0!
0%
#54145000000
1!
1%
#54150000000
0!
0%
#54155000000
1!
1%
#54160000000
0!
0%
#54165000000
1!
1%
#54170000000
0!
0%
#54175000000
1!
1%
#54180000000
0!
0%
#54185000000
1!
1%
#54190000000
0!
0%
#54195000000
1!
1%
#54200000000
0!
0%
#54205000000
1!
1%
#54210000000
0!
0%
#54215000000
1!
1%
#54220000000
0!
0%
#54225000000
1!
1%
#54230000000
0!
0%
#54235000000
1!
1%
#54240000000
0!
0%
#54245000000
1!
1%
#54250000000
0!
0%
#54255000000
1!
1%
#54260000000
0!
0%
#54265000000
1!
1%
#54270000000
0!
0%
#54275000000
1!
1%
#54280000000
0!
0%
#54285000000
1!
1%
#54290000000
0!
0%
#54295000000
1!
1%
#54300000000
0!
0%
#54305000000
1!
1%
#54310000000
0!
0%
#54315000000
1!
1%
#54320000000
0!
0%
#54325000000
1!
1%
#54330000000
0!
0%
#54335000000
1!
1%
#54340000000
0!
0%
#54345000000
1!
1%
#54350000000
0!
0%
#54355000000
1!
1%
#54360000000
0!
0%
#54365000000
1!
1%
#54370000000
0!
0%
#54375000000
1!
1%
#54380000000
0!
0%
#54385000000
1!
1%
#54390000000
0!
0%
#54395000000
1!
1%
#54400000000
0!
0%
#54405000000
1!
1%
#54410000000
0!
0%
#54415000000
1!
1%
#54420000000
0!
0%
#54425000000
1!
1%
#54430000000
0!
0%
#54435000000
1!
1%
#54440000000
0!
0%
#54445000000
1!
1%
#54450000000
0!
0%
#54455000000
1!
1%
#54460000000
0!
0%
#54465000000
1!
1%
#54470000000
0!
0%
#54475000000
1!
1%
#54480000000
0!
0%
#54485000000
1!
1%
#54490000000
0!
0%
#54495000000
1!
1%
#54500000000
0!
0%
#54505000000
1!
1%
#54510000000
0!
0%
#54515000000
1!
1%
#54520000000
0!
0%
#54525000000
1!
1%
#54530000000
0!
0%
#54535000000
1!
1%
#54540000000
0!
0%
#54545000000
1!
1%
#54550000000
0!
0%
#54555000000
1!
1%
#54560000000
0!
0%
#54565000000
1!
1%
#54570000000
0!
0%
#54575000000
1!
1%
#54580000000
0!
0%
#54585000000
1!
1%
#54590000000
0!
0%
#54595000000
1!
1%
#54600000000
0!
0%
#54605000000
1!
1%
#54610000000
0!
0%
#54615000000
1!
1%
#54620000000
0!
0%
#54625000000
1!
1%
#54630000000
0!
0%
#54635000000
1!
1%
#54640000000
0!
0%
#54645000000
1!
1%
#54650000000
0!
0%
#54655000000
1!
1%
#54660000000
0!
0%
#54665000000
1!
1%
#54670000000
0!
0%
#54675000000
1!
1%
#54680000000
0!
0%
#54685000000
1!
1%
#54690000000
0!
0%
#54695000000
1!
1%
#54700000000
0!
0%
#54705000000
1!
1%
#54710000000
0!
0%
#54715000000
1!
1%
#54720000000
0!
0%
#54725000000
1!
1%
#54730000000
0!
0%
#54735000000
1!
1%
#54740000000
0!
0%
#54745000000
1!
1%
#54750000000
0!
0%
#54755000000
1!
1%
#54760000000
0!
0%
#54765000000
1!
1%
#54770000000
0!
0%
#54775000000
1!
1%
#54780000000
0!
0%
#54785000000
1!
1%
#54790000000
0!
0%
#54795000000
1!
1%
#54800000000
0!
0%
#54805000000
1!
1%
#54810000000
0!
0%
#54815000000
1!
1%
#54820000000
0!
0%
#54825000000
1!
1%
#54830000000
0!
0%
#54835000000
1!
1%
#54840000000
0!
0%
#54845000000
1!
1%
#54850000000
0!
0%
#54855000000
1!
1%
#54860000000
0!
0%
#54865000000
1!
1%
#54870000000
0!
0%
#54875000000
1!
1%
#54880000000
0!
0%
#54885000000
1!
1%
#54890000000
0!
0%
#54895000000
1!
1%
#54900000000
0!
0%
#54905000000
1!
1%
#54910000000
0!
0%
#54915000000
1!
1%
#54920000000
0!
0%
#54925000000
1!
1%
#54930000000
0!
0%
#54935000000
1!
1%
#54940000000
0!
0%
#54945000000
1!
1%
#54950000000
0!
0%
#54955000000
1!
1%
#54960000000
0!
0%
#54965000000
1!
1%
#54970000000
0!
0%
#54975000000
1!
1%
#54980000000
0!
0%
#54985000000
1!
1%
#54990000000
0!
0%
#54995000000
1!
1%
#55000000000
0!
0%
#55005000000
1!
1%
#55010000000
0!
0%
#55015000000
1!
1%
#55020000000
0!
0%
#55025000000
1!
1%
#55030000000
0!
0%
#55035000000
1!
1%
#55040000000
0!
0%
#55045000000
1!
1%
#55050000000
0!
0%
#55055000000
1!
1%
#55060000000
0!
0%
#55065000000
1!
1%
#55070000000
0!
0%
#55075000000
1!
1%
#55080000000
0!
0%
#55085000000
1!
1%
#55090000000
0!
0%
#55095000000
1!
1%
#55100000000
0!
0%
#55105000000
1!
1%
#55110000000
0!
0%
#55115000000
1!
1%
#55120000000
0!
0%
#55125000000
1!
1%
#55130000000
0!
0%
#55135000000
1!
1%
#55140000000
0!
0%
#55145000000
1!
1%
#55150000000
0!
0%
#55155000000
1!
1%
#55160000000
0!
0%
#55165000000
1!
1%
#55170000000
0!
0%
#55175000000
1!
1%
#55180000000
0!
0%
#55185000000
1!
1%
#55190000000
0!
0%
#55195000000
1!
1%
#55200000000
0!
0%
#55205000000
1!
1%
#55210000000
0!
0%
#55215000000
1!
1%
#55220000000
0!
0%
#55225000000
1!
1%
#55230000000
0!
0%
#55235000000
1!
1%
#55240000000
0!
0%
#55245000000
1!
1%
#55250000000
0!
0%
#55255000000
1!
1%
#55260000000
0!
0%
#55265000000
1!
1%
#55270000000
0!
0%
#55275000000
1!
1%
#55280000000
0!
0%
#55285000000
1!
1%
#55290000000
0!
0%
#55295000000
1!
1%
#55300000000
0!
0%
#55305000000
1!
1%
#55310000000
0!
0%
#55315000000
1!
1%
#55320000000
0!
0%
#55325000000
1!
1%
#55330000000
0!
0%
#55335000000
1!
1%
#55340000000
0!
0%
#55345000000
1!
1%
#55350000000
0!
0%
#55355000000
1!
1%
#55360000000
0!
0%
#55365000000
1!
1%
#55370000000
0!
0%
#55375000000
1!
1%
#55380000000
0!
0%
#55385000000
1!
1%
#55390000000
0!
0%
#55395000000
1!
1%
#55400000000
0!
0%
#55405000000
1!
1%
#55410000000
0!
0%
#55415000000
1!
1%
#55420000000
0!
0%
#55425000000
1!
1%
#55430000000
0!
0%
#55435000000
1!
1%
#55440000000
0!
0%
#55445000000
1!
1%
#55450000000
0!
0%
#55455000000
1!
1%
#55460000000
0!
0%
#55465000000
1!
1%
#55470000000
0!
0%
#55475000000
1!
1%
#55480000000
0!
0%
#55485000000
1!
1%
#55490000000
0!
0%
#55495000000
1!
1%
#55500000000
0!
0%
#55505000000
1!
1%
#55510000000
0!
0%
#55515000000
1!
1%
#55520000000
0!
0%
#55525000000
1!
1%
#55530000000
0!
0%
#55535000000
1!
1%
#55540000000
0!
0%
#55545000000
1!
1%
#55550000000
0!
0%
#55555000000
1!
1%
#55560000000
0!
0%
#55565000000
1!
1%
#55570000000
0!
0%
#55575000000
1!
1%
#55580000000
0!
0%
#55585000000
1!
1%
#55590000000
0!
0%
#55595000000
1!
1%
#55600000000
0!
0%
#55605000000
1!
1%
#55610000000
0!
0%
#55615000000
1!
1%
#55620000000
0!
0%
#55625000000
1!
1%
#55630000000
0!
0%
#55635000000
1!
1%
#55640000000
0!
0%
#55645000000
1!
1%
#55650000000
0!
0%
#55655000000
1!
1%
#55660000000
0!
0%
#55665000000
1!
1%
#55670000000
0!
0%
#55675000000
1!
1%
#55680000000
0!
0%
#55685000000
1!
1%
#55690000000
0!
0%
#55695000000
1!
1%
#55700000000
0!
0%
#55705000000
1!
1%
#55710000000
0!
0%
#55715000000
1!
1%
#55720000000
0!
0%
#55725000000
1!
1%
#55730000000
0!
0%
#55735000000
1!
1%
#55740000000
0!
0%
#55745000000
1!
1%
#55750000000
0!
0%
#55755000000
1!
1%
#55760000000
0!
0%
#55765000000
1!
1%
#55770000000
0!
0%
#55775000000
1!
1%
#55780000000
0!
0%
#55785000000
1!
1%
#55790000000
0!
0%
#55795000000
1!
1%
#55800000000
0!
0%
#55805000000
1!
1%
#55810000000
0!
0%
#55815000000
1!
1%
#55820000000
0!
0%
#55825000000
1!
1%
#55830000000
0!
0%
#55835000000
1!
1%
#55840000000
0!
0%
#55845000000
1!
1%
#55850000000
0!
0%
#55855000000
1!
1%
#55860000000
0!
0%
#55865000000
1!
1%
#55870000000
0!
0%
#55875000000
1!
1%
#55880000000
0!
0%
#55885000000
1!
1%
#55890000000
0!
0%
#55895000000
1!
1%
#55900000000
0!
0%
#55905000000
1!
1%
#55910000000
0!
0%
#55915000000
1!
1%
#55920000000
0!
0%
#55925000000
1!
1%
#55930000000
0!
0%
#55935000000
1!
1%
#55940000000
0!
0%
#55945000000
1!
1%
#55950000000
0!
0%
#55955000000
1!
1%
#55960000000
0!
0%
#55965000000
1!
1%
#55970000000
0!
0%
#55975000000
1!
1%
#55980000000
0!
0%
#55985000000
1!
1%
#55990000000
0!
0%
#55995000000
1!
1%
#56000000000
0!
0%
#56005000000
1!
1%
#56010000000
0!
0%
#56015000000
1!
1%
#56020000000
0!
0%
#56025000000
1!
1%
#56030000000
0!
0%
#56035000000
1!
1%
#56040000000
0!
0%
#56045000000
1!
1%
#56050000000
0!
0%
#56055000000
1!
1%
#56060000000
0!
0%
#56065000000
1!
1%
#56070000000
0!
0%
#56075000000
1!
1%
#56080000000
0!
0%
#56085000000
1!
1%
#56090000000
0!
0%
#56095000000
1!
1%
#56100000000
0!
0%
#56105000000
1!
1%
#56110000000
0!
0%
#56115000000
1!
1%
#56120000000
0!
0%
#56125000000
1!
1%
#56130000000
0!
0%
#56135000000
1!
1%
#56140000000
0!
0%
#56145000000
1!
1%
#56150000000
0!
0%
#56155000000
1!
1%
#56160000000
0!
0%
#56165000000
1!
1%
#56170000000
0!
0%
#56175000000
1!
1%
#56180000000
0!
0%
#56185000000
1!
1%
#56190000000
0!
0%
#56195000000
1!
1%
#56200000000
0!
0%
#56205000000
1!
1%
#56210000000
0!
0%
#56215000000
1!
1%
#56220000000
0!
0%
#56225000000
1!
1%
#56230000000
0!
0%
#56235000000
1!
1%
#56240000000
0!
0%
#56245000000
1!
1%
#56250000000
0!
0%
#56255000000
1!
1%
#56260000000
0!
0%
#56265000000
1!
1%
#56270000000
0!
0%
#56275000000
1!
1%
#56280000000
0!
0%
#56285000000
1!
1%
#56290000000
0!
0%
#56295000000
1!
1%
#56300000000
0!
0%
#56305000000
1!
1%
#56310000000
0!
0%
#56315000000
1!
1%
#56320000000
0!
0%
#56325000000
1!
1%
#56330000000
0!
0%
#56335000000
1!
1%
#56340000000
0!
0%
#56345000000
1!
1%
#56350000000
0!
0%
#56355000000
1!
1%
#56360000000
0!
0%
#56365000000
1!
1%
#56370000000
0!
0%
#56375000000
1!
1%
#56380000000
0!
0%
#56385000000
1!
1%
#56390000000
0!
0%
#56395000000
1!
1%
#56400000000
0!
0%
#56405000000
1!
1%
#56410000000
0!
0%
#56415000000
1!
1%
#56420000000
0!
0%
#56425000000
1!
1%
#56430000000
0!
0%
#56435000000
1!
1%
#56440000000
0!
0%
#56445000000
1!
1%
#56450000000
0!
0%
#56455000000
1!
1%
#56460000000
0!
0%
#56465000000
1!
1%
#56470000000
0!
0%
#56475000000
1!
1%
#56480000000
0!
0%
#56485000000
1!
1%
#56490000000
0!
0%
#56495000000
1!
1%
#56500000000
0!
0%
#56505000000
1!
1%
#56510000000
0!
0%
#56515000000
1!
1%
#56520000000
0!
0%
#56525000000
1!
1%
#56530000000
0!
0%
#56535000000
1!
1%
#56540000000
0!
0%
#56545000000
1!
1%
#56550000000
0!
0%
#56555000000
1!
1%
#56560000000
0!
0%
#56565000000
1!
1%
#56570000000
0!
0%
#56575000000
1!
1%
#56580000000
0!
0%
#56585000000
1!
1%
#56590000000
0!
0%
#56595000000
1!
1%
#56600000000
0!
0%
#56605000000
1!
1%
#56610000000
0!
0%
#56615000000
1!
1%
#56620000000
0!
0%
#56625000000
1!
1%
#56630000000
0!
0%
#56635000000
1!
1%
#56640000000
0!
0%
#56645000000
1!
1%
#56650000000
0!
0%
#56655000000
1!
1%
#56660000000
0!
0%
#56665000000
1!
1%
#56670000000
0!
0%
#56675000000
1!
1%
#56680000000
0!
0%
#56685000000
1!
1%
#56690000000
0!
0%
#56695000000
1!
1%
#56700000000
0!
0%
#56705000000
1!
1%
#56710000000
0!
0%
#56715000000
1!
1%
#56720000000
0!
0%
#56725000000
1!
1%
#56730000000
0!
0%
#56735000000
1!
1%
#56740000000
0!
0%
#56745000000
1!
1%
#56750000000
0!
0%
#56755000000
1!
1%
#56760000000
0!
0%
#56765000000
1!
1%
#56770000000
0!
0%
#56775000000
1!
1%
#56780000000
0!
0%
#56785000000
1!
1%
#56790000000
0!
0%
#56795000000
1!
1%
#56800000000
0!
0%
#56805000000
1!
1%
#56810000000
0!
0%
#56815000000
1!
1%
#56820000000
0!
0%
#56825000000
1!
1%
#56830000000
0!
0%
#56835000000
1!
1%
#56840000000
0!
0%
#56845000000
1!
1%
#56850000000
0!
0%
#56855000000
1!
1%
#56860000000
0!
0%
#56865000000
1!
1%
#56870000000
0!
0%
#56875000000
1!
1%
#56880000000
0!
0%
#56885000000
1!
1%
#56890000000
0!
0%
#56895000000
1!
1%
#56900000000
0!
0%
#56905000000
1!
1%
#56910000000
0!
0%
#56915000000
1!
1%
#56920000000
0!
0%
#56925000000
1!
1%
#56930000000
0!
0%
#56935000000
1!
1%
#56940000000
0!
0%
#56945000000
1!
1%
#56950000000
0!
0%
#56955000000
1!
1%
#56960000000
0!
0%
#56965000000
1!
1%
#56970000000
0!
0%
#56975000000
1!
1%
#56980000000
0!
0%
#56985000000
1!
1%
#56990000000
0!
0%
#56995000000
1!
1%
#57000000000
0!
0%
#57005000000
1!
1%
#57010000000
0!
0%
#57015000000
1!
1%
#57020000000
0!
0%
#57025000000
1!
1%
#57030000000
0!
0%
#57035000000
1!
1%
#57040000000
0!
0%
#57045000000
1!
1%
#57050000000
0!
0%
#57055000000
1!
1%
#57060000000
0!
0%
#57065000000
1!
1%
#57070000000
0!
0%
#57075000000
1!
1%
#57080000000
0!
0%
#57085000000
1!
1%
#57090000000
0!
0%
#57095000000
1!
1%
#57100000000
0!
0%
#57105000000
1!
1%
#57110000000
0!
0%
#57115000000
1!
1%
#57120000000
0!
0%
#57125000000
1!
1%
#57130000000
0!
0%
#57135000000
1!
1%
#57140000000
0!
0%
#57145000000
1!
1%
#57150000000
0!
0%
#57155000000
1!
1%
#57160000000
0!
0%
#57165000000
1!
1%
#57170000000
0!
0%
#57175000000
1!
1%
#57180000000
0!
0%
#57185000000
1!
1%
#57190000000
0!
0%
#57195000000
1!
1%
#57200000000
0!
0%
#57205000000
1!
1%
#57210000000
0!
0%
#57215000000
1!
1%
#57220000000
0!
0%
#57225000000
1!
1%
#57230000000
0!
0%
#57235000000
1!
1%
#57240000000
0!
0%
#57245000000
1!
1%
#57250000000
0!
0%
#57255000000
1!
1%
#57260000000
0!
0%
#57265000000
1!
1%
#57270000000
0!
0%
#57275000000
1!
1%
#57280000000
0!
0%
#57285000000
1!
1%
#57290000000
0!
0%
#57295000000
1!
1%
#57300000000
0!
0%
#57305000000
1!
1%
#57310000000
0!
0%
#57315000000
1!
1%
#57320000000
0!
0%
#57325000000
1!
1%
#57330000000
0!
0%
#57335000000
1!
1%
#57340000000
0!
0%
#57345000000
1!
1%
#57350000000
0!
0%
#57355000000
1!
1%
#57360000000
0!
0%
#57365000000
1!
1%
#57370000000
0!
0%
#57375000000
1!
1%
#57380000000
0!
0%
#57385000000
1!
1%
#57390000000
0!
0%
#57395000000
1!
1%
#57400000000
0!
0%
#57405000000
1!
1%
#57410000000
0!
0%
#57415000000
1!
1%
#57420000000
0!
0%
#57425000000
1!
1%
#57430000000
0!
0%
#57435000000
1!
1%
#57440000000
0!
0%
#57445000000
1!
1%
#57450000000
0!
0%
#57455000000
1!
1%
#57460000000
0!
0%
#57465000000
1!
1%
#57470000000
0!
0%
#57475000000
1!
1%
#57480000000
0!
0%
#57485000000
1!
1%
#57490000000
0!
0%
#57495000000
1!
1%
#57500000000
0!
0%
#57505000000
1!
1%
#57510000000
0!
0%
#57515000000
1!
1%
#57520000000
0!
0%
#57525000000
1!
1%
#57530000000
0!
0%
#57535000000
1!
1%
#57540000000
0!
0%
#57545000000
1!
1%
#57550000000
0!
0%
#57555000000
1!
1%
#57560000000
0!
0%
#57565000000
1!
1%
#57570000000
0!
0%
#57575000000
1!
1%
#57580000000
0!
0%
#57585000000
1!
1%
#57590000000
0!
0%
#57595000000
1!
1%
#57600000000
0!
0%
#57605000000
1!
1%
#57610000000
0!
0%
#57615000000
1!
1%
#57620000000
0!
0%
#57625000000
1!
1%
#57630000000
0!
0%
#57635000000
1!
1%
#57640000000
0!
0%
#57645000000
1!
1%
#57650000000
0!
0%
#57655000000
1!
1%
#57660000000
0!
0%
#57665000000
1!
1%
#57670000000
0!
0%
#57675000000
1!
1%
#57680000000
0!
0%
#57685000000
1!
1%
#57690000000
0!
0%
#57695000000
1!
1%
#57700000000
0!
0%
#57705000000
1!
1%
#57710000000
0!
0%
#57715000000
1!
1%
#57720000000
0!
0%
#57725000000
1!
1%
#57730000000
0!
0%
#57735000000
1!
1%
#57740000000
0!
0%
#57745000000
1!
1%
#57750000000
0!
0%
#57755000000
1!
1%
#57760000000
0!
0%
#57765000000
1!
1%
#57770000000
0!
0%
#57775000000
1!
1%
#57780000000
0!
0%
#57785000000
1!
1%
#57790000000
0!
0%
#57795000000
1!
1%
#57800000000
0!
0%
#57805000000
1!
1%
#57810000000
0!
0%
#57815000000
1!
1%
#57820000000
0!
0%
#57825000000
1!
1%
#57830000000
0!
0%
#57835000000
1!
1%
#57840000000
0!
0%
#57845000000
1!
1%
#57850000000
0!
0%
#57855000000
1!
1%
#57860000000
0!
0%
#57865000000
1!
1%
#57870000000
0!
0%
#57875000000
1!
1%
#57880000000
0!
0%
#57885000000
1!
1%
#57890000000
0!
0%
#57895000000
1!
1%
#57900000000
0!
0%
#57905000000
1!
1%
#57910000000
0!
0%
#57915000000
1!
1%
#57920000000
0!
0%
#57925000000
1!
1%
#57930000000
0!
0%
#57935000000
1!
1%
#57940000000
0!
0%
#57945000000
1!
1%
#57950000000
0!
0%
#57955000000
1!
1%
#57960000000
0!
0%
#57965000000
1!
1%
#57970000000
0!
0%
#57975000000
1!
1%
#57980000000
0!
0%
#57985000000
1!
1%
#57990000000
0!
0%
#57995000000
1!
1%
#58000000000
0!
0%
#58005000000
1!
1%
#58010000000
0!
0%
#58015000000
1!
1%
#58020000000
0!
0%
#58025000000
1!
1%
#58030000000
0!
0%
#58035000000
1!
1%
#58040000000
0!
0%
#58045000000
1!
1%
#58050000000
0!
0%
#58055000000
1!
1%
#58060000000
0!
0%
#58065000000
1!
1%
#58070000000
0!
0%
#58075000000
1!
1%
#58080000000
0!
0%
#58085000000
1!
1%
#58090000000
0!
0%
#58095000000
1!
1%
#58100000000
0!
0%
#58105000000
1!
1%
#58110000000
0!
0%
#58115000000
1!
1%
#58120000000
0!
0%
#58125000000
1!
1%
#58130000000
0!
0%
#58135000000
1!
1%
#58140000000
0!
0%
#58145000000
1!
1%
#58150000000
0!
0%
#58155000000
1!
1%
#58160000000
0!
0%
#58165000000
1!
1%
#58170000000
0!
0%
#58175000000
1!
1%
#58180000000
0!
0%
#58185000000
1!
1%
#58190000000
0!
0%
#58195000000
1!
1%
#58200000000
0!
0%
#58205000000
1!
1%
#58210000000
0!
0%
#58215000000
1!
1%
#58220000000
0!
0%
#58225000000
1!
1%
#58230000000
0!
0%
#58235000000
1!
1%
#58240000000
0!
0%
#58245000000
1!
1%
#58250000000
0!
0%
#58255000000
1!
1%
#58260000000
0!
0%
#58265000000
1!
1%
#58270000000
0!
0%
#58275000000
1!
1%
#58280000000
0!
0%
#58285000000
1!
1%
#58290000000
0!
0%
#58295000000
1!
1%
#58300000000
0!
0%
#58305000000
1!
1%
#58310000000
0!
0%
#58315000000
1!
1%
#58320000000
0!
0%
#58325000000
1!
1%
#58330000000
0!
0%
#58335000000
1!
1%
#58340000000
0!
0%
#58345000000
1!
1%
#58350000000
0!
0%
#58355000000
1!
1%
#58360000000
0!
0%
#58365000000
1!
1%
#58370000000
0!
0%
#58375000000
1!
1%
#58380000000
0!
0%
#58385000000
1!
1%
#58390000000
0!
0%
#58395000000
1!
1%
#58400000000
0!
0%
#58405000000
1!
1%
#58410000000
0!
0%
#58415000000
1!
1%
#58420000000
0!
0%
#58425000000
1!
1%
#58430000000
0!
0%
#58435000000
1!
1%
#58440000000
0!
0%
#58445000000
1!
1%
#58450000000
0!
0%
#58455000000
1!
1%
#58460000000
0!
0%
#58465000000
1!
1%
#58470000000
0!
0%
#58475000000
1!
1%
#58480000000
0!
0%
#58485000000
1!
1%
#58490000000
0!
0%
#58495000000
1!
1%
#58500000000
0!
0%
#58505000000
1!
1%
#58510000000
0!
0%
#58515000000
1!
1%
#58520000000
0!
0%
#58525000000
1!
1%
#58530000000
0!
0%
#58535000000
1!
1%
#58540000000
0!
0%
#58545000000
1!
1%
#58550000000
0!
0%
#58555000000
1!
1%
#58560000000
0!
0%
#58565000000
1!
1%
#58570000000
0!
0%
#58575000000
1!
1%
#58580000000
0!
0%
#58585000000
1!
1%
#58590000000
0!
0%
#58595000000
1!
1%
#58600000000
0!
0%
#58605000000
1!
1%
#58610000000
0!
0%
#58615000000
1!
1%
#58620000000
0!
0%
#58625000000
1!
1%
#58630000000
0!
0%
#58635000000
1!
1%
#58640000000
0!
0%
#58645000000
1!
1%
#58650000000
0!
0%
#58655000000
1!
1%
#58660000000
0!
0%
#58665000000
1!
1%
#58670000000
0!
0%
#58675000000
1!
1%
#58680000000
0!
0%
#58685000000
1!
1%
#58690000000
0!
0%
#58695000000
1!
1%
#58700000000
0!
0%
#58705000000
1!
1%
#58710000000
0!
0%
#58715000000
1!
1%
#58720000000
0!
0%
#58725000000
1!
1%
#58730000000
0!
0%
#58735000000
1!
1%
#58740000000
0!
0%
#58745000000
1!
1%
#58750000000
0!
0%
#58755000000
1!
1%
#58760000000
0!
0%
#58765000000
1!
1%
#58770000000
0!
0%
#58775000000
1!
1%
#58780000000
0!
0%
#58785000000
1!
1%
#58790000000
0!
0%
#58795000000
1!
1%
#58800000000
0!
0%
#58805000000
1!
1%
#58810000000
0!
0%
#58815000000
1!
1%
#58820000000
0!
0%
#58825000000
1!
1%
#58830000000
0!
0%
#58835000000
1!
1%
#58840000000
0!
0%
#58845000000
1!
1%
#58850000000
0!
0%
#58855000000
1!
1%
#58860000000
0!
0%
#58865000000
1!
1%
#58870000000
0!
0%
#58875000000
1!
1%
#58880000000
0!
0%
#58885000000
1!
1%
#58890000000
0!
0%
#58895000000
1!
1%
#58900000000
0!
0%
#58905000000
1!
1%
#58910000000
0!
0%
#58915000000
1!
1%
#58920000000
0!
0%
#58925000000
1!
1%
#58930000000
0!
0%
#58935000000
1!
1%
#58940000000
0!
0%
#58945000000
1!
1%
#58950000000
0!
0%
#58955000000
1!
1%
#58960000000
0!
0%
#58965000000
1!
1%
#58970000000
0!
0%
#58975000000
1!
1%
#58980000000
0!
0%
#58985000000
1!
1%
#58990000000
0!
0%
#58995000000
1!
1%
#59000000000
0!
0%
#59005000000
1!
1%
#59010000000
0!
0%
#59015000000
1!
1%
#59020000000
0!
0%
#59025000000
1!
1%
#59030000000
0!
0%
#59035000000
1!
1%
#59040000000
0!
0%
#59045000000
1!
1%
#59050000000
0!
0%
#59055000000
1!
1%
#59060000000
0!
0%
#59065000000
1!
1%
#59070000000
0!
0%
#59075000000
1!
1%
#59080000000
0!
0%
#59085000000
1!
1%
#59090000000
0!
0%
#59095000000
1!
1%
#59100000000
0!
0%
#59105000000
1!
1%
#59110000000
0!
0%
#59115000000
1!
1%
#59120000000
0!
0%
#59125000000
1!
1%
#59130000000
0!
0%
#59135000000
1!
1%
#59140000000
0!
0%
#59145000000
1!
1%
#59150000000
0!
0%
#59155000000
1!
1%
#59160000000
0!
0%
#59165000000
1!
1%
#59170000000
0!
0%
#59175000000
1!
1%
#59180000000
0!
0%
#59185000000
1!
1%
#59190000000
0!
0%
#59195000000
1!
1%
#59200000000
0!
0%
#59205000000
1!
1%
#59210000000
0!
0%
#59215000000
1!
1%
#59220000000
0!
0%
#59225000000
1!
1%
#59230000000
0!
0%
#59235000000
1!
1%
#59240000000
0!
0%
#59245000000
1!
1%
#59250000000
0!
0%
#59255000000
1!
1%
#59260000000
0!
0%
#59265000000
1!
1%
#59270000000
0!
0%
#59275000000
1!
1%
#59280000000
0!
0%
#59285000000
1!
1%
#59290000000
0!
0%
#59295000000
1!
1%
#59300000000
0!
0%
#59305000000
1!
1%
#59310000000
0!
0%
#59315000000
1!
1%
#59320000000
0!
0%
#59325000000
1!
1%
#59330000000
0!
0%
#59335000000
1!
1%
#59340000000
0!
0%
#59345000000
1!
1%
#59350000000
0!
0%
#59355000000
1!
1%
#59360000000
0!
0%
#59365000000
1!
1%
#59370000000
0!
0%
#59375000000
1!
1%
#59380000000
0!
0%
#59385000000
1!
1%
#59390000000
0!
0%
#59395000000
1!
1%
#59400000000
0!
0%
#59405000000
1!
1%
#59410000000
0!
0%
#59415000000
1!
1%
#59420000000
0!
0%
#59425000000
1!
1%
#59430000000
0!
0%
#59435000000
1!
1%
#59440000000
0!
0%
#59445000000
1!
1%
#59450000000
0!
0%
#59455000000
1!
1%
#59460000000
0!
0%
#59465000000
1!
1%
#59470000000
0!
0%
#59475000000
1!
1%
#59480000000
0!
0%
#59485000000
1!
1%
#59490000000
0!
0%
#59495000000
1!
1%
#59500000000
0!
0%
#59505000000
1!
1%
#59510000000
0!
0%
#59515000000
1!
1%
#59520000000
0!
0%
#59525000000
1!
1%
#59530000000
0!
0%
#59535000000
1!
1%
#59540000000
0!
0%
#59545000000
1!
1%
#59550000000
0!
0%
#59555000000
1!
1%
#59560000000
0!
0%
#59565000000
1!
1%
#59570000000
0!
0%
#59575000000
1!
1%
#59580000000
0!
0%
#59585000000
1!
1%
#59590000000
0!
0%
#59595000000
1!
1%
#59600000000
0!
0%
#59605000000
1!
1%
#59610000000
0!
0%
#59615000000
1!
1%
#59620000000
0!
0%
#59625000000
1!
1%
#59630000000
0!
0%
#59635000000
1!
1%
#59640000000
0!
0%
#59645000000
1!
1%
#59650000000
0!
0%
#59655000000
1!
1%
#59660000000
0!
0%
#59665000000
1!
1%
#59670000000
0!
0%
#59675000000
1!
1%
#59680000000
0!
0%
#59685000000
1!
1%
#59690000000
0!
0%
#59695000000
1!
1%
#59700000000
0!
0%
#59705000000
1!
1%
#59710000000
0!
0%
#59715000000
1!
1%
#59720000000
0!
0%
#59725000000
1!
1%
#59730000000
0!
0%
#59735000000
1!
1%
#59740000000
0!
0%
#59745000000
1!
1%
#59750000000
0!
0%
#59755000000
1!
1%
#59760000000
0!
0%
#59765000000
1!
1%
#59770000000
0!
0%
#59775000000
1!
1%
#59780000000
0!
0%
#59785000000
1!
1%
#59790000000
0!
0%
#59795000000
1!
1%
#59800000000
0!
0%
#59805000000
1!
1%
#59810000000
0!
0%
#59815000000
1!
1%
#59820000000
0!
0%
#59825000000
1!
1%
#59830000000
0!
0%
#59835000000
1!
1%
#59840000000
0!
0%
#59845000000
1!
1%
#59850000000
0!
0%
#59855000000
1!
1%
#59860000000
0!
0%
#59865000000
1!
1%
#59870000000
0!
0%
#59875000000
1!
1%
#59880000000
0!
0%
#59885000000
1!
1%
#59890000000
0!
0%
#59895000000
1!
1%
#59900000000
0!
0%
#59905000000
1!
1%
#59910000000
0!
0%
#59915000000
1!
1%
#59920000000
0!
0%
#59925000000
1!
1%
#59930000000
0!
0%
#59935000000
1!
1%
#59940000000
0!
0%
#59945000000
1!
1%
#59950000000
0!
0%
#59955000000
1!
1%
#59960000000
0!
0%
#59965000000
1!
1%
#59970000000
0!
0%
#59975000000
1!
1%
#59980000000
0!
0%
#59985000000
1!
1%
#59990000000
0!
0%
#59995000000
1!
1%
#60000000000
0!
0%
#60005000000
1!
1%
#60010000000
0!
0%
#60015000000
1!
1%
#60020000000
0!
0%
#60025000000
1!
1%
#60030000000
0!
0%
#60035000000
1!
1%
#60040000000
0!
0%
#60045000000
1!
1%
#60050000000
0!
0%
#60055000000
1!
1%
#60060000000
0!
0%
#60065000000
1!
1%
#60070000000
0!
0%
#60075000000
1!
1%
#60080000000
0!
0%
#60085000000
1!
1%
#60090000000
0!
0%
#60095000000
1!
1%
#60100000000
0!
0%
#60105000000
1!
1%
#60110000000
0!
0%
#60115000000
1!
1%
#60120000000
0!
0%
#60125000000
1!
1%
#60130000000
0!
0%
#60135000000
1!
1%
#60140000000
0!
0%
#60145000000
1!
1%
#60150000000
0!
0%
#60155000000
1!
1%
#60160000000
0!
0%
#60165000000
1!
1%
#60170000000
0!
0%
#60175000000
1!
1%
#60180000000
0!
0%
#60185000000
1!
1%
#60190000000
0!
0%
#60195000000
1!
1%
#60200000000
0!
0%
#60205000000
1!
1%
#60210000000
0!
0%
#60215000000
1!
1%
#60220000000
0!
0%
#60225000000
1!
1%
#60230000000
0!
0%
#60235000000
1!
1%
#60240000000
0!
0%
#60245000000
1!
1%
#60250000000
0!
0%
#60255000000
1!
1%
#60260000000
0!
0%
#60265000000
1!
1%
#60270000000
0!
0%
#60275000000
1!
1%
#60280000000
0!
0%
#60285000000
1!
1%
#60290000000
0!
0%
#60295000000
1!
1%
#60300000000
0!
0%
#60305000000
1!
1%
#60310000000
0!
0%
#60315000000
1!
1%
#60320000000
0!
0%
#60325000000
1!
1%
#60330000000
0!
0%
#60335000000
1!
1%
#60340000000
0!
0%
#60345000000
1!
1%
#60350000000
0!
0%
#60355000000
1!
1%
#60360000000
0!
0%
#60365000000
1!
1%
#60370000000
0!
0%
#60375000000
1!
1%
#60380000000
0!
0%
#60385000000
1!
1%
#60390000000
0!
0%
#60395000000
1!
1%
#60400000000
0!
0%
#60405000000
1!
1%
#60410000000
0!
0%
#60415000000
1!
1%
#60420000000
0!
0%
#60425000000
1!
1%
#60430000000
0!
0%
#60435000000
1!
1%
#60440000000
0!
0%
#60445000000
1!
1%
#60450000000
0!
0%
#60455000000
1!
1%
#60460000000
0!
0%
#60465000000
1!
1%
#60470000000
0!
0%
#60475000000
1!
1%
#60480000000
0!
0%
#60485000000
1!
1%
#60490000000
0!
0%
#60495000000
1!
1%
#60500000000
0!
0%
#60505000000
1!
1%
#60510000000
0!
0%
#60515000000
1!
1%
#60520000000
0!
0%
#60525000000
1!
1%
#60530000000
0!
0%
#60535000000
1!
1%
#60540000000
0!
0%
#60545000000
1!
1%
#60550000000
0!
0%
#60555000000
1!
1%
#60560000000
0!
0%
#60565000000
1!
1%
#60570000000
0!
0%
#60575000000
1!
1%
#60580000000
0!
0%
#60585000000
1!
1%
#60590000000
0!
0%
#60595000000
1!
1%
#60600000000
0!
0%
#60605000000
1!
1%
#60610000000
0!
0%
#60615000000
1!
1%
#60620000000
0!
0%
#60625000000
1!
1%
#60630000000
0!
0%
#60635000000
1!
1%
#60640000000
0!
0%
#60645000000
1!
1%
#60650000000
0!
0%
#60655000000
1!
1%
#60660000000
0!
0%
#60665000000
1!
1%
#60670000000
0!
0%
#60675000000
1!
1%
#60680000000
0!
0%
#60685000000
1!
1%
#60690000000
0!
0%
#60695000000
1!
1%
#60700000000
0!
0%
#60705000000
1!
1%
#60710000000
0!
0%
#60715000000
1!
1%
#60720000000
0!
0%
#60725000000
1!
1%
#60730000000
0!
0%
#60735000000
1!
1%
#60740000000
0!
0%
#60745000000
1!
1%
#60750000000
0!
0%
#60755000000
1!
1%
#60760000000
0!
0%
#60765000000
1!
1%
#60770000000
0!
0%
#60775000000
1!
1%
#60780000000
0!
0%
#60785000000
1!
1%
#60790000000
0!
0%
#60795000000
1!
1%
#60800000000
0!
0%
#60805000000
1!
1%
#60810000000
0!
0%
#60815000000
1!
1%
#60820000000
0!
0%
#60825000000
1!
1%
#60830000000
0!
0%
#60835000000
1!
1%
#60840000000
0!
0%
#60845000000
1!
1%
#60850000000
0!
0%
#60855000000
1!
1%
#60860000000
0!
0%
#60865000000
1!
1%
#60870000000
0!
0%
#60875000000
1!
1%
#60880000000
0!
0%
#60885000000
1!
1%
#60890000000
0!
0%
#60895000000
1!
1%
#60900000000
0!
0%
#60905000000
1!
1%
#60910000000
0!
0%
#60915000000
1!
1%
#60920000000
0!
0%
#60925000000
1!
1%
#60930000000
0!
0%
#60935000000
1!
1%
#60940000000
0!
0%
#60945000000
1!
1%
#60950000000
0!
0%
#60955000000
1!
1%
#60960000000
0!
0%
#60965000000
1!
1%
#60970000000
0!
0%
#60975000000
1!
1%
#60980000000
0!
0%
#60985000000
1!
1%
#60990000000
0!
0%
#60995000000
1!
1%
#61000000000
0!
0%
#61005000000
1!
1%
#61010000000
0!
0%
#61015000000
1!
1%
#61020000000
0!
0%
#61025000000
1!
1%
#61030000000
0!
0%
#61035000000
1!
1%
#61040000000
0!
0%
#61045000000
1!
1%
#61050000000
0!
0%
#61055000000
1!
1%
#61060000000
0!
0%
#61065000000
1!
1%
#61070000000
0!
0%
#61075000000
1!
1%
#61080000000
0!
0%
#61085000000
1!
1%
#61090000000
0!
0%
#61095000000
1!
1%
#61100000000
0!
0%
#61105000000
1!
1%
#61110000000
0!
0%
#61115000000
1!
1%
#61120000000
0!
0%
#61125000000
1!
1%
#61130000000
0!
0%
#61135000000
1!
1%
#61140000000
0!
0%
#61145000000
1!
1%
#61150000000
0!
0%
#61155000000
1!
1%
#61160000000
0!
0%
#61165000000
1!
1%
#61170000000
0!
0%
#61175000000
1!
1%
#61180000000
0!
0%
#61185000000
1!
1%
#61190000000
0!
0%
#61195000000
1!
1%
#61200000000
0!
0%
#61205000000
1!
1%
#61210000000
0!
0%
#61215000000
1!
1%
#61220000000
0!
0%
#61225000000
1!
1%
#61230000000
0!
0%
#61235000000
1!
1%
#61240000000
0!
0%
#61245000000
1!
1%
#61250000000
0!
0%
#61255000000
1!
1%
#61260000000
0!
0%
#61265000000
1!
1%
#61270000000
0!
0%
#61275000000
1!
1%
#61280000000
0!
0%
#61285000000
1!
1%
#61290000000
0!
0%
#61295000000
1!
1%
#61300000000
0!
0%
#61305000000
1!
1%
#61310000000
0!
0%
#61315000000
1!
1%
#61320000000
0!
0%
#61325000000
1!
1%
#61330000000
0!
0%
#61335000000
1!
1%
#61340000000
0!
0%
#61345000000
1!
1%
#61350000000
0!
0%
#61355000000
1!
1%
#61360000000
0!
0%
#61365000000
1!
1%
#61370000000
0!
0%
#61375000000
1!
1%
#61380000000
0!
0%
#61385000000
1!
1%
#61390000000
0!
0%
#61395000000
1!
1%
#61400000000
0!
0%
#61405000000
1!
1%
#61410000000
0!
0%
#61415000000
1!
1%
#61420000000
0!
0%
#61425000000
1!
1%
#61430000000
0!
0%
#61435000000
1!
1%
#61440000000
0!
0%
#61445000000
1!
1%
#61450000000
0!
0%
#61455000000
1!
1%
#61460000000
0!
0%
#61465000000
1!
1%
#61470000000
0!
0%
#61475000000
1!
1%
#61480000000
0!
0%
#61485000000
1!
1%
#61490000000
0!
0%
#61495000000
1!
1%
#61500000000
0!
0%
#61505000000
1!
1%
#61510000000
0!
0%
#61515000000
1!
1%
#61520000000
0!
0%
#61525000000
1!
1%
#61530000000
0!
0%
#61535000000
1!
1%
#61540000000
0!
0%
#61545000000
1!
1%
#61550000000
0!
0%
#61555000000
1!
1%
#61560000000
0!
0%
#61565000000
1!
1%
#61570000000
0!
0%
#61575000000
1!
1%
#61580000000
0!
0%
#61585000000
1!
1%
#61590000000
0!
0%
#61595000000
1!
1%
#61600000000
0!
0%
#61605000000
1!
1%
#61610000000
0!
0%
#61615000000
1!
1%
#61620000000
0!
0%
#61625000000
1!
1%
#61630000000
0!
0%
#61635000000
1!
1%
#61640000000
0!
0%
#61645000000
1!
1%
#61650000000
0!
0%
#61655000000
1!
1%
#61660000000
0!
0%
#61665000000
1!
1%
#61670000000
0!
0%
#61675000000
1!
1%
#61680000000
0!
0%
#61685000000
1!
1%
#61690000000
0!
0%
#61695000000
1!
1%
#61700000000
0!
0%
#61705000000
1!
1%
#61710000000
0!
0%
#61715000000
1!
1%
#61720000000
0!
0%
#61725000000
1!
1%
#61730000000
0!
0%
#61735000000
1!
1%
#61740000000
0!
0%
#61745000000
1!
1%
#61750000000
0!
0%
#61755000000
1!
1%
#61760000000
0!
0%
#61765000000
1!
1%
#61770000000
0!
0%
#61775000000
1!
1%
#61780000000
0!
0%
#61785000000
1!
1%
#61790000000
0!
0%
#61795000000
1!
1%
#61800000000
0!
0%
#61805000000
1!
1%
#61810000000
0!
0%
#61815000000
1!
1%
#61820000000
0!
0%
#61825000000
1!
1%
#61830000000
0!
0%
#61835000000
1!
1%
#61840000000
0!
0%
#61845000000
1!
1%
#61850000000
0!
0%
#61855000000
1!
1%
#61860000000
0!
0%
#61865000000
1!
1%
#61870000000
0!
0%
#61875000000
1!
1%
#61880000000
0!
0%
#61885000000
1!
1%
#61890000000
0!
0%
#61895000000
1!
1%
#61900000000
0!
0%
#61905000000
1!
1%
#61910000000
0!
0%
#61915000000
1!
1%
#61920000000
0!
0%
#61925000000
1!
1%
#61930000000
0!
0%
#61935000000
1!
1%
#61940000000
0!
0%
#61945000000
1!
1%
#61950000000
0!
0%
#61955000000
1!
1%
#61960000000
0!
0%
#61965000000
1!
1%
#61970000000
0!
0%
#61975000000
1!
1%
#61980000000
0!
0%
#61985000000
1!
1%
#61990000000
0!
0%
#61995000000
1!
1%
#62000000000
0!
0%
#62005000000
1!
1%
#62010000000
0!
0%
#62015000000
1!
1%
#62020000000
0!
0%
#62025000000
1!
1%
#62030000000
0!
0%
#62035000000
1!
1%
#62040000000
0!
0%
#62045000000
1!
1%
#62050000000
0!
0%
#62055000000
1!
1%
#62060000000
0!
0%
#62065000000
1!
1%
#62070000000
0!
0%
#62075000000
1!
1%
#62080000000
0!
0%
#62085000000
1!
1%
#62090000000
0!
0%
#62095000000
1!
1%
#62100000000
0!
0%
#62105000000
1!
1%
#62110000000
0!
0%
#62115000000
1!
1%
#62120000000
0!
0%
#62125000000
1!
1%
#62130000000
0!
0%
#62135000000
1!
1%
#62140000000
0!
0%
#62145000000
1!
1%
#62150000000
0!
0%
#62155000000
1!
1%
#62160000000
0!
0%
#62165000000
1!
1%
#62170000000
0!
0%
#62175000000
1!
1%
#62180000000
0!
0%
#62185000000
1!
1%
#62190000000
0!
0%
#62195000000
1!
1%
#62200000000
0!
0%
#62205000000
1!
1%
#62210000000
0!
0%
#62215000000
1!
1%
#62220000000
0!
0%
#62225000000
1!
1%
#62230000000
0!
0%
#62235000000
1!
1%
#62240000000
0!
0%
#62245000000
1!
1%
#62250000000
0!
0%
#62255000000
1!
1%
#62260000000
0!
0%
#62265000000
1!
1%
#62270000000
0!
0%
#62275000000
1!
1%
#62280000000
0!
0%
#62285000000
1!
1%
#62290000000
0!
0%
#62295000000
1!
1%
#62300000000
0!
0%
#62305000000
1!
1%
#62310000000
0!
0%
#62315000000
1!
1%
#62320000000
0!
0%
#62325000000
1!
1%
#62330000000
0!
0%
#62335000000
1!
1%
#62340000000
0!
0%
#62345000000
1!
1%
#62350000000
0!
0%
#62355000000
1!
1%
#62360000000
0!
0%
#62365000000
1!
1%
#62370000000
0!
0%
#62375000000
1!
1%
#62380000000
0!
0%
#62385000000
1!
1%
#62390000000
0!
0%
#62395000000
1!
1%
#62400000000
0!
0%
#62405000000
1!
1%
#62410000000
0!
0%
#62415000000
1!
1%
#62420000000
0!
0%
#62425000000
1!
1%
#62430000000
0!
0%
#62435000000
1!
1%
#62440000000
0!
0%
#62445000000
1!
1%
#62450000000
0!
0%
#62455000000
1!
1%
#62460000000
0!
0%
#62465000000
1!
1%
#62470000000
0!
0%
#62475000000
1!
1%
#62480000000
0!
0%
#62485000000
1!
1%
#62490000000
0!
0%
#62495000000
1!
1%
#62500000000
0!
0%
#62505000000
1!
1%
#62510000000
0!
0%
#62515000000
1!
1%
#62520000000
0!
0%
#62525000000
1!
1%
#62530000000
0!
0%
#62535000000
1!
1%
#62540000000
0!
0%
#62545000000
1!
1%
#62550000000
0!
0%
#62555000000
1!
1%
#62560000000
0!
0%
#62565000000
1!
1%
#62570000000
0!
0%
#62575000000
1!
1%
#62580000000
0!
0%
#62585000000
1!
1%
#62590000000
0!
0%
#62595000000
1!
1%
#62600000000
0!
0%
#62605000000
1!
1%
#62610000000
0!
0%
#62615000000
1!
1%
#62620000000
0!
0%
#62625000000
1!
1%
#62630000000
0!
0%
#62635000000
1!
1%
#62640000000
0!
0%
#62645000000
1!
1%
#62650000000
0!
0%
#62655000000
1!
1%
#62660000000
0!
0%
#62665000000
1!
1%
#62670000000
0!
0%
#62675000000
1!
1%
#62680000000
0!
0%
#62685000000
1!
1%
#62690000000
0!
0%
#62695000000
1!
1%
#62700000000
0!
0%
#62705000000
1!
1%
#62710000000
0!
0%
#62715000000
1!
1%
#62720000000
0!
0%
#62725000000
1!
1%
#62730000000
0!
0%
#62735000000
1!
1%
#62740000000
0!
0%
#62745000000
1!
1%
#62750000000
0!
0%
#62755000000
1!
1%
#62760000000
0!
0%
#62765000000
1!
1%
#62770000000
0!
0%
#62775000000
1!
1%
#62780000000
0!
0%
#62785000000
1!
1%
#62790000000
0!
0%
#62795000000
1!
1%
#62800000000
0!
0%
#62805000000
1!
1%
#62810000000
0!
0%
#62815000000
1!
1%
#62820000000
0!
0%
#62825000000
1!
1%
#62830000000
0!
0%
#62835000000
1!
1%
#62840000000
0!
0%
#62845000000
1!
1%
#62850000000
0!
0%
#62855000000
1!
1%
#62860000000
0!
0%
#62865000000
1!
1%
#62870000000
0!
0%
#62875000000
1!
1%
#62880000000
0!
0%
#62885000000
1!
1%
#62890000000
0!
0%
#62895000000
1!
1%
#62900000000
0!
0%
#62905000000
1!
1%
#62910000000
0!
0%
#62915000000
1!
1%
#62920000000
0!
0%
#62925000000
1!
1%
#62930000000
0!
0%
#62935000000
1!
1%
#62940000000
0!
0%
#62945000000
1!
1%
#62950000000
0!
0%
#62955000000
1!
1%
#62960000000
0!
0%
#62965000000
1!
1%
#62970000000
0!
0%
#62975000000
1!
1%
#62980000000
0!
0%
#62985000000
1!
1%
#62990000000
0!
0%
#62995000000
1!
1%
#63000000000
0!
0%
#63005000000
1!
1%
#63010000000
0!
0%
#63015000000
1!
1%
#63020000000
0!
0%
#63025000000
1!
1%
#63030000000
0!
0%
#63035000000
1!
1%
#63040000000
0!
0%
#63045000000
1!
1%
#63050000000
0!
0%
#63055000000
1!
1%
#63060000000
0!
0%
#63065000000
1!
1%
#63070000000
0!
0%
#63075000000
1!
1%
#63080000000
0!
0%
#63085000000
1!
1%
#63090000000
0!
0%
#63095000000
1!
1%
#63100000000
0!
0%
#63105000000
1!
1%
#63110000000
0!
0%
#63115000000
1!
1%
#63120000000
0!
0%
#63125000000
1!
1%
#63130000000
0!
0%
#63135000000
1!
1%
#63140000000
0!
0%
#63145000000
1!
1%
#63150000000
0!
0%
#63155000000
1!
1%
#63160000000
0!
0%
#63165000000
1!
1%
#63170000000
0!
0%
#63175000000
1!
1%
#63180000000
0!
0%
#63185000000
1!
1%
#63190000000
0!
0%
#63195000000
1!
1%
#63200000000
0!
0%
#63205000000
1!
1%
#63210000000
0!
0%
#63215000000
1!
1%
#63220000000
0!
0%
#63225000000
1!
1%
#63230000000
0!
0%
#63235000000
1!
1%
#63240000000
0!
0%
#63245000000
1!
1%
#63250000000
0!
0%
#63255000000
1!
1%
#63260000000
0!
0%
#63265000000
1!
1%
#63270000000
0!
0%
#63275000000
1!
1%
#63280000000
0!
0%
#63285000000
1!
1%
#63290000000
0!
0%
#63295000000
1!
1%
#63300000000
0!
0%
#63305000000
1!
1%
#63310000000
0!
0%
#63315000000
1!
1%
#63320000000
0!
0%
#63325000000
1!
1%
#63330000000
0!
0%
#63335000000
1!
1%
#63340000000
0!
0%
#63345000000
1!
1%
#63350000000
0!
0%
#63355000000
1!
1%
#63360000000
0!
0%
#63365000000
1!
1%
#63370000000
0!
0%
#63375000000
1!
1%
#63380000000
0!
0%
#63385000000
1!
1%
#63390000000
0!
0%
#63395000000
1!
1%
#63400000000
0!
0%
#63405000000
1!
1%
#63410000000
0!
0%
#63415000000
1!
1%
#63420000000
0!
0%
#63425000000
1!
1%
#63430000000
0!
0%
#63435000000
1!
1%
#63440000000
0!
0%
#63445000000
1!
1%
#63450000000
0!
0%
#63455000000
1!
1%
#63460000000
0!
0%
#63465000000
1!
1%
#63470000000
0!
0%
#63475000000
1!
1%
#63480000000
0!
0%
#63485000000
1!
1%
#63490000000
0!
0%
#63495000000
1!
1%
#63500000000
0!
0%
#63505000000
1!
1%
#63510000000
0!
0%
#63515000000
1!
1%
#63520000000
0!
0%
#63525000000
1!
1%
#63530000000
0!
0%
#63535000000
1!
1%
#63540000000
0!
0%
#63545000000
1!
1%
#63550000000
0!
0%
#63555000000
1!
1%
#63560000000
0!
0%
#63565000000
1!
1%
#63570000000
0!
0%
#63575000000
1!
1%
#63580000000
0!
0%
#63585000000
1!
1%
#63590000000
0!
0%
#63595000000
1!
1%
#63600000000
0!
0%
#63605000000
1!
1%
#63610000000
0!
0%
#63615000000
1!
1%
#63620000000
0!
0%
#63625000000
1!
1%
#63630000000
0!
0%
#63635000000
1!
1%
#63640000000
0!
0%
#63645000000
1!
1%
#63650000000
0!
0%
#63655000000
1!
1%
#63660000000
0!
0%
#63665000000
1!
1%
#63670000000
0!
0%
#63675000000
1!
1%
#63680000000
0!
0%
#63685000000
1!
1%
#63690000000
0!
0%
#63695000000
1!
1%
#63700000000
0!
0%
#63705000000
1!
1%
#63710000000
0!
0%
#63715000000
1!
1%
#63720000000
0!
0%
#63725000000
1!
1%
#63730000000
0!
0%
#63735000000
1!
1%
#63740000000
0!
0%
#63745000000
1!
1%
#63750000000
0!
0%
#63755000000
1!
1%
#63760000000
0!
0%
#63765000000
1!
1%
#63770000000
0!
0%
#63775000000
1!
1%
#63780000000
0!
0%
#63785000000
1!
1%
#63790000000
0!
0%
#63795000000
1!
1%
#63800000000
0!
0%
#63805000000
1!
1%
#63810000000
0!
0%
#63815000000
1!
1%
#63820000000
0!
0%
#63825000000
1!
1%
#63830000000
0!
0%
#63835000000
1!
1%
#63840000000
0!
0%
#63845000000
1!
1%
#63850000000
0!
0%
#63855000000
1!
1%
#63860000000
0!
0%
#63865000000
1!
1%
#63870000000
0!
0%
#63875000000
1!
1%
#63880000000
0!
0%
#63885000000
1!
1%
#63890000000
0!
0%
#63895000000
1!
1%
#63900000000
0!
0%
#63905000000
1!
1%
#63910000000
0!
0%
#63915000000
1!
1%
#63920000000
0!
0%
#63925000000
1!
1%
#63930000000
0!
0%
#63935000000
1!
1%
#63940000000
0!
0%
#63945000000
1!
1%
#63950000000
0!
0%
#63955000000
1!
1%
#63960000000
0!
0%
#63965000000
1!
1%
#63970000000
0!
0%
#63975000000
1!
1%
#63980000000
0!
0%
#63985000000
1!
1%
#63990000000
0!
0%
#63995000000
1!
1%
#64000000000
0!
0%
#64005000000
1!
1%
#64010000000
0!
0%
#64015000000
1!
1%
#64020000000
0!
0%
#64025000000
1!
1%
#64030000000
0!
0%
#64035000000
1!
1%
#64040000000
0!
0%
#64045000000
1!
1%
#64050000000
0!
0%
#64055000000
1!
1%
#64060000000
0!
0%
#64065000000
1!
1%
#64070000000
0!
0%
#64075000000
1!
1%
#64080000000
0!
0%
#64085000000
1!
1%
#64090000000
0!
0%
#64095000000
1!
1%
#64100000000
0!
0%
#64105000000
1!
1%
#64110000000
0!
0%
#64115000000
1!
1%
#64120000000
0!
0%
#64125000000
1!
1%
#64130000000
0!
0%
#64135000000
1!
1%
#64140000000
0!
0%
#64145000000
1!
1%
#64150000000
0!
0%
#64155000000
1!
1%
#64160000000
0!
0%
#64165000000
1!
1%
#64170000000
0!
0%
#64175000000
1!
1%
#64180000000
0!
0%
#64185000000
1!
1%
#64190000000
0!
0%
#64195000000
1!
1%
#64200000000
0!
0%
#64205000000
1!
1%
#64210000000
0!
0%
#64215000000
1!
1%
#64220000000
0!
0%
#64225000000
1!
1%
#64230000000
0!
0%
#64235000000
1!
1%
#64240000000
0!
0%
#64245000000
1!
1%
#64250000000
0!
0%
#64255000000
1!
1%
#64260000000
0!
0%
#64265000000
1!
1%
#64270000000
0!
0%
#64275000000
1!
1%
#64280000000
0!
0%
#64285000000
1!
1%
#64290000000
0!
0%
#64295000000
1!
1%
#64300000000
0!
0%
#64305000000
1!
1%
#64310000000
0!
0%
#64315000000
1!
1%
#64320000000
0!
0%
#64325000000
1!
1%
#64330000000
0!
0%
#64335000000
1!
1%
#64340000000
0!
0%
#64345000000
1!
1%
#64350000000
0!
0%
#64355000000
1!
1%
#64360000000
0!
0%
#64365000000
1!
1%
#64370000000
0!
0%
#64375000000
1!
1%
#64380000000
0!
0%
#64385000000
1!
1%
#64390000000
0!
0%
#64395000000
1!
1%
#64400000000
0!
0%
#64405000000
1!
1%
#64410000000
0!
0%
#64415000000
1!
1%
#64420000000
0!
0%
#64425000000
1!
1%
#64430000000
0!
0%
#64435000000
1!
1%
#64440000000
0!
0%
#64445000000
1!
1%
#64450000000
0!
0%
#64455000000
1!
1%
#64460000000
0!
0%
#64465000000
1!
1%
#64470000000
0!
0%
#64475000000
1!
1%
#64480000000
0!
0%
#64485000000
1!
1%
#64490000000
0!
0%
#64495000000
1!
1%
#64500000000
0!
0%
#64505000000
1!
1%
#64510000000
0!
0%
#64515000000
1!
1%
#64520000000
0!
0%
#64525000000
1!
1%
#64530000000
0!
0%
#64535000000
1!
1%
#64540000000
0!
0%
#64545000000
1!
1%
#64550000000
0!
0%
#64555000000
1!
1%
#64560000000
0!
0%
#64565000000
1!
1%
#64570000000
0!
0%
#64575000000
1!
1%
#64580000000
0!
0%
#64585000000
1!
1%
#64590000000
0!
0%
#64595000000
1!
1%
#64600000000
0!
0%
#64605000000
1!
1%
#64610000000
0!
0%
#64615000000
1!
1%
#64620000000
0!
0%
#64625000000
1!
1%
#64630000000
0!
0%
#64635000000
1!
1%
#64640000000
0!
0%
#64645000000
1!
1%
#64650000000
0!
0%
#64655000000
1!
1%
#64660000000
0!
0%
#64665000000
1!
1%
#64670000000
0!
0%
#64675000000
1!
1%
#64680000000
0!
0%
#64685000000
1!
1%
#64690000000
0!
0%
#64695000000
1!
1%
#64700000000
0!
0%
#64705000000
1!
1%
#64710000000
0!
0%
#64715000000
1!
1%
#64720000000
0!
0%
#64725000000
1!
1%
#64730000000
0!
0%
#64735000000
1!
1%
#64740000000
0!
0%
#64745000000
1!
1%
#64750000000
0!
0%
#64755000000
1!
1%
#64760000000
0!
0%
#64765000000
1!
1%
#64770000000
0!
0%
#64775000000
1!
1%
#64780000000
0!
0%
#64785000000
1!
1%
#64790000000
0!
0%
#64795000000
1!
1%
#64800000000
0!
0%
#64805000000
1!
1%
#64810000000
0!
0%
#64815000000
1!
1%
#64820000000
0!
0%
#64825000000
1!
1%
#64830000000
0!
0%
#64835000000
1!
1%
#64840000000
0!
0%
#64845000000
1!
1%
#64850000000
0!
0%
#64855000000
1!
1%
#64860000000
0!
0%
#64865000000
1!
1%
#64870000000
0!
0%
#64875000000
1!
1%
#64880000000
0!
0%
#64885000000
1!
1%
#64890000000
0!
0%
#64895000000
1!
1%
#64900000000
0!
0%
#64905000000
1!
1%
#64910000000
0!
0%
#64915000000
1!
1%
#64920000000
0!
0%
#64925000000
1!
1%
#64930000000
0!
0%
#64935000000
1!
1%
#64940000000
0!
0%
#64945000000
1!
1%
#64950000000
0!
0%
#64955000000
1!
1%
#64960000000
0!
0%
#64965000000
1!
1%
#64970000000
0!
0%
#64975000000
1!
1%
#64980000000
0!
0%
#64985000000
1!
1%
#64990000000
0!
0%
#64995000000
1!
1%
#65000000000
0!
0%
#65005000000
1!
1%
#65010000000
0!
0%
#65015000000
1!
1%
#65020000000
0!
0%
#65025000000
1!
1%
#65030000000
0!
0%
#65035000000
1!
1%
#65040000000
0!
0%
#65045000000
1!
1%
#65050000000
0!
0%
#65055000000
1!
1%
#65060000000
0!
0%
#65065000000
1!
1%
#65070000000
0!
0%
#65075000000
1!
1%
#65080000000
0!
0%
#65085000000
1!
1%
#65090000000
0!
0%
#65095000000
1!
1%
#65100000000
0!
0%
#65105000000
1!
1%
#65110000000
0!
0%
#65115000000
1!
1%
#65120000000
0!
0%
#65125000000
1!
1%
#65130000000
0!
0%
#65135000000
1!
1%
#65140000000
0!
0%
#65145000000
1!
1%
#65150000000
0!
0%
#65155000000
1!
1%
#65160000000
0!
0%
#65165000000
1!
1%
#65170000000
0!
0%
#65175000000
1!
1%
#65180000000
0!
0%
#65185000000
1!
1%
#65190000000
0!
0%
#65195000000
1!
1%
#65200000000
0!
0%
#65205000000
1!
1%
#65210000000
0!
0%
#65215000000
1!
1%
#65220000000
0!
0%
#65225000000
1!
1%
#65230000000
0!
0%
#65235000000
1!
1%
#65240000000
0!
0%
#65245000000
1!
1%
#65250000000
0!
0%
#65255000000
1!
1%
#65260000000
0!
0%
#65265000000
1!
1%
#65270000000
0!
0%
#65275000000
1!
1%
#65280000000
0!
0%
#65285000000
1!
1%
#65290000000
0!
0%
#65295000000
1!
1%
#65300000000
0!
0%
#65305000000
1!
1%
#65310000000
0!
0%
#65315000000
1!
1%
#65320000000
0!
0%
#65325000000
1!
1%
#65330000000
0!
0%
#65335000000
1!
1%
#65340000000
0!
0%
#65345000000
1!
1%
#65350000000
0!
0%
#65355000000
1!
1%
#65360000000
0!
0%
#65365000000
1!
1%
#65370000000
0!
0%
#65375000000
1!
1%
#65380000000
0!
0%
#65385000000
1!
1%
#65390000000
0!
0%
#65395000000
1!
1%
#65400000000
0!
0%
#65405000000
1!
1%
#65410000000
0!
0%
#65415000000
1!
1%
#65420000000
0!
0%
#65425000000
1!
1%
#65430000000
0!
0%
#65435000000
1!
1%
#65440000000
0!
0%
#65445000000
1!
1%
#65450000000
0!
0%
#65455000000
1!
1%
#65460000000
0!
0%
#65465000000
1!
1%
#65470000000
0!
0%
#65475000000
1!
1%
#65480000000
0!
0%
#65485000000
1!
1%
#65490000000
0!
0%
#65495000000
1!
1%
#65500000000
0!
0%
#65505000000
1!
1%
#65510000000
0!
0%
#65515000000
1!
1%
#65520000000
0!
0%
#65525000000
1!
1%
#65530000000
0!
0%
#65535000000
1!
1%
#65540000000
0!
0%
#65545000000
1!
1%
#65550000000
0!
0%
#65555000000
1!
1%
#65560000000
0!
0%
#65565000000
1!
1%
#65570000000
0!
0%
#65575000000
1!
1%
#65580000000
0!
0%
#65585000000
1!
1%
#65590000000
0!
0%
#65595000000
1!
1%
#65600000000
0!
0%
#65605000000
1!
1%
#65610000000
0!
0%
#65615000000
1!
1%
#65620000000
0!
0%
#65625000000
1!
1%
#65630000000
0!
0%
#65635000000
1!
1%
#65640000000
0!
0%
#65645000000
1!
1%
#65650000000
0!
0%
#65655000000
1!
1%
#65660000000
0!
0%
#65665000000
1!
1%
#65670000000
0!
0%
#65675000000
1!
1%
#65680000000
0!
0%
#65685000000
1!
1%
#65690000000
0!
0%
#65695000000
1!
1%
#65700000000
0!
0%
#65705000000
1!
1%
#65710000000
0!
0%
#65715000000
1!
1%
#65720000000
0!
0%
#65725000000
1!
1%
#65730000000
0!
0%
#65735000000
1!
1%
#65740000000
0!
0%
#65745000000
1!
1%
#65750000000
0!
0%
#65755000000
1!
1%
#65760000000
0!
0%
#65765000000
1!
1%
#65770000000
0!
0%
#65775000000
1!
1%
#65780000000
0!
0%
#65785000000
1!
1%
#65790000000
0!
0%
#65795000000
1!
1%
#65800000000
0!
0%
#65805000000
1!
1%
#65810000000
0!
0%
#65815000000
1!
1%
#65820000000
0!
0%
#65825000000
1!
1%
#65830000000
0!
0%
#65835000000
1!
1%
#65840000000
0!
0%
#65845000000
1!
1%
#65850000000
0!
0%
#65855000000
1!
1%
#65860000000
0!
0%
#65865000000
1!
1%
#65870000000
0!
0%
#65875000000
1!
1%
#65880000000
0!
0%
#65885000000
1!
1%
#65890000000
0!
0%
#65895000000
1!
1%
#65900000000
0!
0%
#65905000000
1!
1%
#65910000000
0!
0%
#65915000000
1!
1%
#65920000000
0!
0%
#65925000000
1!
1%
#65930000000
0!
0%
#65935000000
1!
1%
#65940000000
0!
0%
#65945000000
1!
1%
#65950000000
0!
0%
#65955000000
1!
1%
#65960000000
0!
0%
#65965000000
1!
1%
#65970000000
0!
0%
#65975000000
1!
1%
#65980000000
0!
0%
#65985000000
1!
1%
#65990000000
0!
0%
#65995000000
1!
1%
#66000000000
0!
0%
#66005000000
1!
1%
#66010000000
0!
0%
#66015000000
1!
1%
#66020000000
0!
0%
#66025000000
1!
1%
#66030000000
0!
0%
#66035000000
1!
1%
#66040000000
0!
0%
#66045000000
1!
1%
#66050000000
0!
0%
#66055000000
1!
1%
#66060000000
0!
0%
#66065000000
1!
1%
#66070000000
0!
0%
#66075000000
1!
1%
#66080000000
0!
0%
#66085000000
1!
1%
#66090000000
0!
0%
#66095000000
1!
1%
#66100000000
0!
0%
#66105000000
1!
1%
#66110000000
0!
0%
#66115000000
1!
1%
#66120000000
0!
0%
#66125000000
1!
1%
#66130000000
0!
0%
#66135000000
1!
1%
#66140000000
0!
0%
#66145000000
1!
1%
#66150000000
0!
0%
#66155000000
1!
1%
#66160000000
0!
0%
#66165000000
1!
1%
#66170000000
0!
0%
#66175000000
1!
1%
#66180000000
0!
0%
#66185000000
1!
1%
#66190000000
0!
0%
#66195000000
1!
1%
#66200000000
0!
0%
#66205000000
1!
1%
#66210000000
0!
0%
#66215000000
1!
1%
#66220000000
0!
0%
#66225000000
1!
1%
#66230000000
0!
0%
#66235000000
1!
1%
#66240000000
0!
0%
#66245000000
1!
1%
#66250000000
0!
0%
#66255000000
1!
1%
#66260000000
0!
0%
#66265000000
1!
1%
#66270000000
0!
0%
#66275000000
1!
1%
#66280000000
0!
0%
#66285000000
1!
1%
#66290000000
0!
0%
#66295000000
1!
1%
#66300000000
0!
0%
#66305000000
1!
1%
#66310000000
0!
0%
#66315000000
1!
1%
#66320000000
0!
0%
#66325000000
1!
1%
#66330000000
0!
0%
#66335000000
1!
1%
#66340000000
0!
0%
#66345000000
1!
1%
#66350000000
0!
0%
#66355000000
1!
1%
#66360000000
0!
0%
#66365000000
1!
1%
#66370000000
0!
0%
#66375000000
1!
1%
#66380000000
0!
0%
#66385000000
1!
1%
#66390000000
0!
0%
#66395000000
1!
1%
#66400000000
0!
0%
#66405000000
1!
1%
#66410000000
0!
0%
#66415000000
1!
1%
#66420000000
0!
0%
#66425000000
1!
1%
#66430000000
0!
0%
#66435000000
1!
1%
#66440000000
0!
0%
#66445000000
1!
1%
#66450000000
0!
0%
#66455000000
1!
1%
#66460000000
0!
0%
#66465000000
1!
1%
#66470000000
0!
0%
#66475000000
1!
1%
#66480000000
0!
0%
#66485000000
1!
1%
#66490000000
0!
0%
#66495000000
1!
1%
#66500000000
0!
0%
#66505000000
1!
1%
#66510000000
0!
0%
#66515000000
1!
1%
#66520000000
0!
0%
#66525000000
1!
1%
#66530000000
0!
0%
#66535000000
1!
1%
#66540000000
0!
0%
#66545000000
1!
1%
#66550000000
0!
0%
#66555000000
1!
1%
#66560000000
0!
0%
#66565000000
1!
1%
#66570000000
0!
0%
#66575000000
1!
1%
#66580000000
0!
0%
#66585000000
1!
1%
#66590000000
0!
0%
#66595000000
1!
1%
#66600000000
0!
0%
#66605000000
1!
1%
#66610000000
0!
0%
#66615000000
1!
1%
#66620000000
0!
0%
#66625000000
1!
1%
#66630000000
0!
0%
#66635000000
1!
1%
#66640000000
0!
0%
#66645000000
1!
1%
#66650000000
0!
0%
#66655000000
1!
1%
#66660000000
0!
0%
#66665000000
1!
1%
#66670000000
0!
0%
#66675000000
1!
1%
#66680000000
0!
0%
#66685000000
1!
1%
#66690000000
0!
0%
#66695000000
1!
1%
#66700000000
0!
0%
#66705000000
1!
1%
#66710000000
0!
0%
#66715000000
1!
1%
#66720000000
0!
0%
#66725000000
1!
1%
#66730000000
0!
0%
#66735000000
1!
1%
#66740000000
0!
0%
#66745000000
1!
1%
#66750000000
0!
0%
#66755000000
1!
1%
#66760000000
0!
0%
#66765000000
1!
1%
#66770000000
0!
0%
#66775000000
1!
1%
#66780000000
0!
0%
#66785000000
1!
1%
#66790000000
0!
0%
#66795000000
1!
1%
#66800000000
0!
0%
#66805000000
1!
1%
#66810000000
0!
0%
#66815000000
1!
1%
#66820000000
0!
0%
#66825000000
1!
1%
#66830000000
0!
0%
#66835000000
1!
1%
#66840000000
0!
0%
#66845000000
1!
1%
#66850000000
0!
0%
#66855000000
1!
1%
#66860000000
0!
0%
#66865000000
1!
1%
#66870000000
0!
0%
#66875000000
1!
1%
#66880000000
0!
0%
#66885000000
1!
1%
#66890000000
0!
0%
#66895000000
1!
1%
#66900000000
0!
0%
#66905000000
1!
1%
#66910000000
0!
0%
#66915000000
1!
1%
#66920000000
0!
0%
#66925000000
1!
1%
#66930000000
0!
0%
#66935000000
1!
1%
#66940000000
0!
0%
#66945000000
1!
1%
#66950000000
0!
0%
#66955000000
1!
1%
#66960000000
0!
0%
#66965000000
1!
1%
#66970000000
0!
0%
#66975000000
1!
1%
#66980000000
0!
0%
#66985000000
1!
1%
#66990000000
0!
0%
#66995000000
1!
1%
#67000000000
0!
0%
#67005000000
1!
1%
#67010000000
0!
0%
#67015000000
1!
1%
#67020000000
0!
0%
#67025000000
1!
1%
#67030000000
0!
0%
#67035000000
1!
1%
#67040000000
0!
0%
#67045000000
1!
1%
#67050000000
0!
0%
#67055000000
1!
1%
#67060000000
0!
0%
#67065000000
1!
1%
#67070000000
0!
0%
#67075000000
1!
1%
#67080000000
0!
0%
#67085000000
1!
1%
#67090000000
0!
0%
#67095000000
1!
1%
#67100000000
0!
0%
#67105000000
1!
1%
#67110000000
0!
0%
#67115000000
1!
1%
#67120000000
0!
0%
#67125000000
1!
1%
#67130000000
0!
0%
#67135000000
1!
1%
#67140000000
0!
0%
#67145000000
1!
1%
#67150000000
0!
0%
#67155000000
1!
1%
#67160000000
0!
0%
#67165000000
1!
1%
#67170000000
0!
0%
#67175000000
1!
1%
#67180000000
0!
0%
#67185000000
1!
1%
#67190000000
0!
0%
#67195000000
1!
1%
#67200000000
0!
0%
#67205000000
1!
1%
#67210000000
0!
0%
#67215000000
1!
1%
#67220000000
0!
0%
#67225000000
1!
1%
#67230000000
0!
0%
#67235000000
1!
1%
#67240000000
0!
0%
#67245000000
1!
1%
#67250000000
0!
0%
#67255000000
1!
1%
#67260000000
0!
0%
#67265000000
1!
1%
#67270000000
0!
0%
#67275000000
1!
1%
#67280000000
0!
0%
#67285000000
1!
1%
#67290000000
0!
0%
#67295000000
1!
1%
#67300000000
0!
0%
#67305000000
1!
1%
#67310000000
0!
0%
#67315000000
1!
1%
#67320000000
0!
0%
#67325000000
1!
1%
#67330000000
0!
0%
#67335000000
1!
1%
#67340000000
0!
0%
#67345000000
1!
1%
#67350000000
0!
0%
#67355000000
1!
1%
#67360000000
0!
0%
#67365000000
1!
1%
#67370000000
0!
0%
#67375000000
1!
1%
#67380000000
0!
0%
#67385000000
1!
1%
#67390000000
0!
0%
#67395000000
1!
1%
#67400000000
0!
0%
#67405000000
1!
1%
#67410000000
0!
0%
#67415000000
1!
1%
#67420000000
0!
0%
#67425000000
1!
1%
#67430000000
0!
0%
#67435000000
1!
1%
#67440000000
0!
0%
#67445000000
1!
1%
#67450000000
0!
0%
#67455000000
1!
1%
#67460000000
0!
0%
#67465000000
1!
1%
#67470000000
0!
0%
#67475000000
1!
1%
#67480000000
0!
0%
#67485000000
1!
1%
#67490000000
0!
0%
#67495000000
1!
1%
#67500000000
0!
0%
#67505000000
1!
1%
#67510000000
0!
0%
#67515000000
1!
1%
#67520000000
0!
0%
#67525000000
1!
1%
#67530000000
0!
0%
#67535000000
1!
1%
#67540000000
0!
0%
#67545000000
1!
1%
#67550000000
0!
0%
#67555000000
1!
1%
#67560000000
0!
0%
#67565000000
1!
1%
#67570000000
0!
0%
#67575000000
1!
1%
#67580000000
0!
0%
#67585000000
1!
1%
#67590000000
0!
0%
#67595000000
1!
1%
#67600000000
0!
0%
#67605000000
1!
1%
#67610000000
0!
0%
#67615000000
1!
1%
#67620000000
0!
0%
#67625000000
1!
1%
#67630000000
0!
0%
#67635000000
1!
1%
#67640000000
0!
0%
#67645000000
1!
1%
#67650000000
0!
0%
#67655000000
1!
1%
#67660000000
0!
0%
#67665000000
1!
1%
#67670000000
0!
0%
#67675000000
1!
1%
#67680000000
0!
0%
#67685000000
1!
1%
#67690000000
0!
0%
#67695000000
1!
1%
#67700000000
0!
0%
#67705000000
1!
1%
#67710000000
0!
0%
#67715000000
1!
1%
#67720000000
0!
0%
#67725000000
1!
1%
#67730000000
0!
0%
#67735000000
1!
1%
#67740000000
0!
0%
#67745000000
1!
1%
#67750000000
0!
0%
#67755000000
1!
1%
#67760000000
0!
0%
#67765000000
1!
1%
#67770000000
0!
0%
#67775000000
1!
1%
#67780000000
0!
0%
#67785000000
1!
1%
#67790000000
0!
0%
#67795000000
1!
1%
#67800000000
0!
0%
#67805000000
1!
1%
#67810000000
0!
0%
#67815000000
1!
1%
#67820000000
0!
0%
#67825000000
1!
1%
#67830000000
0!
0%
#67835000000
1!
1%
#67840000000
0!
0%
#67845000000
1!
1%
#67850000000
0!
0%
#67855000000
1!
1%
#67860000000
0!
0%
#67865000000
1!
1%
#67870000000
0!
0%
#67875000000
1!
1%
#67880000000
0!
0%
#67885000000
1!
1%
#67890000000
0!
0%
#67895000000
1!
1%
#67900000000
0!
0%
#67905000000
1!
1%
#67910000000
0!
0%
#67915000000
1!
1%
#67920000000
0!
0%
#67925000000
1!
1%
#67930000000
0!
0%
#67935000000
1!
1%
#67940000000
0!
0%
#67945000000
1!
1%
#67950000000
0!
0%
#67955000000
1!
1%
#67960000000
0!
0%
#67965000000
1!
1%
#67970000000
0!
0%
#67975000000
1!
1%
#67980000000
0!
0%
#67985000000
1!
1%
#67990000000
0!
0%
#67995000000
1!
1%
#68000000000
0!
0%
#68005000000
1!
1%
#68010000000
0!
0%
#68015000000
1!
1%
#68020000000
0!
0%
#68025000000
1!
1%
#68030000000
0!
0%
#68035000000
1!
1%
#68040000000
0!
0%
#68045000000
1!
1%
#68050000000
0!
0%
#68055000000
1!
1%
#68060000000
0!
0%
#68065000000
1!
1%
#68070000000
0!
0%
#68075000000
1!
1%
#68080000000
0!
0%
#68085000000
1!
1%
#68090000000
0!
0%
#68095000000
1!
1%
#68100000000
0!
0%
#68105000000
1!
1%
#68110000000
0!
0%
#68115000000
1!
1%
#68120000000
0!
0%
#68125000000
1!
1%
#68130000000
0!
0%
#68135000000
1!
1%
#68140000000
0!
0%
#68145000000
1!
1%
#68150000000
0!
0%
#68155000000
1!
1%
#68160000000
0!
0%
#68165000000
1!
1%
#68170000000
0!
0%
#68175000000
1!
1%
#68180000000
0!
0%
#68185000000
1!
1%
#68190000000
0!
0%
#68195000000
1!
1%
#68200000000
0!
0%
#68205000000
1!
1%
#68210000000
0!
0%
#68215000000
1!
1%
#68220000000
0!
0%
#68225000000
1!
1%
#68230000000
0!
0%
#68235000000
1!
1%
#68240000000
0!
0%
#68245000000
1!
1%
#68250000000
0!
0%
#68255000000
1!
1%
#68260000000
0!
0%
#68265000000
1!
1%
#68270000000
0!
0%
#68275000000
1!
1%
#68280000000
0!
0%
#68285000000
1!
1%
#68290000000
0!
0%
#68295000000
1!
1%
#68300000000
0!
0%
#68305000000
1!
1%
#68310000000
0!
0%
#68315000000
1!
1%
#68320000000
0!
0%
#68325000000
1!
1%
#68330000000
0!
0%
#68335000000
1!
1%
#68340000000
0!
0%
#68345000000
1!
1%
#68350000000
0!
0%
#68355000000
1!
1%
#68360000000
0!
0%
#68365000000
1!
1%
#68370000000
0!
0%
#68375000000
1!
1%
#68380000000
0!
0%
#68385000000
1!
1%
#68390000000
0!
0%
#68395000000
1!
1%
#68400000000
0!
0%
#68405000000
1!
1%
#68410000000
0!
0%
#68415000000
1!
1%
#68420000000
0!
0%
#68425000000
1!
1%
#68430000000
0!
0%
#68435000000
1!
1%
#68440000000
0!
0%
#68445000000
1!
1%
#68450000000
0!
0%
#68455000000
1!
1%
#68460000000
0!
0%
#68465000000
1!
1%
#68470000000
0!
0%
#68475000000
1!
1%
#68480000000
0!
0%
#68485000000
1!
1%
#68490000000
0!
0%
#68495000000
1!
1%
#68500000000
0!
0%
#68505000000
1!
1%
#68510000000
0!
0%
#68515000000
1!
1%
#68520000000
0!
0%
#68525000000
1!
1%
#68530000000
0!
0%
#68535000000
1!
1%
#68540000000
0!
0%
#68545000000
1!
1%
#68550000000
0!
0%
#68555000000
1!
1%
#68560000000
0!
0%
#68565000000
1!
1%
#68570000000
0!
0%
#68575000000
1!
1%
#68580000000
0!
0%
#68585000000
1!
1%
#68590000000
0!
0%
#68595000000
1!
1%
#68600000000
0!
0%
#68605000000
1!
1%
#68610000000
0!
0%
#68615000000
1!
1%
#68620000000
0!
0%
#68625000000
1!
1%
#68630000000
0!
0%
#68635000000
1!
1%
#68640000000
0!
0%
#68645000000
1!
1%
#68650000000
0!
0%
#68655000000
1!
1%
#68660000000
0!
0%
#68665000000
1!
1%
#68670000000
0!
0%
#68675000000
1!
1%
#68680000000
0!
0%
#68685000000
1!
1%
#68690000000
0!
0%
#68695000000
1!
1%
#68700000000
0!
0%
#68705000000
1!
1%
#68710000000
0!
0%
#68715000000
1!
1%
#68720000000
0!
0%
#68725000000
1!
1%
#68730000000
0!
0%
#68735000000
1!
1%
#68740000000
0!
0%
#68745000000
1!
1%
#68750000000
0!
0%
#68755000000
1!
1%
#68760000000
0!
0%
#68765000000
1!
1%
#68770000000
0!
0%
#68775000000
1!
1%
#68780000000
0!
0%
#68785000000
1!
1%
#68790000000
0!
0%
#68795000000
1!
1%
#68800000000
0!
0%
#68805000000
1!
1%
#68810000000
0!
0%
#68815000000
1!
1%
#68820000000
0!
0%
#68825000000
1!
1%
#68830000000
0!
0%
#68835000000
1!
1%
#68840000000
0!
0%
#68845000000
1!
1%
#68850000000
0!
0%
#68855000000
1!
1%
#68860000000
0!
0%
#68865000000
1!
1%
#68870000000
0!
0%
#68875000000
1!
1%
#68880000000
0!
0%
#68885000000
1!
1%
#68890000000
0!
0%
#68895000000
1!
1%
#68900000000
0!
0%
#68905000000
1!
1%
#68910000000
0!
0%
#68915000000
1!
1%
#68920000000
0!
0%
#68925000000
1!
1%
#68930000000
0!
0%
#68935000000
1!
1%
#68940000000
0!
0%
#68945000000
1!
1%
#68950000000
0!
0%
#68955000000
1!
1%
#68960000000
0!
0%
#68965000000
1!
1%
#68970000000
0!
0%
#68975000000
1!
1%
#68980000000
0!
0%
#68985000000
1!
1%
#68990000000
0!
0%
#68995000000
1!
1%
#69000000000
0!
0%
#69005000000
1!
1%
#69010000000
0!
0%
#69015000000
1!
1%
#69020000000
0!
0%
#69025000000
1!
1%
#69030000000
0!
0%
#69035000000
1!
1%
#69040000000
0!
0%
#69045000000
1!
1%
#69050000000
0!
0%
#69055000000
1!
1%
#69060000000
0!
0%
#69065000000
1!
1%
#69070000000
0!
0%
#69075000000
1!
1%
#69080000000
0!
0%
#69085000000
1!
1%
#69090000000
0!
0%
#69095000000
1!
1%
#69100000000
0!
0%
#69105000000
1!
1%
#69110000000
0!
0%
#69115000000
1!
1%
#69120000000
0!
0%
#69125000000
1!
1%
#69130000000
0!
0%
#69135000000
1!
1%
#69140000000
0!
0%
#69145000000
1!
1%
#69150000000
0!
0%
#69155000000
1!
1%
#69160000000
0!
0%
#69165000000
1!
1%
#69170000000
0!
0%
#69175000000
1!
1%
#69180000000
0!
0%
#69185000000
1!
1%
#69190000000
0!
0%
#69195000000
1!
1%
#69200000000
0!
0%
#69205000000
1!
1%
#69210000000
0!
0%
#69215000000
1!
1%
#69220000000
0!
0%
#69225000000
1!
1%
#69230000000
0!
0%
#69235000000
1!
1%
#69240000000
0!
0%
#69245000000
1!
1%
#69250000000
0!
0%
#69255000000
1!
1%
#69260000000
0!
0%
#69265000000
1!
1%
#69270000000
0!
0%
#69275000000
1!
1%
#69280000000
0!
0%
#69285000000
1!
1%
#69290000000
0!
0%
#69295000000
1!
1%
#69300000000
0!
0%
#69305000000
1!
1%
#69310000000
0!
0%
#69315000000
1!
1%
#69320000000
0!
0%
#69325000000
1!
1%
#69330000000
0!
0%
#69335000000
1!
1%
#69340000000
0!
0%
#69345000000
1!
1%
#69350000000
0!
0%
#69355000000
1!
1%
#69360000000
0!
0%
#69365000000
1!
1%
#69370000000
0!
0%
#69375000000
1!
1%
#69380000000
0!
0%
#69385000000
1!
1%
#69390000000
0!
0%
#69395000000
1!
1%
#69400000000
0!
0%
#69405000000
1!
1%
#69410000000
0!
0%
#69415000000
1!
1%
#69420000000
0!
0%
#69425000000
1!
1%
#69430000000
0!
0%
#69435000000
1!
1%
#69440000000
0!
0%
#69445000000
1!
1%
#69450000000
0!
0%
#69455000000
1!
1%
#69460000000
0!
0%
#69465000000
1!
1%
#69470000000
0!
0%
#69475000000
1!
1%
#69480000000
0!
0%
#69485000000
1!
1%
#69490000000
0!
0%
#69495000000
1!
1%
#69500000000
0!
0%
#69505000000
1!
1%
#69510000000
0!
0%
#69515000000
1!
1%
#69520000000
0!
0%
#69525000000
1!
1%
#69530000000
0!
0%
#69535000000
1!
1%
#69540000000
0!
0%
#69545000000
1!
1%
#69550000000
0!
0%
#69555000000
1!
1%
#69560000000
0!
0%
#69565000000
1!
1%
#69570000000
0!
0%
#69575000000
1!
1%
#69580000000
0!
0%
#69585000000
1!
1%
#69590000000
0!
0%
#69595000000
1!
1%
#69600000000
0!
0%
#69605000000
1!
1%
#69610000000
0!
0%
#69615000000
1!
1%
#69620000000
0!
0%
#69625000000
1!
1%
#69630000000
0!
0%
#69635000000
1!
1%
#69640000000
0!
0%
#69645000000
1!
1%
#69650000000
0!
0%
#69655000000
1!
1%
#69660000000
0!
0%
#69665000000
1!
1%
#69670000000
0!
0%
#69675000000
1!
1%
#69680000000
0!
0%
#69685000000
1!
1%
#69690000000
0!
0%
#69695000000
1!
1%
#69700000000
0!
0%
#69705000000
1!
1%
#69710000000
0!
0%
#69715000000
1!
1%
#69720000000
0!
0%
#69725000000
1!
1%
#69730000000
0!
0%
#69735000000
1!
1%
#69740000000
0!
0%
#69745000000
1!
1%
#69750000000
0!
0%
#69755000000
1!
1%
#69760000000
0!
0%
#69765000000
1!
1%
#69770000000
0!
0%
#69775000000
1!
1%
#69780000000
0!
0%
#69785000000
1!
1%
#69790000000
0!
0%
#69795000000
1!
1%
#69800000000
0!
0%
#69805000000
1!
1%
#69810000000
0!
0%
#69815000000
1!
1%
#69820000000
0!
0%
#69825000000
1!
1%
#69830000000
0!
0%
#69835000000
1!
1%
#69840000000
0!
0%
#69845000000
1!
1%
#69850000000
0!
0%
#69855000000
1!
1%
#69860000000
0!
0%
#69865000000
1!
1%
#69870000000
0!
0%
#69875000000
1!
1%
#69880000000
0!
0%
#69885000000
1!
1%
#69890000000
0!
0%
#69895000000
1!
1%
#69900000000
0!
0%
#69905000000
1!
1%
#69910000000
0!
0%
#69915000000
1!
1%
#69920000000
0!
0%
#69925000000
1!
1%
#69930000000
0!
0%
#69935000000
1!
1%
#69940000000
0!
0%
#69945000000
1!
1%
#69950000000
0!
0%
#69955000000
1!
1%
#69960000000
0!
0%
#69965000000
1!
1%
#69970000000
0!
0%
#69975000000
1!
1%
#69980000000
0!
0%
#69985000000
1!
1%
#69990000000
0!
0%
#69995000000
1!
1%
#70000000000
0!
0%
#70005000000
1!
1%
#70010000000
0!
0%
#70015000000
1!
1%
#70020000000
0!
0%
#70025000000
1!
1%
#70030000000
0!
0%
#70035000000
1!
1%
#70040000000
0!
0%
#70045000000
1!
1%
#70050000000
0!
0%
#70055000000
1!
1%
#70060000000
0!
0%
#70065000000
1!
1%
#70070000000
0!
0%
#70075000000
1!
1%
#70080000000
0!
0%
#70085000000
1!
1%
#70090000000
0!
0%
#70095000000
1!
1%
#70100000000
0!
0%
#70105000000
1!
1%
#70110000000
0!
0%
#70115000000
1!
1%
#70120000000
0!
0%
#70125000000
1!
1%
#70130000000
0!
0%
#70135000000
1!
1%
#70140000000
0!
0%
#70145000000
1!
1%
#70150000000
0!
0%
#70155000000
1!
1%
#70160000000
0!
0%
#70165000000
1!
1%
#70170000000
0!
0%
#70175000000
1!
1%
#70180000000
0!
0%
#70185000000
1!
1%
#70190000000
0!
0%
#70195000000
1!
1%
#70200000000
0!
0%
#70205000000
1!
1%
#70210000000
0!
0%
#70215000000
1!
1%
#70220000000
0!
0%
#70225000000
1!
1%
#70230000000
0!
0%
#70235000000
1!
1%
#70240000000
0!
0%
#70245000000
1!
1%
#70250000000
0!
0%
#70255000000
1!
1%
#70260000000
0!
0%
#70265000000
1!
1%
#70270000000
0!
0%
#70275000000
1!
1%
#70280000000
0!
0%
#70285000000
1!
1%
#70290000000
0!
0%
#70295000000
1!
1%
#70300000000
0!
0%
#70305000000
1!
1%
#70310000000
0!
0%
#70315000000
1!
1%
#70320000000
0!
0%
#70325000000
1!
1%
#70330000000
0!
0%
#70335000000
1!
1%
#70340000000
0!
0%
#70345000000
1!
1%
#70350000000
0!
0%
#70355000000
1!
1%
#70360000000
0!
0%
#70365000000
1!
1%
#70370000000
0!
0%
#70375000000
1!
1%
#70380000000
0!
0%
#70385000000
1!
1%
#70390000000
0!
0%
#70395000000
1!
1%
#70400000000
0!
0%
#70405000000
1!
1%
#70410000000
0!
0%
#70415000000
1!
1%
#70420000000
0!
0%
#70425000000
1!
1%
#70430000000
0!
0%
#70435000000
1!
1%
#70440000000
0!
0%
#70445000000
1!
1%
#70450000000
0!
0%
#70455000000
1!
1%
#70460000000
0!
0%
#70465000000
1!
1%
#70470000000
0!
0%
#70475000000
1!
1%
#70480000000
0!
0%
#70485000000
1!
1%
#70490000000
0!
0%
#70495000000
1!
1%
#70500000000
0!
0%
#70505000000
1!
1%
#70510000000
0!
0%
#70515000000
1!
1%
#70520000000
0!
0%
#70525000000
1!
1%
#70530000000
0!
0%
#70535000000
1!
1%
#70540000000
0!
0%
#70545000000
1!
1%
#70550000000
0!
0%
#70555000000
1!
1%
#70560000000
0!
0%
#70565000000
1!
1%
#70570000000
0!
0%
#70575000000
1!
1%
#70580000000
0!
0%
#70585000000
1!
1%
#70590000000
0!
0%
#70595000000
1!
1%
#70600000000
0!
0%
#70605000000
1!
1%
#70610000000
0!
0%
#70615000000
1!
1%
#70620000000
0!
0%
#70625000000
1!
1%
#70630000000
0!
0%
#70635000000
1!
1%
#70640000000
0!
0%
#70645000000
1!
1%
#70650000000
0!
0%
#70655000000
1!
1%
#70660000000
0!
0%
#70665000000
1!
1%
#70670000000
0!
0%
#70675000000
1!
1%
#70680000000
0!
0%
#70685000000
1!
1%
#70690000000
0!
0%
#70695000000
1!
1%
#70700000000
0!
0%
#70705000000
1!
1%
#70710000000
0!
0%
#70715000000
1!
1%
#70720000000
0!
0%
#70725000000
1!
1%
#70730000000
0!
0%
#70735000000
1!
1%
#70740000000
0!
0%
#70745000000
1!
1%
#70750000000
0!
0%
#70755000000
1!
1%
#70760000000
0!
0%
#70765000000
1!
1%
#70770000000
0!
0%
#70775000000
1!
1%
#70780000000
0!
0%
#70785000000
1!
1%
#70790000000
0!
0%
#70795000000
1!
1%
#70800000000
0!
0%
#70805000000
1!
1%
#70810000000
0!
0%
#70815000000
1!
1%
#70820000000
0!
0%
#70825000000
1!
1%
#70830000000
0!
0%
#70835000000
1!
1%
#70840000000
0!
0%
#70845000000
1!
1%
#70850000000
0!
0%
#70855000000
1!
1%
#70860000000
0!
0%
#70865000000
1!
1%
#70870000000
0!
0%
#70875000000
1!
1%
#70880000000
0!
0%
#70885000000
1!
1%
#70890000000
0!
0%
#70895000000
1!
1%
#70900000000
0!
0%
#70905000000
1!
1%
#70910000000
0!
0%
#70915000000
1!
1%
#70920000000
0!
0%
#70925000000
1!
1%
#70930000000
0!
0%
#70935000000
1!
1%
#70940000000
0!
0%
#70945000000
1!
1%
#70950000000
0!
0%
#70955000000
1!
1%
#70960000000
0!
0%
#70965000000
1!
1%
#70970000000
0!
0%
#70975000000
1!
1%
#70980000000
0!
0%
#70985000000
1!
1%
#70990000000
0!
0%
#70995000000
1!
1%
#71000000000
0!
0%
#71005000000
1!
1%
#71010000000
0!
0%
#71015000000
1!
1%
#71020000000
0!
0%
#71025000000
1!
1%
#71030000000
0!
0%
#71035000000
1!
1%
#71040000000
0!
0%
#71045000000
1!
1%
#71050000000
0!
0%
#71055000000
1!
1%
#71060000000
0!
0%
#71065000000
1!
1%
#71070000000
0!
0%
#71075000000
1!
1%
#71080000000
0!
0%
#71085000000
1!
1%
#71090000000
0!
0%
#71095000000
1!
1%
#71100000000
0!
0%
#71105000000
1!
1%
#71110000000
0!
0%
#71115000000
1!
1%
#71120000000
0!
0%
#71125000000
1!
1%
#71130000000
0!
0%
#71135000000
1!
1%
#71140000000
0!
0%
#71145000000
1!
1%
#71150000000
0!
0%
#71155000000
1!
1%
#71160000000
0!
0%
#71165000000
1!
1%
#71170000000
0!
0%
#71175000000
1!
1%
#71180000000
0!
0%
#71185000000
1!
1%
#71190000000
0!
0%
#71195000000
1!
1%
#71200000000
0!
0%
#71205000000
1!
1%
#71210000000
0!
0%
#71215000000
1!
1%
#71220000000
0!
0%
#71225000000
1!
1%
#71230000000
0!
0%
#71235000000
1!
1%
#71240000000
0!
0%
#71245000000
1!
1%
#71250000000
0!
0%
#71255000000
1!
1%
#71260000000
0!
0%
#71265000000
1!
1%
#71270000000
0!
0%
#71275000000
1!
1%
#71280000000
0!
0%
#71285000000
1!
1%
#71290000000
0!
0%
#71295000000
1!
1%
#71300000000
0!
0%
#71305000000
1!
1%
#71310000000
0!
0%
#71315000000
1!
1%
#71320000000
0!
0%
#71325000000
1!
1%
#71330000000
0!
0%
#71335000000
1!
1%
#71340000000
0!
0%
#71345000000
1!
1%
#71350000000
0!
0%
#71355000000
1!
1%
#71360000000
0!
0%
#71365000000
1!
1%
#71370000000
0!
0%
#71375000000
1!
1%
#71380000000
0!
0%
#71385000000
1!
1%
#71390000000
0!
0%
#71395000000
1!
1%
#71400000000
0!
0%
#71405000000
1!
1%
#71410000000
0!
0%
#71415000000
1!
1%
#71420000000
0!
0%
#71425000000
1!
1%
#71430000000
0!
0%
#71435000000
1!
1%
#71440000000
0!
0%
#71445000000
1!
1%
#71450000000
0!
0%
#71455000000
1!
1%
#71460000000
0!
0%
#71465000000
1!
1%
#71470000000
0!
0%
#71475000000
1!
1%
#71480000000
0!
0%
#71485000000
1!
1%
#71490000000
0!
0%
#71495000000
1!
1%
#71500000000
0!
0%
#71505000000
1!
1%
#71510000000
0!
0%
#71515000000
1!
1%
#71520000000
0!
0%
#71525000000
1!
1%
#71530000000
0!
0%
#71535000000
1!
1%
#71540000000
0!
0%
#71545000000
1!
1%
#71550000000
0!
0%
#71555000000
1!
1%
#71560000000
0!
0%
#71565000000
1!
1%
#71570000000
0!
0%
#71575000000
1!
1%
#71580000000
0!
0%
#71585000000
1!
1%
#71590000000
0!
0%
#71595000000
1!
1%
#71600000000
0!
0%
#71605000000
1!
1%
#71610000000
0!
0%
#71615000000
1!
1%
#71620000000
0!
0%
#71625000000
1!
1%
#71630000000
0!
0%
#71635000000
1!
1%
#71640000000
0!
0%
#71645000000
1!
1%
#71650000000
0!
0%
#71655000000
1!
1%
#71660000000
0!
0%
#71665000000
1!
1%
#71670000000
0!
0%
#71675000000
1!
1%
#71680000000
0!
0%
#71685000000
1!
1%
#71690000000
0!
0%
#71695000000
1!
1%
#71700000000
0!
0%
#71705000000
1!
1%
#71710000000
0!
0%
#71715000000
1!
1%
#71720000000
0!
0%
#71725000000
1!
1%
#71730000000
0!
0%
#71735000000
1!
1%
#71740000000
0!
0%
#71745000000
1!
1%
#71750000000
0!
0%
#71755000000
1!
1%
#71760000000
0!
0%
#71765000000
1!
1%
#71770000000
0!
0%
#71775000000
1!
1%
#71780000000
0!
0%
#71785000000
1!
1%
#71790000000
0!
0%
#71795000000
1!
1%
#71800000000
0!
0%
#71805000000
1!
1%
#71810000000
0!
0%
#71815000000
1!
1%
#71820000000
0!
0%
#71825000000
1!
1%
#71830000000
0!
0%
#71835000000
1!
1%
#71840000000
0!
0%
#71845000000
1!
1%
#71850000000
0!
0%
#71855000000
1!
1%
#71860000000
0!
0%
#71865000000
1!
1%
#71870000000
0!
0%
#71875000000
1!
1%
#71880000000
0!
0%
#71885000000
1!
1%
#71890000000
0!
0%
#71895000000
1!
1%
#71900000000
0!
0%
#71905000000
1!
1%
#71910000000
0!
0%
#71915000000
1!
1%
#71920000000
0!
0%
#71925000000
1!
1%
#71930000000
0!
0%
#71935000000
1!
1%
#71940000000
0!
0%
#71945000000
1!
1%
#71950000000
0!
0%
#71955000000
1!
1%
#71960000000
0!
0%
#71965000000
1!
1%
#71970000000
0!
0%
#71975000000
1!
1%
#71980000000
0!
0%
#71985000000
1!
1%
#71990000000
0!
0%
#71995000000
1!
1%
#72000000000
0!
0%
#72005000000
1!
1%
#72010000000
0!
0%
#72015000000
1!
1%
#72020000000
0!
0%
#72025000000
1!
1%
#72030000000
0!
0%
#72035000000
1!
1%
#72040000000
0!
0%
#72045000000
1!
1%
#72050000000
0!
0%
#72055000000
1!
1%
#72060000000
0!
0%
#72065000000
1!
1%
#72070000000
0!
0%
#72075000000
1!
1%
#72080000000
0!
0%
#72085000000
1!
1%
#72090000000
0!
0%
#72095000000
1!
1%
#72100000000
0!
0%
#72105000000
1!
1%
#72110000000
0!
0%
#72115000000
1!
1%
#72120000000
0!
0%
#72125000000
1!
1%
#72130000000
0!
0%
#72135000000
1!
1%
#72140000000
0!
0%
#72145000000
1!
1%
#72150000000
0!
0%
#72155000000
1!
1%
#72160000000
0!
0%
#72165000000
1!
1%
#72170000000
0!
0%
#72175000000
1!
1%
#72180000000
0!
0%
#72185000000
1!
1%
#72190000000
0!
0%
#72195000000
1!
1%
#72200000000
0!
0%
#72205000000
1!
1%
#72210000000
0!
0%
#72215000000
1!
1%
#72220000000
0!
0%
#72225000000
1!
1%
#72230000000
0!
0%
#72235000000
1!
1%
#72240000000
0!
0%
#72245000000
1!
1%
#72250000000
0!
0%
#72255000000
1!
1%
#72260000000
0!
0%
#72265000000
1!
1%
#72270000000
0!
0%
#72275000000
1!
1%
#72280000000
0!
0%
#72285000000
1!
1%
#72290000000
0!
0%
#72295000000
1!
1%
#72300000000
0!
0%
#72305000000
1!
1%
#72310000000
0!
0%
#72315000000
1!
1%
#72320000000
0!
0%
#72325000000
1!
1%
#72330000000
0!
0%
#72335000000
1!
1%
#72340000000
0!
0%
#72345000000
1!
1%
#72350000000
0!
0%
#72355000000
1!
1%
#72360000000
0!
0%
#72365000000
1!
1%
#72370000000
0!
0%
#72375000000
1!
1%
#72380000000
0!
0%
#72385000000
1!
1%
#72390000000
0!
0%
#72395000000
1!
1%
#72400000000
0!
0%
#72405000000
1!
1%
#72410000000
0!
0%
#72415000000
1!
1%
#72420000000
0!
0%
#72425000000
1!
1%
#72430000000
0!
0%
#72435000000
1!
1%
#72440000000
0!
0%
#72445000000
1!
1%
#72450000000
0!
0%
#72455000000
1!
1%
#72460000000
0!
0%
#72465000000
1!
1%
#72470000000
0!
0%
#72475000000
1!
1%
#72480000000
0!
0%
#72485000000
1!
1%
#72490000000
0!
0%
#72495000000
1!
1%
#72500000000
0!
0%
#72505000000
1!
1%
#72510000000
0!
0%
#72515000000
1!
1%
#72520000000
0!
0%
#72525000000
1!
1%
#72530000000
0!
0%
#72535000000
1!
1%
#72540000000
0!
0%
#72545000000
1!
1%
#72550000000
0!
0%
#72555000000
1!
1%
#72560000000
0!
0%
#72565000000
1!
1%
#72570000000
0!
0%
#72575000000
1!
1%
#72580000000
0!
0%
#72585000000
1!
1%
#72590000000
0!
0%
#72595000000
1!
1%
#72600000000
0!
0%
#72605000000
1!
1%
#72610000000
0!
0%
#72615000000
1!
1%
#72620000000
0!
0%
#72625000000
1!
1%
#72630000000
0!
0%
#72635000000
1!
1%
#72640000000
0!
0%
#72645000000
1!
1%
#72650000000
0!
0%
#72655000000
1!
1%
#72660000000
0!
0%
#72665000000
1!
1%
#72670000000
0!
0%
#72675000000
1!
1%
#72680000000
0!
0%
#72685000000
1!
1%
#72690000000
0!
0%
#72695000000
1!
1%
#72700000000
0!
0%
#72705000000
1!
1%
#72710000000
0!
0%
#72715000000
1!
1%
#72720000000
0!
0%
#72725000000
1!
1%
#72730000000
0!
0%
#72735000000
1!
1%
#72740000000
0!
0%
#72745000000
1!
1%
#72750000000
0!
0%
#72755000000
1!
1%
#72760000000
0!
0%
#72765000000
1!
1%
#72770000000
0!
0%
#72775000000
1!
1%
#72780000000
0!
0%
#72785000000
1!
1%
#72790000000
0!
0%
#72795000000
1!
1%
#72800000000
0!
0%
#72805000000
1!
1%
#72810000000
0!
0%
#72815000000
1!
1%
#72820000000
0!
0%
#72825000000
1!
1%
#72830000000
0!
0%
#72835000000
1!
1%
#72840000000
0!
0%
#72845000000
1!
1%
#72850000000
0!
0%
#72855000000
1!
1%
#72860000000
0!
0%
#72865000000
1!
1%
#72870000000
0!
0%
#72875000000
1!
1%
#72880000000
0!
0%
#72885000000
1!
1%
#72890000000
0!
0%
#72895000000
1!
1%
#72900000000
0!
0%
#72905000000
1!
1%
#72910000000
0!
0%
#72915000000
1!
1%
#72920000000
0!
0%
#72925000000
1!
1%
#72930000000
0!
0%
#72935000000
1!
1%
#72940000000
0!
0%
#72945000000
1!
1%
#72950000000
0!
0%
#72955000000
1!
1%
#72960000000
0!
0%
#72965000000
1!
1%
#72970000000
0!
0%
#72975000000
1!
1%
#72980000000
0!
0%
#72985000000
1!
1%
#72990000000
0!
0%
#72995000000
1!
1%
#73000000000
0!
0%
#73005000000
1!
1%
#73010000000
0!
0%
#73015000000
1!
1%
#73020000000
0!
0%
#73025000000
1!
1%
#73030000000
0!
0%
#73035000000
1!
1%
#73040000000
0!
0%
#73045000000
1!
1%
#73050000000
0!
0%
#73055000000
1!
1%
#73060000000
0!
0%
#73065000000
1!
1%
#73070000000
0!
0%
#73075000000
1!
1%
#73080000000
0!
0%
#73085000000
1!
1%
#73090000000
0!
0%
#73095000000
1!
1%
#73100000000
0!
0%
#73105000000
1!
1%
#73110000000
0!
0%
#73115000000
1!
1%
#73120000000
0!
0%
#73125000000
1!
1%
#73130000000
0!
0%
#73135000000
1!
1%
#73140000000
0!
0%
#73145000000
1!
1%
#73150000000
0!
0%
#73155000000
1!
1%
#73160000000
0!
0%
#73165000000
1!
1%
#73170000000
0!
0%
#73175000000
1!
1%
#73180000000
0!
0%
#73185000000
1!
1%
#73190000000
0!
0%
#73195000000
1!
1%
#73200000000
0!
0%
#73205000000
1!
1%
#73210000000
0!
0%
#73215000000
1!
1%
#73220000000
0!
0%
#73225000000
1!
1%
#73230000000
0!
0%
#73235000000
1!
1%
#73240000000
0!
0%
#73245000000
1!
1%
#73250000000
0!
0%
#73255000000
1!
1%
#73260000000
0!
0%
#73265000000
1!
1%
#73270000000
0!
0%
#73275000000
1!
1%
#73280000000
0!
0%
#73285000000
1!
1%
#73290000000
0!
0%
#73295000000
1!
1%
#73300000000
0!
0%
#73305000000
1!
1%
#73310000000
0!
0%
#73315000000
1!
1%
#73320000000
0!
0%
#73325000000
1!
1%
#73330000000
0!
0%
#73335000000
1!
1%
#73340000000
0!
0%
#73345000000
1!
1%
#73350000000
0!
0%
#73355000000
1!
1%
#73360000000
0!
0%
#73365000000
1!
1%
#73370000000
0!
0%
#73375000000
1!
1%
#73380000000
0!
0%
#73385000000
1!
1%
#73390000000
0!
0%
#73395000000
1!
1%
#73400000000
0!
0%
#73405000000
1!
1%
#73410000000
0!
0%
#73415000000
1!
1%
#73420000000
0!
0%
#73425000000
1!
1%
#73430000000
0!
0%
#73435000000
1!
1%
#73440000000
0!
0%
#73445000000
1!
1%
#73450000000
0!
0%
#73455000000
1!
1%
#73460000000
0!
0%
#73465000000
1!
1%
#73470000000
0!
0%
#73475000000
1!
1%
#73480000000
0!
0%
#73485000000
1!
1%
#73490000000
0!
0%
#73495000000
1!
1%
#73500000000
0!
0%
#73505000000
1!
1%
#73510000000
0!
0%
#73515000000
1!
1%
#73520000000
0!
0%
#73525000000
1!
1%
#73530000000
0!
0%
#73535000000
1!
1%
#73540000000
0!
0%
#73545000000
1!
1%
#73550000000
0!
0%
#73555000000
1!
1%
#73560000000
0!
0%
#73565000000
1!
1%
#73570000000
0!
0%
#73575000000
1!
1%
#73580000000
0!
0%
#73585000000
1!
1%
#73590000000
0!
0%
#73595000000
1!
1%
#73600000000
0!
0%
#73605000000
1!
1%
#73610000000
0!
0%
#73615000000
1!
1%
#73620000000
0!
0%
#73625000000
1!
1%
#73630000000
0!
0%
#73635000000
1!
1%
#73640000000
0!
0%
#73645000000
1!
1%
#73650000000
0!
0%
#73655000000
1!
1%
#73660000000
0!
0%
#73665000000
1!
1%
#73670000000
0!
0%
#73675000000
1!
1%
#73680000000
0!
0%
#73685000000
1!
1%
#73690000000
0!
0%
#73695000000
1!
1%
#73700000000
0!
0%
#73705000000
1!
1%
#73710000000
0!
0%
#73715000000
1!
1%
#73720000000
0!
0%
#73725000000
1!
1%
#73730000000
0!
0%
#73735000000
1!
1%
#73740000000
0!
0%
#73745000000
1!
1%
#73750000000
0!
0%
#73755000000
1!
1%
#73760000000
0!
0%
#73765000000
1!
1%
#73770000000
0!
0%
#73775000000
1!
1%
#73780000000
0!
0%
#73785000000
1!
1%
#73790000000
0!
0%
#73795000000
1!
1%
#73800000000
0!
0%
#73805000000
1!
1%
#73810000000
0!
0%
#73815000000
1!
1%
#73820000000
0!
0%
#73825000000
1!
1%
#73830000000
0!
0%
#73835000000
1!
1%
#73840000000
0!
0%
#73845000000
1!
1%
#73850000000
0!
0%
#73855000000
1!
1%
#73860000000
0!
0%
#73865000000
1!
1%
#73870000000
0!
0%
#73875000000
1!
1%
#73880000000
0!
0%
#73885000000
1!
1%
#73890000000
0!
0%
#73895000000
1!
1%
#73900000000
0!
0%
#73905000000
1!
1%
#73910000000
0!
0%
#73915000000
1!
1%
#73920000000
0!
0%
#73925000000
1!
1%
#73930000000
0!
0%
#73935000000
1!
1%
#73940000000
0!
0%
#73945000000
1!
1%
#73950000000
0!
0%
#73955000000
1!
1%
#73960000000
0!
0%
#73965000000
1!
1%
#73970000000
0!
0%
#73975000000
1!
1%
#73980000000
0!
0%
#73985000000
1!
1%
#73990000000
0!
0%
#73995000000
1!
1%
#74000000000
0!
0%
#74005000000
1!
1%
#74010000000
0!
0%
#74015000000
1!
1%
#74020000000
0!
0%
#74025000000
1!
1%
#74030000000
0!
0%
#74035000000
1!
1%
#74040000000
0!
0%
#74045000000
1!
1%
#74050000000
0!
0%
#74055000000
1!
1%
#74060000000
0!
0%
#74065000000
1!
1%
#74070000000
0!
0%
#74075000000
1!
1%
#74080000000
0!
0%
#74085000000
1!
1%
#74090000000
0!
0%
#74095000000
1!
1%
#74100000000
0!
0%
#74105000000
1!
1%
#74110000000
0!
0%
#74115000000
1!
1%
#74120000000
0!
0%
#74125000000
1!
1%
#74130000000
0!
0%
#74135000000
1!
1%
#74140000000
0!
0%
#74145000000
1!
1%
#74150000000
0!
0%
#74155000000
1!
1%
#74160000000
0!
0%
#74165000000
1!
1%
#74170000000
0!
0%
#74175000000
1!
1%
#74180000000
0!
0%
#74185000000
1!
1%
#74190000000
0!
0%
#74195000000
1!
1%
#74200000000
0!
0%
#74205000000
1!
1%
#74210000000
0!
0%
#74215000000
1!
1%
#74220000000
0!
0%
#74225000000
1!
1%
#74230000000
0!
0%
#74235000000
1!
1%
#74240000000
0!
0%
#74245000000
1!
1%
#74250000000
0!
0%
#74255000000
1!
1%
#74260000000
0!
0%
#74265000000
1!
1%
#74270000000
0!
0%
#74275000000
1!
1%
#74280000000
0!
0%
#74285000000
1!
1%
#74290000000
0!
0%
#74295000000
1!
1%
#74300000000
0!
0%
#74305000000
1!
1%
#74310000000
0!
0%
#74315000000
1!
1%
#74320000000
0!
0%
#74325000000
1!
1%
#74330000000
0!
0%
#74335000000
1!
1%
#74340000000
0!
0%
#74345000000
1!
1%
#74350000000
0!
0%
#74355000000
1!
1%
#74360000000
0!
0%
#74365000000
1!
1%
#74370000000
0!
0%
#74375000000
1!
1%
#74380000000
0!
0%
#74385000000
1!
1%
#74390000000
0!
0%
#74395000000
1!
1%
#74400000000
0!
0%
#74405000000
1!
1%
#74410000000
0!
0%
#74415000000
1!
1%
#74420000000
0!
0%
#74425000000
1!
1%
#74430000000
0!
0%
#74435000000
1!
1%
#74440000000
0!
0%
#74445000000
1!
1%
#74450000000
0!
0%
#74455000000
1!
1%
#74460000000
0!
0%
#74465000000
1!
1%
#74470000000
0!
0%
#74475000000
1!
1%
#74480000000
0!
0%
#74485000000
1!
1%
#74490000000
0!
0%
#74495000000
1!
1%
#74500000000
0!
0%
#74505000000
1!
1%
#74510000000
0!
0%
#74515000000
1!
1%
#74520000000
0!
0%
#74525000000
1!
1%
#74530000000
0!
0%
#74535000000
1!
1%
#74540000000
0!
0%
#74545000000
1!
1%
#74550000000
0!
0%
#74555000000
1!
1%
#74560000000
0!
0%
#74565000000
1!
1%
#74570000000
0!
0%
#74575000000
1!
1%
#74580000000
0!
0%
#74585000000
1!
1%
#74590000000
0!
0%
#74595000000
1!
1%
#74600000000
0!
0%
#74605000000
1!
1%
#74610000000
0!
0%
#74615000000
1!
1%
#74620000000
0!
0%
#74625000000
1!
1%
#74630000000
0!
0%
#74635000000
1!
1%
#74640000000
0!
0%
#74645000000
1!
1%
#74650000000
0!
0%
#74655000000
1!
1%
#74660000000
0!
0%
#74665000000
1!
1%
#74670000000
0!
0%
#74675000000
1!
1%
#74680000000
0!
0%
#74685000000
1!
1%
#74690000000
0!
0%
#74695000000
1!
1%
#74700000000
0!
0%
#74705000000
1!
1%
#74710000000
0!
0%
#74715000000
1!
1%
#74720000000
0!
0%
#74725000000
1!
1%
#74730000000
0!
0%
#74735000000
1!
1%
#74740000000
0!
0%
#74745000000
1!
1%
#74750000000
0!
0%
#74755000000
1!
1%
#74760000000
0!
0%
#74765000000
1!
1%
#74770000000
0!
0%
#74775000000
1!
1%
#74780000000
0!
0%
#74785000000
1!
1%
#74790000000
0!
0%
#74795000000
1!
1%
#74800000000
0!
0%
#74805000000
1!
1%
#74810000000
0!
0%
#74815000000
1!
1%
#74820000000
0!
0%
#74825000000
1!
1%
#74830000000
0!
0%
#74835000000
1!
1%
#74840000000
0!
0%
#74845000000
1!
1%
#74850000000
0!
0%
#74855000000
1!
1%
#74860000000
0!
0%
#74865000000
1!
1%
#74870000000
0!
0%
#74875000000
1!
1%
#74880000000
0!
0%
#74885000000
1!
1%
#74890000000
0!
0%
#74895000000
1!
1%
#74900000000
0!
0%
#74905000000
1!
1%
#74910000000
0!
0%
#74915000000
1!
1%
#74920000000
0!
0%
#74925000000
1!
1%
#74930000000
0!
0%
#74935000000
1!
1%
#74940000000
0!
0%
#74945000000
1!
1%
#74950000000
0!
0%
#74955000000
1!
1%
#74960000000
0!
0%
#74965000000
1!
1%
#74970000000
0!
0%
#74975000000
1!
1%
#74980000000
0!
0%
#74985000000
1!
1%
#74990000000
0!
0%
#74995000000
1!
1%
#75000000000
0!
0%
#75005000000
1!
1%
#75010000000
0!
0%
#75015000000
1!
1%
#75020000000
0!
0%
#75025000000
1!
1%
#75030000000
0!
0%
#75035000000
1!
1%
#75040000000
0!
0%
#75045000000
1!
1%
#75050000000
0!
0%
#75055000000
1!
1%
#75060000000
0!
0%
#75065000000
1!
1%
#75070000000
0!
0%
#75075000000
1!
1%
#75080000000
0!
0%
#75085000000
1!
1%
#75090000000
0!
0%
#75095000000
1!
1%
#75100000000
0!
0%
#75105000000
1!
1%
#75110000000
0!
0%
#75115000000
1!
1%
#75120000000
0!
0%
#75125000000
1!
1%
#75130000000
0!
0%
#75135000000
1!
1%
#75140000000
0!
0%
#75145000000
1!
1%
#75150000000
0!
0%
#75155000000
1!
1%
#75160000000
0!
0%
#75165000000
1!
1%
#75170000000
0!
0%
#75175000000
1!
1%
#75180000000
0!
0%
#75185000000
1!
1%
#75190000000
0!
0%
#75195000000
1!
1%
#75200000000
0!
0%
#75205000000
1!
1%
#75210000000
0!
0%
#75215000000
1!
1%
#75220000000
0!
0%
#75225000000
1!
1%
#75230000000
0!
0%
#75235000000
1!
1%
#75240000000
0!
0%
#75245000000
1!
1%
#75250000000
0!
0%
#75255000000
1!
1%
#75260000000
0!
0%
#75265000000
1!
1%
#75270000000
0!
0%
#75275000000
1!
1%
#75280000000
0!
0%
#75285000000
1!
1%
#75290000000
0!
0%
#75295000000
1!
1%
#75300000000
0!
0%
#75305000000
1!
1%
#75310000000
0!
0%
#75315000000
1!
1%
#75320000000
0!
0%
#75325000000
1!
1%
#75330000000
0!
0%
#75335000000
1!
1%
#75340000000
0!
0%
#75345000000
1!
1%
#75350000000
0!
0%
#75355000000
1!
1%
#75360000000
0!
0%
#75365000000
1!
1%
#75370000000
0!
0%
#75375000000
1!
1%
#75380000000
0!
0%
#75385000000
1!
1%
#75390000000
0!
0%
#75395000000
1!
1%
#75400000000
0!
0%
#75405000000
1!
1%
#75410000000
0!
0%
#75415000000
1!
1%
#75420000000
0!
0%
#75425000000
1!
1%
#75430000000
0!
0%
#75435000000
1!
1%
#75440000000
0!
0%
#75445000000
1!
1%
#75450000000
0!
0%
#75455000000
1!
1%
#75460000000
0!
0%
#75465000000
1!
1%
#75470000000
0!
0%
#75475000000
1!
1%
#75480000000
0!
0%
#75485000000
1!
1%
#75490000000
0!
0%
#75495000000
1!
1%
#75500000000
0!
0%
#75505000000
1!
1%
#75510000000
0!
0%
#75515000000
1!
1%
#75520000000
0!
0%
#75525000000
1!
1%
#75530000000
0!
0%
#75535000000
1!
1%
#75540000000
0!
0%
#75545000000
1!
1%
#75550000000
0!
0%
#75555000000
1!
1%
#75560000000
0!
0%
#75565000000
1!
1%
#75570000000
0!
0%
#75575000000
1!
1%
#75580000000
0!
0%
#75585000000
1!
1%
#75590000000
0!
0%
#75595000000
1!
1%
#75600000000
0!
0%
#75605000000
1!
1%
#75610000000
0!
0%
#75615000000
1!
1%
#75620000000
0!
0%
#75625000000
1!
1%
#75630000000
0!
0%
#75635000000
1!
1%
#75640000000
0!
0%
#75645000000
1!
1%
#75650000000
0!
0%
#75655000000
1!
1%
#75660000000
0!
0%
#75665000000
1!
1%
#75670000000
0!
0%
#75675000000
1!
1%
#75680000000
0!
0%
#75685000000
1!
1%
#75690000000
0!
0%
#75695000000
1!
1%
#75700000000
0!
0%
#75705000000
1!
1%
#75710000000
0!
0%
#75715000000
1!
1%
#75720000000
0!
0%
#75725000000
1!
1%
#75730000000
0!
0%
#75735000000
1!
1%
#75740000000
0!
0%
#75745000000
1!
1%
#75750000000
0!
0%
#75755000000
1!
1%
#75760000000
0!
0%
#75765000000
1!
1%
#75770000000
0!
0%
#75775000000
1!
1%
#75780000000
0!
0%
#75785000000
1!
1%
#75790000000
0!
0%
#75795000000
1!
1%
#75800000000
0!
0%
#75805000000
1!
1%
#75810000000
0!
0%
#75815000000
1!
1%
#75820000000
0!
0%
#75825000000
1!
1%
#75830000000
0!
0%
#75835000000
1!
1%
#75840000000
0!
0%
#75845000000
1!
1%
#75850000000
0!
0%
#75855000000
1!
1%
#75860000000
0!
0%
#75865000000
1!
1%
#75870000000
0!
0%
#75875000000
1!
1%
#75880000000
0!
0%
#75885000000
1!
1%
#75890000000
0!
0%
#75895000000
1!
1%
#75900000000
0!
0%
#75905000000
1!
1%
#75910000000
0!
0%
#75915000000
1!
1%
#75920000000
0!
0%
#75925000000
1!
1%
#75930000000
0!
0%
#75935000000
1!
1%
#75940000000
0!
0%
#75945000000
1!
1%
#75950000000
0!
0%
#75955000000
1!
1%
#75960000000
0!
0%
#75965000000
1!
1%
#75970000000
0!
0%
#75975000000
1!
1%
#75980000000
0!
0%
#75985000000
1!
1%
#75990000000
0!
0%
#75995000000
1!
1%
#76000000000
0!
0%
#76005000000
1!
1%
#76010000000
0!
0%
#76015000000
1!
1%
#76020000000
0!
0%
#76025000000
1!
1%
#76030000000
0!
0%
#76035000000
1!
1%
#76040000000
0!
0%
#76045000000
1!
1%
#76050000000
0!
0%
#76055000000
1!
1%
#76060000000
0!
0%
#76065000000
1!
1%
#76070000000
0!
0%
#76075000000
1!
1%
#76080000000
0!
0%
#76085000000
1!
1%
#76090000000
0!
0%
#76095000000
1!
1%
#76100000000
0!
0%
#76105000000
1!
1%
#76110000000
0!
0%
#76115000000
1!
1%
#76120000000
0!
0%
#76125000000
1!
1%
#76130000000
0!
0%
#76135000000
1!
1%
#76140000000
0!
0%
#76145000000
1!
1%
#76150000000
0!
0%
#76155000000
1!
1%
#76160000000
0!
0%
#76165000000
1!
1%
#76170000000
0!
0%
#76175000000
1!
1%
#76180000000
0!
0%
#76185000000
1!
1%
#76190000000
0!
0%
#76195000000
1!
1%
#76200000000
0!
0%
#76205000000
1!
1%
#76210000000
0!
0%
#76215000000
1!
1%
#76220000000
0!
0%
#76225000000
1!
1%
#76230000000
0!
0%
#76235000000
1!
1%
#76240000000
0!
0%
#76245000000
1!
1%
#76250000000
0!
0%
#76255000000
1!
1%
#76260000000
0!
0%
#76265000000
1!
1%
#76270000000
0!
0%
#76275000000
1!
1%
#76280000000
0!
0%
#76285000000
1!
1%
#76290000000
0!
0%
#76295000000
1!
1%
#76300000000
0!
0%
#76305000000
1!
1%
#76310000000
0!
0%
#76315000000
1!
1%
#76320000000
0!
0%
#76325000000
1!
1%
#76330000000
0!
0%
#76335000000
1!
1%
#76340000000
0!
0%
#76345000000
1!
1%
#76350000000
0!
0%
#76355000000
1!
1%
#76360000000
0!
0%
#76365000000
1!
1%
#76370000000
0!
0%
#76375000000
1!
1%
#76380000000
0!
0%
#76385000000
1!
1%
#76390000000
0!
0%
#76395000000
1!
1%
#76400000000
0!
0%
#76405000000
1!
1%
#76410000000
0!
0%
#76415000000
1!
1%
#76420000000
0!
0%
#76425000000
1!
1%
#76430000000
0!
0%
#76435000000
1!
1%
#76440000000
0!
0%
#76445000000
1!
1%
#76450000000
0!
0%
#76455000000
1!
1%
#76460000000
0!
0%
#76465000000
1!
1%
#76470000000
0!
0%
#76475000000
1!
1%
#76480000000
0!
0%
#76485000000
1!
1%
#76490000000
0!
0%
#76495000000
1!
1%
#76500000000
0!
0%
#76505000000
1!
1%
#76510000000
0!
0%
#76515000000
1!
1%
#76520000000
0!
0%
#76525000000
1!
1%
#76530000000
0!
0%
#76535000000
1!
1%
#76540000000
0!
0%
#76545000000
1!
1%
#76550000000
0!
0%
#76555000000
1!
1%
#76560000000
0!
0%
#76565000000
1!
1%
#76570000000
0!
0%
#76575000000
1!
1%
#76580000000
0!
0%
#76585000000
1!
1%
#76590000000
0!
0%
#76595000000
1!
1%
#76600000000
0!
0%
#76605000000
1!
1%
#76610000000
0!
0%
#76615000000
1!
1%
#76620000000
0!
0%
#76625000000
1!
1%
#76630000000
0!
0%
#76635000000
1!
1%
#76640000000
0!
0%
#76645000000
1!
1%
#76650000000
0!
0%
#76655000000
1!
1%
#76660000000
0!
0%
#76665000000
1!
1%
#76670000000
0!
0%
#76675000000
1!
1%
#76680000000
0!
0%
#76685000000
1!
1%
#76690000000
0!
0%
#76695000000
1!
1%
#76700000000
0!
0%
#76705000000
1!
1%
#76710000000
0!
0%
#76715000000
1!
1%
#76720000000
0!
0%
#76725000000
1!
1%
#76730000000
0!
0%
#76735000000
1!
1%
#76740000000
0!
0%
#76745000000
1!
1%
#76750000000
0!
0%
#76755000000
1!
1%
#76760000000
0!
0%
#76765000000
1!
1%
#76770000000
0!
0%
#76775000000
1!
1%
#76780000000
0!
0%
#76785000000
1!
1%
#76790000000
0!
0%
#76795000000
1!
1%
#76800000000
0!
0%
#76805000000
1!
1%
#76810000000
0!
0%
#76815000000
1!
1%
#76820000000
0!
0%
#76825000000
1!
1%
#76830000000
0!
0%
#76835000000
1!
1%
#76840000000
0!
0%
#76845000000
1!
1%
#76850000000
0!
0%
#76855000000
1!
1%
#76860000000
0!
0%
#76865000000
1!
1%
#76870000000
0!
0%
#76875000000
1!
1%
#76880000000
0!
0%
#76885000000
1!
1%
#76890000000
0!
0%
#76895000000
1!
1%
#76900000000
0!
0%
#76905000000
1!
1%
#76910000000
0!
0%
#76915000000
1!
1%
#76920000000
0!
0%
#76925000000
1!
1%
#76930000000
0!
0%
#76935000000
1!
1%
#76940000000
0!
0%
#76945000000
1!
1%
#76950000000
0!
0%
#76955000000
1!
1%
#76960000000
0!
0%
#76965000000
1!
1%
#76970000000
0!
0%
#76975000000
1!
1%
#76980000000
0!
0%
#76985000000
1!
1%
#76990000000
0!
0%
#76995000000
1!
1%
#77000000000
0!
0%
#77005000000
1!
1%
#77010000000
0!
0%
#77015000000
1!
1%
#77020000000
0!
0%
#77025000000
1!
1%
#77030000000
0!
0%
#77035000000
1!
1%
#77040000000
0!
0%
#77045000000
1!
1%
#77050000000
0!
0%
#77055000000
1!
1%
#77060000000
0!
0%
#77065000000
1!
1%
#77070000000
0!
0%
#77075000000
1!
1%
#77080000000
0!
0%
#77085000000
1!
1%
#77090000000
0!
0%
#77095000000
1!
1%
#77100000000
0!
0%
#77105000000
1!
1%
#77110000000
0!
0%
#77115000000
1!
1%
#77120000000
0!
0%
#77125000000
1!
1%
#77130000000
0!
0%
#77135000000
1!
1%
#77140000000
0!
0%
#77145000000
1!
1%
#77150000000
0!
0%
#77155000000
1!
1%
#77160000000
0!
0%
#77165000000
1!
1%
#77170000000
0!
0%
#77175000000
1!
1%
#77180000000
0!
0%
#77185000000
1!
1%
#77190000000
0!
0%
#77195000000
1!
1%
#77200000000
0!
0%
#77205000000
1!
1%
#77210000000
0!
0%
#77215000000
1!
1%
#77220000000
0!
0%
#77225000000
1!
1%
#77230000000
0!
0%
#77235000000
1!
1%
#77240000000
0!
0%
#77245000000
1!
1%
#77250000000
0!
0%
#77255000000
1!
1%
#77260000000
0!
0%
#77265000000
1!
1%
#77270000000
0!
0%
#77275000000
1!
1%
#77280000000
0!
0%
#77285000000
1!
1%
#77290000000
0!
0%
#77295000000
1!
1%
#77300000000
0!
0%
#77305000000
1!
1%
#77310000000
0!
0%
#77315000000
1!
1%
#77320000000
0!
0%
#77325000000
1!
1%
#77330000000
0!
0%
#77335000000
1!
1%
#77340000000
0!
0%
#77345000000
1!
1%
#77350000000
0!
0%
#77355000000
1!
1%
#77360000000
0!
0%
#77365000000
1!
1%
#77370000000
0!
0%
#77375000000
1!
1%
#77380000000
0!
0%
#77385000000
1!
1%
#77390000000
0!
0%
#77395000000
1!
1%
#77400000000
0!
0%
#77405000000
1!
1%
#77410000000
0!
0%
#77415000000
1!
1%
#77420000000
0!
0%
#77425000000
1!
1%
#77430000000
0!
0%
#77435000000
1!
1%
#77440000000
0!
0%
#77445000000
1!
1%
#77450000000
0!
0%
#77455000000
1!
1%
#77460000000
0!
0%
#77465000000
1!
1%
#77470000000
0!
0%
#77475000000
1!
1%
#77480000000
0!
0%
#77485000000
1!
1%
#77490000000
0!
0%
#77495000000
1!
1%
#77500000000
0!
0%
#77505000000
1!
1%
#77510000000
0!
0%
#77515000000
1!
1%
#77520000000
0!
0%
#77525000000
1!
1%
#77530000000
0!
0%
#77535000000
1!
1%
#77540000000
0!
0%
#77545000000
1!
1%
#77550000000
0!
0%
#77555000000
1!
1%
#77560000000
0!
0%
#77565000000
1!
1%
#77570000000
0!
0%
#77575000000
1!
1%
#77580000000
0!
0%
#77585000000
1!
1%
#77590000000
0!
0%
#77595000000
1!
1%
#77600000000
0!
0%
#77605000000
1!
1%
#77610000000
0!
0%
#77615000000
1!
1%
#77620000000
0!
0%
#77625000000
1!
1%
#77630000000
0!
0%
#77635000000
1!
1%
#77640000000
0!
0%
#77645000000
1!
1%
#77650000000
0!
0%
#77655000000
1!
1%
#77660000000
0!
0%
#77665000000
1!
1%
#77670000000
0!
0%
#77675000000
1!
1%
#77680000000
0!
0%
#77685000000
1!
1%
#77690000000
0!
0%
#77695000000
1!
1%
#77700000000
0!
0%
#77705000000
1!
1%
#77710000000
0!
0%
#77715000000
1!
1%
#77720000000
0!
0%
#77725000000
1!
1%
#77730000000
0!
0%
#77735000000
1!
1%
#77740000000
0!
0%
#77745000000
1!
1%
#77750000000
0!
0%
#77755000000
1!
1%
#77760000000
0!
0%
#77765000000
1!
1%
#77770000000
0!
0%
#77775000000
1!
1%
#77780000000
0!
0%
#77785000000
1!
1%
#77790000000
0!
0%
#77795000000
1!
1%
#77800000000
0!
0%
#77805000000
1!
1%
#77810000000
0!
0%
#77815000000
1!
1%
#77820000000
0!
0%
#77825000000
1!
1%
#77830000000
0!
0%
#77835000000
1!
1%
#77840000000
0!
0%
#77845000000
1!
1%
#77850000000
0!
0%
#77855000000
1!
1%
#77860000000
0!
0%
#77865000000
1!
1%
#77870000000
0!
0%
#77875000000
1!
1%
#77880000000
0!
0%
#77885000000
1!
1%
#77890000000
0!
0%
#77895000000
1!
1%
#77900000000
0!
0%
#77905000000
1!
1%
#77910000000
0!
0%
#77915000000
1!
1%
#77920000000
0!
0%
#77925000000
1!
1%
#77930000000
0!
0%
#77935000000
1!
1%
#77940000000
0!
0%
#77945000000
1!
1%
#77950000000
0!
0%
#77955000000
1!
1%
#77960000000
0!
0%
#77965000000
1!
1%
#77970000000
0!
0%
#77975000000
1!
1%
#77980000000
0!
0%
#77985000000
1!
1%
#77990000000
0!
0%
#77995000000
1!
1%
#78000000000
0!
0%
#78005000000
1!
1%
#78010000000
0!
0%
#78015000000
1!
1%
#78020000000
0!
0%
#78025000000
1!
1%
#78030000000
0!
0%
#78035000000
1!
1%
#78040000000
0!
0%
#78045000000
1!
1%
#78050000000
0!
0%
#78055000000
1!
1%
#78060000000
0!
0%
#78065000000
1!
1%
#78070000000
0!
0%
#78075000000
1!
1%
#78080000000
0!
0%
#78085000000
1!
1%
#78090000000
0!
0%
#78095000000
1!
1%
#78100000000
0!
0%
#78105000000
1!
1%
#78110000000
0!
0%
#78115000000
1!
1%
#78120000000
0!
0%
#78125000000
1!
1%
#78130000000
0!
0%
#78135000000
1!
1%
#78140000000
0!
0%
#78145000000
1!
1%
#78150000000
0!
0%
#78155000000
1!
1%
#78160000000
0!
0%
#78165000000
1!
1%
#78170000000
0!
0%
#78175000000
1!
1%
#78180000000
0!
0%
#78185000000
1!
1%
#78190000000
0!
0%
#78195000000
1!
1%
#78200000000
0!
0%
#78205000000
1!
1%
#78210000000
0!
0%
#78215000000
1!
1%
#78220000000
0!
0%
#78225000000
1!
1%
#78230000000
0!
0%
#78235000000
1!
1%
#78240000000
0!
0%
#78245000000
1!
1%
#78250000000
0!
0%
#78255000000
1!
1%
#78260000000
0!
0%
#78265000000
1!
1%
#78270000000
0!
0%
#78275000000
1!
1%
#78280000000
0!
0%
#78285000000
1!
1%
#78290000000
0!
0%
#78295000000
1!
1%
#78300000000
0!
0%
#78305000000
1!
1%
#78310000000
0!
0%
#78315000000
1!
1%
#78320000000
0!
0%
#78325000000
1!
1%
#78330000000
0!
0%
#78335000000
1!
1%
#78340000000
0!
0%
#78345000000
1!
1%
#78350000000
0!
0%
#78355000000
1!
1%
#78360000000
0!
0%
#78365000000
1!
1%
#78370000000
0!
0%
#78375000000
1!
1%
#78380000000
0!
0%
#78385000000
1!
1%
#78390000000
0!
0%
#78395000000
1!
1%
#78400000000
0!
0%
#78405000000
1!
1%
#78410000000
0!
0%
#78415000000
1!
1%
#78420000000
0!
0%
#78425000000
1!
1%
#78430000000
0!
0%
#78435000000
1!
1%
#78440000000
0!
0%
#78445000000
1!
1%
#78450000000
0!
0%
#78455000000
1!
1%
#78460000000
0!
0%
#78465000000
1!
1%
#78470000000
0!
0%
#78475000000
1!
1%
#78480000000
0!
0%
#78485000000
1!
1%
#78490000000
0!
0%
#78495000000
1!
1%
#78500000000
0!
0%
#78505000000
1!
1%
#78510000000
0!
0%
#78515000000
1!
1%
#78520000000
0!
0%
#78525000000
1!
1%
#78530000000
0!
0%
#78535000000
1!
1%
#78540000000
0!
0%
#78545000000
1!
1%
#78550000000
0!
0%
#78555000000
1!
1%
#78560000000
0!
0%
#78565000000
1!
1%
#78570000000
0!
0%
#78575000000
1!
1%
#78580000000
0!
0%
#78585000000
1!
1%
#78590000000
0!
0%
#78595000000
1!
1%
#78600000000
0!
0%
#78605000000
1!
1%
#78610000000
0!
0%
#78615000000
1!
1%
#78620000000
0!
0%
#78625000000
1!
1%
#78630000000
0!
0%
#78635000000
1!
1%
#78640000000
0!
0%
#78645000000
1!
1%
#78650000000
0!
0%
#78655000000
1!
1%
#78660000000
0!
0%
#78665000000
1!
1%
#78670000000
0!
0%
#78675000000
1!
1%
#78680000000
0!
0%
#78685000000
1!
1%
#78690000000
0!
0%
#78695000000
1!
1%
#78700000000
0!
0%
#78705000000
1!
1%
#78710000000
0!
0%
#78715000000
1!
1%
#78720000000
0!
0%
#78725000000
1!
1%
#78730000000
0!
0%
#78735000000
1!
1%
#78740000000
0!
0%
#78745000000
1!
1%
#78750000000
0!
0%
#78755000000
1!
1%
#78760000000
0!
0%
#78765000000
1!
1%
#78770000000
0!
0%
#78775000000
1!
1%
#78780000000
0!
0%
#78785000000
1!
1%
#78790000000
0!
0%
#78795000000
1!
1%
#78800000000
0!
0%
#78805000000
1!
1%
#78810000000
0!
0%
#78815000000
1!
1%
#78820000000
0!
0%
#78825000000
1!
1%
#78830000000
0!
0%
#78835000000
1!
1%
#78840000000
0!
0%
#78845000000
1!
1%
#78850000000
0!
0%
#78855000000
1!
1%
#78860000000
0!
0%
#78865000000
1!
1%
#78870000000
0!
0%
#78875000000
1!
1%
#78880000000
0!
0%
#78885000000
1!
1%
#78890000000
0!
0%
#78895000000
1!
1%
#78900000000
0!
0%
#78905000000
1!
1%
#78910000000
0!
0%
#78915000000
1!
1%
#78920000000
0!
0%
#78925000000
1!
1%
#78930000000
0!
0%
#78935000000
1!
1%
#78940000000
0!
0%
#78945000000
1!
1%
#78950000000
0!
0%
#78955000000
1!
1%
#78960000000
0!
0%
#78965000000
1!
1%
#78970000000
0!
0%
#78975000000
1!
1%
#78980000000
0!
0%
#78985000000
1!
1%
#78990000000
0!
0%
#78995000000
1!
1%
#79000000000
0!
0%
#79005000000
1!
1%
#79010000000
0!
0%
#79015000000
1!
1%
#79020000000
0!
0%
#79025000000
1!
1%
#79030000000
0!
0%
#79035000000
1!
1%
#79040000000
0!
0%
#79045000000
1!
1%
#79050000000
0!
0%
#79055000000
1!
1%
#79060000000
0!
0%
#79065000000
1!
1%
#79070000000
0!
0%
#79075000000
1!
1%
#79080000000
0!
0%
#79085000000
1!
1%
#79090000000
0!
0%
#79095000000
1!
1%
#79100000000
0!
0%
#79105000000
1!
1%
#79110000000
0!
0%
#79115000000
1!
1%
#79120000000
0!
0%
#79125000000
1!
1%
#79130000000
0!
0%
#79135000000
1!
1%
#79140000000
0!
0%
#79145000000
1!
1%
#79150000000
0!
0%
#79155000000
1!
1%
#79160000000
0!
0%
#79165000000
1!
1%
#79170000000
0!
0%
#79175000000
1!
1%
#79180000000
0!
0%
#79185000000
1!
1%
#79190000000
0!
0%
#79195000000
1!
1%
#79200000000
0!
0%
#79205000000
1!
1%
#79210000000
0!
0%
#79215000000
1!
1%
#79220000000
0!
0%
#79225000000
1!
1%
#79230000000
0!
0%
#79235000000
1!
1%
#79240000000
0!
0%
#79245000000
1!
1%
#79250000000
0!
0%
#79255000000
1!
1%
#79260000000
0!
0%
#79265000000
1!
1%
#79270000000
0!
0%
#79275000000
1!
1%
#79280000000
0!
0%
#79285000000
1!
1%
#79290000000
0!
0%
#79295000000
1!
1%
#79300000000
0!
0%
#79305000000
1!
1%
#79310000000
0!
0%
#79315000000
1!
1%
#79320000000
0!
0%
#79325000000
1!
1%
#79330000000
0!
0%
#79335000000
1!
1%
#79340000000
0!
0%
#79345000000
1!
1%
#79350000000
0!
0%
#79355000000
1!
1%
#79360000000
0!
0%
#79365000000
1!
1%
#79370000000
0!
0%
#79375000000
1!
1%
#79380000000
0!
0%
#79385000000
1!
1%
#79390000000
0!
0%
#79395000000
1!
1%
#79400000000
0!
0%
#79405000000
1!
1%
#79410000000
0!
0%
#79415000000
1!
1%
#79420000000
0!
0%
#79425000000
1!
1%
#79430000000
0!
0%
#79435000000
1!
1%
#79440000000
0!
0%
#79445000000
1!
1%
#79450000000
0!
0%
#79455000000
1!
1%
#79460000000
0!
0%
#79465000000
1!
1%
#79470000000
0!
0%
#79475000000
1!
1%
#79480000000
0!
0%
#79485000000
1!
1%
#79490000000
0!
0%
#79495000000
1!
1%
#79500000000
0!
0%
#79505000000
1!
1%
#79510000000
0!
0%
#79515000000
1!
1%
#79520000000
0!
0%
#79525000000
1!
1%
#79530000000
0!
0%
#79535000000
1!
1%
#79540000000
0!
0%
#79545000000
1!
1%
#79550000000
0!
0%
#79555000000
1!
1%
#79560000000
0!
0%
#79565000000
1!
1%
#79570000000
0!
0%
#79575000000
1!
1%
#79580000000
0!
0%
#79585000000
1!
1%
#79590000000
0!
0%
#79595000000
1!
1%
#79600000000
0!
0%
#79605000000
1!
1%
#79610000000
0!
0%
#79615000000
1!
1%
#79620000000
0!
0%
#79625000000
1!
1%
#79630000000
0!
0%
#79635000000
1!
1%
#79640000000
0!
0%
#79645000000
1!
1%
#79650000000
0!
0%
#79655000000
1!
1%
#79660000000
0!
0%
#79665000000
1!
1%
#79670000000
0!
0%
#79675000000
1!
1%
#79680000000
0!
0%
#79685000000
1!
1%
#79690000000
0!
0%
#79695000000
1!
1%
#79700000000
0!
0%
#79705000000
1!
1%
#79710000000
0!
0%
#79715000000
1!
1%
#79720000000
0!
0%
#79725000000
1!
1%
#79730000000
0!
0%
#79735000000
1!
1%
#79740000000
0!
0%
#79745000000
1!
1%
#79750000000
0!
0%
#79755000000
1!
1%
#79760000000
0!
0%
#79765000000
1!
1%
#79770000000
0!
0%
#79775000000
1!
1%
#79780000000
0!
0%
#79785000000
1!
1%
#79790000000
0!
0%
#79795000000
1!
1%
#79800000000
0!
0%
#79805000000
1!
1%
#79810000000
0!
0%
#79815000000
1!
1%
#79820000000
0!
0%
#79825000000
1!
1%
#79830000000
0!
0%
#79835000000
1!
1%
#79840000000
0!
0%
#79845000000
1!
1%
#79850000000
0!
0%
#79855000000
1!
1%
#79860000000
0!
0%
#79865000000
1!
1%
#79870000000
0!
0%
#79875000000
1!
1%
#79880000000
0!
0%
#79885000000
1!
1%
#79890000000
0!
0%
#79895000000
1!
1%
#79900000000
0!
0%
#79905000000
1!
1%
#79910000000
0!
0%
#79915000000
1!
1%
#79920000000
0!
0%
#79925000000
1!
1%
#79930000000
0!
0%
#79935000000
1!
1%
#79940000000
0!
0%
#79945000000
1!
1%
#79950000000
0!
0%
#79955000000
1!
1%
#79960000000
0!
0%
#79965000000
1!
1%
#79970000000
0!
0%
#79975000000
1!
1%
#79980000000
0!
0%
#79985000000
1!
1%
#79990000000
0!
0%
#79995000000
1!
1%
#80000000000
0!
0%
#80005000000
1!
1%
#80010000000
0!
0%
#80015000000
1!
1%
#80020000000
0!
0%
#80025000000
1!
1%
#80030000000
0!
0%
#80035000000
1!
1%
#80040000000
0!
0%
#80045000000
1!
1%
#80050000000
0!
0%
#80055000000
1!
1%
#80060000000
0!
0%
#80065000000
1!
1%
#80070000000
0!
0%
#80075000000
1!
1%
#80080000000
0!
0%
#80085000000
1!
1%
#80090000000
0!
0%
#80095000000
1!
1%
#80100000000
0!
0%
#80105000000
1!
1%
#80110000000
0!
0%
#80115000000
1!
1%
#80120000000
0!
0%
#80125000000
1!
1%
#80130000000
0!
0%
#80135000000
1!
1%
#80140000000
0!
0%
#80145000000
1!
1%
#80150000000
0!
0%
#80155000000
1!
1%
#80160000000
0!
0%
#80165000000
1!
1%
#80170000000
0!
0%
#80175000000
1!
1%
#80180000000
0!
0%
#80185000000
1!
1%
#80190000000
0!
0%
#80195000000
1!
1%
#80200000000
0!
0%
#80205000000
1!
1%
#80210000000
0!
0%
#80215000000
1!
1%
#80220000000
0!
0%
#80225000000
1!
1%
#80230000000
0!
0%
#80235000000
1!
1%
#80240000000
0!
0%
#80245000000
1!
1%
#80250000000
0!
0%
#80255000000
1!
1%
#80260000000
0!
0%
#80265000000
1!
1%
#80270000000
0!
0%
#80275000000
1!
1%
#80280000000
0!
0%
#80285000000
1!
1%
#80290000000
0!
0%
#80295000000
1!
1%
#80300000000
0!
0%
#80305000000
1!
1%
#80310000000
0!
0%
#80315000000
1!
1%
#80320000000
0!
0%
#80325000000
1!
1%
#80330000000
0!
0%
#80335000000
1!
1%
#80340000000
0!
0%
#80345000000
1!
1%
#80350000000
0!
0%
#80355000000
1!
1%
#80360000000
0!
0%
#80365000000
1!
1%
#80370000000
0!
0%
#80375000000
1!
1%
#80380000000
0!
0%
#80385000000
1!
1%
#80390000000
0!
0%
#80395000000
1!
1%
#80400000000
0!
0%
#80405000000
1!
1%
#80410000000
0!
0%
#80415000000
1!
1%
#80420000000
0!
0%
#80425000000
1!
1%
#80430000000
0!
0%
#80435000000
1!
1%
#80440000000
0!
0%
#80445000000
1!
1%
#80450000000
0!
0%
#80455000000
1!
1%
#80460000000
0!
0%
#80465000000
1!
1%
#80470000000
0!
0%
#80475000000
1!
1%
#80480000000
0!
0%
#80485000000
1!
1%
#80490000000
0!
0%
#80495000000
1!
1%
#80500000000
0!
0%
#80505000000
1!
1%
#80510000000
0!
0%
#80515000000
1!
1%
#80520000000
0!
0%
#80525000000
1!
1%
#80530000000
0!
0%
#80535000000
1!
1%
#80540000000
0!
0%
#80545000000
1!
1%
#80550000000
0!
0%
#80555000000
1!
1%
#80560000000
0!
0%
#80565000000
1!
1%
#80570000000
0!
0%
#80575000000
1!
1%
#80580000000
0!
0%
#80585000000
1!
1%
#80590000000
0!
0%
#80595000000
1!
1%
#80600000000
0!
0%
#80605000000
1!
1%
#80610000000
0!
0%
#80615000000
1!
1%
#80620000000
0!
0%
#80625000000
1!
1%
#80630000000
0!
0%
#80635000000
1!
1%
#80640000000
0!
0%
#80645000000
1!
1%
#80650000000
0!
0%
#80655000000
1!
1%
#80660000000
0!
0%
#80665000000
1!
1%
#80670000000
0!
0%
#80675000000
1!
1%
#80680000000
0!
0%
#80685000000
1!
1%
#80690000000
0!
0%
#80695000000
1!
1%
#80700000000
0!
0%
#80705000000
1!
1%
#80710000000
0!
0%
#80715000000
1!
1%
#80720000000
0!
0%
#80725000000
1!
1%
#80730000000
0!
0%
#80735000000
1!
1%
#80740000000
0!
0%
#80745000000
1!
1%
#80750000000
0!
0%
#80755000000
1!
1%
#80760000000
0!
0%
#80765000000
1!
1%
#80770000000
0!
0%
#80775000000
1!
1%
#80780000000
0!
0%
#80785000000
1!
1%
#80790000000
0!
0%
#80795000000
1!
1%
#80800000000
0!
0%
#80805000000
1!
1%
#80810000000
0!
0%
#80815000000
1!
1%
#80820000000
0!
0%
#80825000000
1!
1%
#80830000000
0!
0%
#80835000000
1!
1%
#80840000000
0!
0%
#80845000000
1!
1%
#80850000000
0!
0%
#80855000000
1!
1%
#80860000000
0!
0%
#80865000000
1!
1%
#80870000000
0!
0%
#80875000000
1!
1%
#80880000000
0!
0%
#80885000000
1!
1%
#80890000000
0!
0%
#80895000000
1!
1%
#80900000000
0!
0%
#80905000000
1!
1%
#80910000000
0!
0%
#80915000000
1!
1%
#80920000000
0!
0%
#80925000000
1!
1%
#80930000000
0!
0%
#80935000000
1!
1%
#80940000000
0!
0%
#80945000000
1!
1%
#80950000000
0!
0%
#80955000000
1!
1%
#80960000000
0!
0%
#80965000000
1!
1%
#80970000000
0!
0%
#80975000000
1!
1%
#80980000000
0!
0%
#80985000000
1!
1%
#80990000000
0!
0%
#80995000000
1!
1%
#81000000000
0!
0%
#81005000000
1!
1%
#81010000000
0!
0%
#81015000000
1!
1%
#81020000000
0!
0%
#81025000000
1!
1%
#81030000000
0!
0%
#81035000000
1!
1%
#81040000000
0!
0%
#81045000000
1!
1%
#81050000000
0!
0%
#81055000000
1!
1%
#81060000000
0!
0%
#81065000000
1!
1%
#81070000000
0!
0%
#81075000000
1!
1%
#81080000000
0!
0%
#81085000000
1!
1%
#81090000000
0!
0%
#81095000000
1!
1%
#81100000000
0!
0%
#81105000000
1!
1%
#81110000000
0!
0%
#81115000000
1!
1%
#81120000000
0!
0%
#81125000000
1!
1%
#81130000000
0!
0%
#81135000000
1!
1%
#81140000000
0!
0%
#81145000000
1!
1%
#81150000000
0!
0%
#81155000000
1!
1%
#81160000000
0!
0%
#81165000000
1!
1%
#81170000000
0!
0%
#81175000000
1!
1%
#81180000000
0!
0%
#81185000000
1!
1%
#81190000000
0!
0%
#81195000000
1!
1%
#81200000000
0!
0%
#81205000000
1!
1%
#81210000000
0!
0%
#81215000000
1!
1%
#81220000000
0!
0%
#81225000000
1!
1%
#81230000000
0!
0%
#81235000000
1!
1%
#81240000000
0!
0%
#81245000000
1!
1%
#81250000000
0!
0%
#81255000000
1!
1%
#81260000000
0!
0%
#81265000000
1!
1%
#81270000000
0!
0%
#81275000000
1!
1%
#81280000000
0!
0%
#81285000000
1!
1%
#81290000000
0!
0%
#81295000000
1!
1%
#81300000000
0!
0%
#81305000000
1!
1%
#81310000000
0!
0%
#81315000000
1!
1%
#81320000000
0!
0%
#81325000000
1!
1%
#81330000000
0!
0%
#81335000000
1!
1%
#81340000000
0!
0%
#81345000000
1!
1%
#81350000000
0!
0%
#81355000000
1!
1%
#81360000000
0!
0%
#81365000000
1!
1%
#81370000000
0!
0%
#81375000000
1!
1%
#81380000000
0!
0%
#81385000000
1!
1%
#81390000000
0!
0%
#81395000000
1!
1%
#81400000000
0!
0%
#81405000000
1!
1%
#81410000000
0!
0%
#81415000000
1!
1%
#81420000000
0!
0%
#81425000000
1!
1%
#81430000000
0!
0%
#81435000000
1!
1%
#81440000000
0!
0%
#81445000000
1!
1%
#81450000000
0!
0%
#81455000000
1!
1%
#81460000000
0!
0%
#81465000000
1!
1%
#81470000000
0!
0%
#81475000000
1!
1%
#81480000000
0!
0%
#81485000000
1!
1%
#81490000000
0!
0%
#81495000000
1!
1%
#81500000000
0!
0%
#81505000000
1!
1%
#81510000000
0!
0%
#81515000000
1!
1%
#81520000000
0!
0%
#81525000000
1!
1%
#81530000000
0!
0%
#81535000000
1!
1%
#81540000000
0!
0%
#81545000000
1!
1%
#81550000000
0!
0%
#81555000000
1!
1%
#81560000000
0!
0%
#81565000000
1!
1%
#81570000000
0!
0%
#81575000000
1!
1%
#81580000000
0!
0%
#81585000000
1!
1%
#81590000000
0!
0%
#81595000000
1!
1%
#81600000000
0!
0%
#81605000000
1!
1%
#81610000000
0!
0%
#81615000000
1!
1%
#81620000000
0!
0%
#81625000000
1!
1%
#81630000000
0!
0%
#81635000000
1!
1%
#81640000000
0!
0%
#81645000000
1!
1%
#81650000000
0!
0%
#81655000000
1!
1%
#81660000000
0!
0%
#81665000000
1!
1%
#81670000000
0!
0%
#81675000000
1!
1%
#81680000000
0!
0%
#81685000000
1!
1%
#81690000000
0!
0%
#81695000000
1!
1%
#81700000000
0!
0%
#81705000000
1!
1%
#81710000000
0!
0%
#81715000000
1!
1%
#81720000000
0!
0%
#81725000000
1!
1%
#81730000000
0!
0%
#81735000000
1!
1%
#81740000000
0!
0%
#81745000000
1!
1%
#81750000000
0!
0%
#81755000000
1!
1%
#81760000000
0!
0%
#81765000000
1!
1%
#81770000000
0!
0%
#81775000000
1!
1%
#81780000000
0!
0%
#81785000000
1!
1%
#81790000000
0!
0%
#81795000000
1!
1%
#81800000000
0!
0%
#81805000000
1!
1%
#81810000000
0!
0%
#81815000000
1!
1%
#81820000000
0!
0%
#81825000000
1!
1%
#81830000000
0!
0%
#81835000000
1!
1%
#81840000000
0!
0%
#81845000000
1!
1%
#81850000000
0!
0%
#81855000000
1!
1%
#81860000000
0!
0%
#81865000000
1!
1%
#81870000000
0!
0%
#81875000000
1!
1%
#81880000000
0!
0%
#81885000000
1!
1%
#81890000000
0!
0%
#81895000000
1!
1%
#81900000000
0!
0%
#81905000000
1!
1%
#81910000000
0!
0%
#81915000000
1!
1%
#81920000000
0!
0%
#81925000000
1!
1%
#81930000000
0!
0%
#81935000000
1!
1%
#81940000000
0!
0%
#81945000000
1!
1%
#81950000000
0!
0%
#81955000000
1!
1%
#81960000000
0!
0%
#81965000000
1!
1%
#81970000000
0!
0%
#81975000000
1!
1%
#81980000000
0!
0%
#81985000000
1!
1%
#81990000000
0!
0%
#81995000000
1!
1%
#82000000000
0!
0%
#82005000000
1!
1%
#82010000000
0!
0%
#82015000000
1!
1%
#82020000000
0!
0%
#82025000000
1!
1%
#82030000000
0!
0%
#82035000000
1!
1%
#82040000000
0!
0%
#82045000000
1!
1%
#82050000000
0!
0%
#82055000000
1!
1%
#82060000000
0!
0%
#82065000000
1!
1%
#82070000000
0!
0%
#82075000000
1!
1%
#82080000000
0!
0%
#82085000000
1!
1%
#82090000000
0!
0%
#82095000000
1!
1%
#82100000000
0!
0%
#82105000000
1!
1%
#82110000000
0!
0%
#82115000000
1!
1%
#82120000000
0!
0%
#82125000000
1!
1%
#82130000000
0!
0%
#82135000000
1!
1%
#82140000000
0!
0%
#82145000000
1!
1%
#82150000000
0!
0%
#82155000000
1!
1%
#82160000000
0!
0%
#82165000000
1!
1%
#82170000000
0!
0%
#82175000000
1!
1%
#82180000000
0!
0%
#82185000000
1!
1%
#82190000000
0!
0%
#82195000000
1!
1%
#82200000000
0!
0%
#82205000000
1!
1%
#82210000000
0!
0%
#82215000000
1!
1%
#82220000000
0!
0%
#82225000000
1!
1%
#82230000000
0!
0%
#82235000000
1!
1%
#82240000000
0!
0%
#82245000000
1!
1%
#82250000000
0!
0%
#82255000000
1!
1%
#82260000000
0!
0%
#82265000000
1!
1%
#82270000000
0!
0%
#82275000000
1!
1%
#82280000000
0!
0%
#82285000000
1!
1%
#82290000000
0!
0%
#82295000000
1!
1%
#82300000000
0!
0%
#82305000000
1!
1%
#82310000000
0!
0%
#82315000000
1!
1%
#82320000000
0!
0%
#82325000000
1!
1%
#82330000000
0!
0%
#82335000000
1!
1%
#82340000000
0!
0%
#82345000000
1!
1%
#82350000000
0!
0%
#82355000000
1!
1%
#82360000000
0!
0%
#82365000000
1!
1%
#82370000000
0!
0%
#82375000000
1!
1%
#82380000000
0!
0%
#82385000000
1!
1%
#82390000000
0!
0%
#82395000000
1!
1%
#82400000000
0!
0%
#82405000000
1!
1%
#82410000000
0!
0%
#82415000000
1!
1%
#82420000000
0!
0%
#82425000000
1!
1%
#82430000000
0!
0%
#82435000000
1!
1%
#82440000000
0!
0%
#82445000000
1!
1%
#82450000000
0!
0%
#82455000000
1!
1%
#82460000000
0!
0%
#82465000000
1!
1%
#82470000000
0!
0%
#82475000000
1!
1%
#82480000000
0!
0%
#82485000000
1!
1%
#82490000000
0!
0%
#82495000000
1!
1%
#82500000000
0!
0%
#82505000000
1!
1%
#82510000000
0!
0%
#82515000000
1!
1%
#82520000000
0!
0%
#82525000000
1!
1%
#82530000000
0!
0%
#82535000000
1!
1%
#82540000000
0!
0%
#82545000000
1!
1%
#82550000000
0!
0%
#82555000000
1!
1%
#82560000000
0!
0%
#82565000000
1!
1%
#82570000000
0!
0%
#82575000000
1!
1%
#82580000000
0!
0%
#82585000000
1!
1%
#82590000000
0!
0%
#82595000000
1!
1%
#82600000000
0!
0%
#82605000000
1!
1%
#82610000000
0!
0%
#82615000000
1!
1%
#82620000000
0!
0%
#82625000000
1!
1%
#82630000000
0!
0%
#82635000000
1!
1%
#82640000000
0!
0%
#82645000000
1!
1%
#82650000000
0!
0%
#82655000000
1!
1%
#82660000000
0!
0%
#82665000000
1!
1%
#82670000000
0!
0%
#82675000000
1!
1%
#82680000000
0!
0%
#82685000000
1!
1%
#82690000000
0!
0%
#82695000000
1!
1%
#82700000000
0!
0%
#82705000000
1!
1%
#82710000000
0!
0%
#82715000000
1!
1%
#82720000000
0!
0%
#82725000000
1!
1%
#82730000000
0!
0%
#82735000000
1!
1%
#82740000000
0!
0%
#82745000000
1!
1%
#82750000000
0!
0%
#82755000000
1!
1%
#82760000000
0!
0%
#82765000000
1!
1%
#82770000000
0!
0%
#82775000000
1!
1%
#82780000000
0!
0%
#82785000000
1!
1%
#82790000000
0!
0%
#82795000000
1!
1%
#82800000000
0!
0%
#82805000000
1!
1%
#82810000000
0!
0%
#82815000000
1!
1%
#82820000000
0!
0%
#82825000000
1!
1%
#82830000000
0!
0%
#82835000000
1!
1%
#82840000000
0!
0%
#82845000000
1!
1%
#82850000000
0!
0%
#82855000000
1!
1%
#82860000000
0!
0%
#82865000000
1!
1%
#82870000000
0!
0%
#82875000000
1!
1%
#82880000000
0!
0%
#82885000000
1!
1%
#82890000000
0!
0%
#82895000000
1!
1%
#82900000000
0!
0%
#82905000000
1!
1%
#82910000000
0!
0%
#82915000000
1!
1%
#82920000000
0!
0%
#82925000000
1!
1%
#82930000000
0!
0%
#82935000000
1!
1%
#82940000000
0!
0%
#82945000000
1!
1%
#82950000000
0!
0%
#82955000000
1!
1%
#82960000000
0!
0%
#82965000000
1!
1%
#82970000000
0!
0%
#82975000000
1!
1%
#82980000000
0!
0%
#82985000000
1!
1%
#82990000000
0!
0%
#82995000000
1!
1%
#83000000000
0!
0%
#83005000000
1!
1%
#83010000000
0!
0%
#83015000000
1!
1%
#83020000000
0!
0%
#83025000000
1!
1%
#83030000000
0!
0%
#83035000000
1!
1%
#83040000000
0!
0%
#83045000000
1!
1%
#83050000000
0!
0%
#83055000000
1!
1%
#83060000000
0!
0%
#83065000000
1!
1%
#83070000000
0!
0%
#83075000000
1!
1%
#83080000000
0!
0%
#83085000000
1!
1%
#83090000000
0!
0%
#83095000000
1!
1%
#83100000000
0!
0%
#83105000000
1!
1%
#83110000000
0!
0%
#83115000000
1!
1%
#83120000000
0!
0%
#83125000000
1!
1%
#83130000000
0!
0%
#83135000000
1!
1%
#83140000000
0!
0%
#83145000000
1!
1%
#83150000000
0!
0%
#83155000000
1!
1%
#83160000000
0!
0%
#83165000000
1!
1%
#83170000000
0!
0%
#83175000000
1!
1%
#83180000000
0!
0%
#83185000000
1!
1%
#83190000000
0!
0%
#83195000000
1!
1%
#83200000000
0!
0%
#83205000000
1!
1%
#83210000000
0!
0%
#83215000000
1!
1%
#83220000000
0!
0%
#83225000000
1!
1%
#83230000000
0!
0%
#83235000000
1!
1%
#83240000000
0!
0%
#83245000000
1!
1%
#83250000000
0!
0%
#83255000000
1!
1%
#83260000000
0!
0%
#83265000000
1!
1%
#83270000000
0!
0%
#83275000000
1!
1%
#83280000000
0!
0%
#83285000000
1!
1%
#83290000000
0!
0%
#83295000000
1!
1%
#83300000000
0!
0%
#83305000000
1!
1%
#83310000000
0!
0%
#83315000000
1!
1%
#83320000000
0!
0%
#83325000000
1!
1%
#83330000000
0!
0%
#83335000000
1!
1%
#83340000000
0!
0%
#83345000000
1!
1%
#83350000000
0!
0%
#83355000000
1!
1%
#83360000000
0!
0%
#83365000000
1!
1%
#83370000000
0!
0%
#83375000000
1!
1%
#83380000000
0!
0%
#83385000000
1!
1%
#83390000000
0!
0%
#83395000000
1!
1%
#83400000000
0!
0%
#83405000000
1!
1%
#83410000000
0!
0%
#83415000000
1!
1%
#83420000000
0!
0%
#83425000000
1!
1%
#83430000000
0!
0%
#83435000000
1!
1%
#83440000000
0!
0%
#83445000000
1!
1%
#83450000000
0!
0%
#83455000000
1!
1%
#83460000000
0!
0%
#83465000000
1!
1%
#83470000000
0!
0%
#83475000000
1!
1%
#83480000000
0!
0%
#83485000000
1!
1%
#83490000000
0!
0%
#83495000000
1!
1%
#83500000000
0!
0%
#83505000000
1!
1%
#83510000000
0!
0%
#83515000000
1!
1%
#83520000000
0!
0%
#83525000000
1!
1%
#83530000000
0!
0%
#83535000000
1!
1%
#83540000000
0!
0%
#83545000000
1!
1%
#83550000000
0!
0%
#83555000000
1!
1%
#83560000000
0!
0%
#83565000000
1!
1%
#83570000000
0!
0%
#83575000000
1!
1%
#83580000000
0!
0%
#83585000000
1!
1%
#83590000000
0!
0%
#83595000000
1!
1%
#83600000000
0!
0%
#83605000000
1!
1%
#83610000000
0!
0%
#83615000000
1!
1%
#83620000000
0!
0%
#83625000000
1!
1%
#83630000000
0!
0%
#83635000000
1!
1%
#83640000000
0!
0%
#83645000000
1!
1%
#83650000000
0!
0%
#83655000000
1!
1%
#83660000000
0!
0%
#83665000000
1!
1%
#83670000000
0!
0%
#83675000000
1!
1%
#83680000000
0!
0%
#83685000000
1!
1%
#83690000000
0!
0%
#83695000000
1!
1%
#83700000000
0!
0%
#83705000000
1!
1%
#83710000000
0!
0%
#83715000000
1!
1%
#83720000000
0!
0%
#83725000000
1!
1%
#83730000000
0!
0%
#83735000000
1!
1%
#83740000000
0!
0%
#83745000000
1!
1%
#83750000000
0!
0%
#83755000000
1!
1%
#83760000000
0!
0%
#83765000000
1!
1%
#83770000000
0!
0%
#83775000000
1!
1%
#83780000000
0!
0%
#83785000000
1!
1%
#83790000000
0!
0%
#83795000000
1!
1%
#83800000000
0!
0%
#83805000000
1!
1%
#83810000000
0!
0%
#83815000000
1!
1%
#83820000000
0!
0%
#83825000000
1!
1%
#83830000000
0!
0%
#83835000000
1!
1%
#83840000000
0!
0%
#83845000000
1!
1%
#83850000000
0!
0%
#83855000000
1!
1%
#83860000000
0!
0%
#83865000000
1!
1%
#83870000000
0!
0%
#83875000000
1!
1%
#83880000000
0!
0%
#83885000000
1!
1%
#83890000000
0!
0%
#83895000000
1!
1%
#83900000000
0!
0%
#83905000000
1!
1%
#83910000000
0!
0%
#83915000000
1!
1%
#83920000000
0!
0%
#83925000000
1!
1%
#83930000000
0!
0%
#83935000000
1!
1%
#83940000000
0!
0%
#83945000000
1!
1%
#83950000000
0!
0%
#83955000000
1!
1%
#83960000000
0!
0%
#83965000000
1!
1%
#83970000000
0!
0%
#83975000000
1!
1%
#83980000000
0!
0%
#83985000000
1!
1%
#83990000000
0!
0%
#83995000000
1!
1%
#84000000000
0!
0%
#84005000000
1!
1%
#84010000000
0!
0%
#84015000000
1!
1%
#84020000000
0!
0%
#84025000000
1!
1%
#84030000000
0!
0%
#84035000000
1!
1%
#84040000000
0!
0%
#84045000000
1!
1%
#84050000000
0!
0%
#84055000000
1!
1%
#84060000000
0!
0%
#84065000000
1!
1%
#84070000000
0!
0%
#84075000000
1!
1%
#84080000000
0!
0%
#84085000000
1!
1%
#84090000000
0!
0%
#84095000000
1!
1%
#84100000000
0!
0%
#84105000000
1!
1%
#84110000000
0!
0%
#84115000000
1!
1%
#84120000000
0!
0%
#84125000000
1!
1%
#84130000000
0!
0%
#84135000000
1!
1%
#84140000000
0!
0%
#84145000000
1!
1%
#84150000000
0!
0%
#84155000000
1!
1%
#84160000000
0!
0%
#84165000000
1!
1%
#84170000000
0!
0%
#84175000000
1!
1%
#84180000000
0!
0%
#84185000000
1!
1%
#84190000000
0!
0%
#84195000000
1!
1%
#84200000000
0!
0%
#84205000000
1!
1%
#84210000000
0!
0%
#84215000000
1!
1%
#84220000000
0!
0%
#84225000000
1!
1%
#84230000000
0!
0%
#84235000000
1!
1%
#84240000000
0!
0%
#84245000000
1!
1%
#84250000000
0!
0%
#84255000000
1!
1%
#84260000000
0!
0%
#84265000000
1!
1%
#84270000000
0!
0%
#84275000000
1!
1%
#84280000000
0!
0%
#84285000000
1!
1%
#84290000000
0!
0%
#84295000000
1!
1%
#84300000000
0!
0%
#84305000000
1!
1%
#84310000000
0!
0%
#84315000000
1!
1%
#84320000000
0!
0%
#84325000000
1!
1%
#84330000000
0!
0%
#84335000000
1!
1%
#84340000000
0!
0%
#84345000000
1!
1%
#84350000000
0!
0%
#84355000000
1!
1%
#84360000000
0!
0%
#84365000000
1!
1%
#84370000000
0!
0%
#84375000000
1!
1%
#84380000000
0!
0%
#84385000000
1!
1%
#84390000000
0!
0%
#84395000000
1!
1%
#84400000000
0!
0%
#84405000000
1!
1%
#84410000000
0!
0%
#84415000000
1!
1%
#84420000000
0!
0%
#84425000000
1!
1%
#84430000000
0!
0%
#84435000000
1!
1%
#84440000000
0!
0%
#84445000000
1!
1%
#84450000000
0!
0%
#84455000000
1!
1%
#84460000000
0!
0%
#84465000000
1!
1%
#84470000000
0!
0%
#84475000000
1!
1%
#84480000000
0!
0%
#84485000000
1!
1%
#84490000000
0!
0%
#84495000000
1!
1%
#84500000000
0!
0%
#84505000000
1!
1%
#84510000000
0!
0%
#84515000000
1!
1%
#84520000000
0!
0%
#84525000000
1!
1%
#84530000000
0!
0%
#84535000000
1!
1%
#84540000000
0!
0%
#84545000000
1!
1%
#84550000000
0!
0%
#84555000000
1!
1%
#84560000000
0!
0%
#84565000000
1!
1%
#84570000000
0!
0%
#84575000000
1!
1%
#84580000000
0!
0%
#84585000000
1!
1%
#84590000000
0!
0%
#84595000000
1!
1%
#84600000000
0!
0%
#84605000000
1!
1%
#84610000000
0!
0%
#84615000000
1!
1%
#84620000000
0!
0%
#84625000000
1!
1%
#84630000000
0!
0%
#84635000000
1!
1%
#84640000000
0!
0%
#84645000000
1!
1%
#84650000000
0!
0%
#84655000000
1!
1%
#84660000000
0!
0%
#84665000000
1!
1%
#84670000000
0!
0%
#84675000000
1!
1%
#84680000000
0!
0%
#84685000000
1!
1%
#84690000000
0!
0%
#84695000000
1!
1%
#84700000000
0!
0%
#84705000000
1!
1%
#84710000000
0!
0%
#84715000000
1!
1%
#84720000000
0!
0%
#84725000000
1!
1%
#84730000000
0!
0%
#84735000000
1!
1%
#84740000000
0!
0%
#84745000000
1!
1%
#84750000000
0!
0%
#84755000000
1!
1%
#84760000000
0!
0%
#84765000000
1!
1%
#84770000000
0!
0%
#84775000000
1!
1%
#84780000000
0!
0%
#84785000000
1!
1%
#84790000000
0!
0%
#84795000000
1!
1%
#84800000000
0!
0%
#84805000000
1!
1%
#84810000000
0!
0%
#84815000000
1!
1%
#84820000000
0!
0%
#84825000000
1!
1%
#84830000000
0!
0%
#84835000000
1!
1%
#84840000000
0!
0%
#84845000000
1!
1%
#84850000000
0!
0%
#84855000000
1!
1%
#84860000000
0!
0%
#84865000000
1!
1%
#84870000000
0!
0%
#84875000000
1!
1%
#84880000000
0!
0%
#84885000000
1!
1%
#84890000000
0!
0%
#84895000000
1!
1%
#84900000000
0!
0%
#84905000000
1!
1%
#84910000000
0!
0%
#84915000000
1!
1%
#84920000000
0!
0%
#84925000000
1!
1%
#84930000000
0!
0%
#84935000000
1!
1%
#84940000000
0!
0%
#84945000000
1!
1%
#84950000000
0!
0%
#84955000000
1!
1%
#84960000000
0!
0%
#84965000000
1!
1%
#84970000000
0!
0%
#84975000000
1!
1%
#84980000000
0!
0%
#84985000000
1!
1%
#84990000000
0!
0%
#84995000000
1!
1%
#85000000000
0!
0%
#85005000000
1!
1%
#85010000000
0!
0%
#85015000000
1!
1%
#85020000000
0!
0%
#85025000000
1!
1%
#85030000000
0!
0%
#85035000000
1!
1%
#85040000000
0!
0%
#85045000000
1!
1%
#85050000000
0!
0%
#85055000000
1!
1%
#85060000000
0!
0%
#85065000000
1!
1%
#85070000000
0!
0%
#85075000000
1!
1%
#85080000000
0!
0%
#85085000000
1!
1%
#85090000000
0!
0%
#85095000000
1!
1%
#85100000000
0!
0%
#85105000000
1!
1%
#85110000000
0!
0%
#85115000000
1!
1%
#85120000000
0!
0%
#85125000000
1!
1%
#85130000000
0!
0%
#85135000000
1!
1%
#85140000000
0!
0%
#85145000000
1!
1%
#85150000000
0!
0%
#85155000000
1!
1%
#85160000000
0!
0%
#85165000000
1!
1%
#85170000000
0!
0%
#85175000000
1!
1%
#85180000000
0!
0%
#85185000000
1!
1%
#85190000000
0!
0%
#85195000000
1!
1%
#85200000000
0!
0%
#85205000000
1!
1%
#85210000000
0!
0%
#85215000000
1!
1%
#85220000000
0!
0%
#85225000000
1!
1%
#85230000000
0!
0%
#85235000000
1!
1%
#85240000000
0!
0%
#85245000000
1!
1%
#85250000000
0!
0%
#85255000000
1!
1%
#85260000000
0!
0%
#85265000000
1!
1%
#85270000000
0!
0%
#85275000000
1!
1%
#85280000000
0!
0%
#85285000000
1!
1%
#85290000000
0!
0%
#85295000000
1!
1%
#85300000000
0!
0%
#85305000000
1!
1%
#85310000000
0!
0%
#85315000000
1!
1%
#85320000000
0!
0%
#85325000000
1!
1%
#85330000000
0!
0%
#85335000000
1!
1%
#85340000000
0!
0%
#85345000000
1!
1%
#85350000000
0!
0%
#85355000000
1!
1%
#85360000000
0!
0%
#85365000000
1!
1%
#85370000000
0!
0%
#85375000000
1!
1%
#85380000000
0!
0%
#85385000000
1!
1%
#85390000000
0!
0%
#85395000000
1!
1%
#85400000000
0!
0%
#85405000000
1!
1%
#85410000000
0!
0%
#85415000000
1!
1%
#85420000000
0!
0%
#85425000000
1!
1%
#85430000000
0!
0%
#85435000000
1!
1%
#85440000000
0!
0%
#85445000000
1!
1%
#85450000000
0!
0%
#85455000000
1!
1%
#85460000000
0!
0%
#85465000000
1!
1%
#85470000000
0!
0%
#85475000000
1!
1%
#85480000000
0!
0%
#85485000000
1!
1%
#85490000000
0!
0%
#85495000000
1!
1%
#85500000000
0!
0%
#85505000000
1!
1%
#85510000000
0!
0%
#85515000000
1!
1%
#85520000000
0!
0%
#85525000000
1!
1%
#85530000000
0!
0%
#85535000000
1!
1%
#85540000000
0!
0%
#85545000000
1!
1%
#85550000000
0!
0%
#85555000000
1!
1%
#85560000000
0!
0%
#85565000000
1!
1%
#85570000000
0!
0%
#85575000000
1!
1%
#85580000000
0!
0%
#85585000000
1!
1%
#85590000000
0!
0%
#85595000000
1!
1%
#85600000000
0!
0%
#85605000000
1!
1%
#85610000000
0!
0%
#85615000000
1!
1%
#85620000000
0!
0%
#85625000000
1!
1%
#85630000000
0!
0%
#85635000000
1!
1%
#85640000000
0!
0%
#85645000000
1!
1%
#85650000000
0!
0%
#85655000000
1!
1%
#85660000000
0!
0%
#85665000000
1!
1%
#85670000000
0!
0%
#85675000000
1!
1%
#85680000000
0!
0%
#85685000000
1!
1%
#85690000000
0!
0%
#85695000000
1!
1%
#85700000000
0!
0%
#85705000000
1!
1%
#85710000000
0!
0%
#85715000000
1!
1%
#85720000000
0!
0%
#85725000000
1!
1%
#85730000000
0!
0%
#85735000000
1!
1%
#85740000000
0!
0%
#85745000000
1!
1%
#85750000000
0!
0%
#85755000000
1!
1%
#85760000000
0!
0%
#85765000000
1!
1%
#85770000000
0!
0%
#85775000000
1!
1%
#85780000000
0!
0%
#85785000000
1!
1%
#85790000000
0!
0%
#85795000000
1!
1%
#85800000000
0!
0%
#85805000000
1!
1%
#85810000000
0!
0%
#85815000000
1!
1%
#85820000000
0!
0%
#85825000000
1!
1%
#85830000000
0!
0%
#85835000000
1!
1%
#85840000000
0!
0%
#85845000000
1!
1%
#85850000000
0!
0%
#85855000000
1!
1%
#85860000000
0!
0%
#85865000000
1!
1%
#85870000000
0!
0%
#85875000000
1!
1%
#85880000000
0!
0%
#85885000000
1!
1%
#85890000000
0!
0%
#85895000000
1!
1%
#85900000000
0!
0%
#85905000000
1!
1%
#85910000000
0!
0%
#85915000000
1!
1%
#85920000000
0!
0%
#85925000000
1!
1%
#85930000000
0!
0%
#85935000000
1!
1%
#85940000000
0!
0%
#85945000000
1!
1%
#85950000000
0!
0%
#85955000000
1!
1%
#85960000000
0!
0%
#85965000000
1!
1%
#85970000000
0!
0%
#85975000000
1!
1%
#85980000000
0!
0%
#85985000000
1!
1%
#85990000000
0!
0%
#85995000000
1!
1%
#86000000000
0!
0%
#86005000000
1!
1%
#86010000000
0!
0%
#86015000000
1!
1%
#86020000000
0!
0%
#86025000000
1!
1%
#86030000000
0!
0%
#86035000000
1!
1%
#86040000000
0!
0%
#86045000000
1!
1%
#86050000000
0!
0%
#86055000000
1!
1%
#86060000000
0!
0%
#86065000000
1!
1%
#86070000000
0!
0%
#86075000000
1!
1%
#86080000000
0!
0%
#86085000000
1!
1%
#86090000000
0!
0%
#86095000000
1!
1%
#86100000000
0!
0%
#86105000000
1!
1%
#86110000000
0!
0%
#86115000000
1!
1%
#86120000000
0!
0%
#86125000000
1!
1%
#86130000000
0!
0%
#86135000000
1!
1%
#86140000000
0!
0%
#86145000000
1!
1%
#86150000000
0!
0%
#86155000000
1!
1%
#86160000000
0!
0%
#86165000000
1!
1%
#86170000000
0!
0%
#86175000000
1!
1%
#86180000000
0!
0%
#86185000000
1!
1%
#86190000000
0!
0%
#86195000000
1!
1%
#86200000000
0!
0%
#86205000000
1!
1%
#86210000000
0!
0%
#86215000000
1!
1%
#86220000000
0!
0%
#86225000000
1!
1%
#86230000000
0!
0%
#86235000000
1!
1%
#86240000000
0!
0%
#86245000000
1!
1%
#86250000000
0!
0%
#86255000000
1!
1%
#86260000000
0!
0%
#86265000000
1!
1%
#86270000000
0!
0%
#86275000000
1!
1%
#86280000000
0!
0%
#86285000000
1!
1%
#86290000000
0!
0%
#86295000000
1!
1%
#86300000000
0!
0%
#86305000000
1!
1%
#86310000000
0!
0%
#86315000000
1!
1%
#86320000000
0!
0%
#86325000000
1!
1%
#86330000000
0!
0%
#86335000000
1!
1%
#86340000000
0!
0%
#86345000000
1!
1%
#86350000000
0!
0%
#86355000000
1!
1%
#86360000000
0!
0%
#86365000000
1!
1%
#86370000000
0!
0%
#86375000000
1!
1%
#86380000000
0!
0%
#86385000000
1!
1%
#86390000000
0!
0%
#86395000000
1!
1%
#86400000000
0!
0%
#86405000000
1!
1%
#86410000000
0!
0%
#86415000000
1!
1%
#86420000000
0!
0%
#86425000000
1!
1%
#86430000000
0!
0%
#86435000000
1!
1%
#86440000000
0!
0%
#86445000000
1!
1%
#86450000000
0!
0%
#86455000000
1!
1%
#86460000000
0!
0%
#86465000000
1!
1%
#86470000000
0!
0%
#86475000000
1!
1%
#86480000000
0!
0%
#86485000000
1!
1%
#86490000000
0!
0%
#86495000000
1!
1%
#86500000000
0!
0%
#86505000000
1!
1%
#86510000000
0!
0%
#86515000000
1!
1%
#86520000000
0!
0%
#86525000000
1!
1%
#86530000000
0!
0%
#86535000000
1!
1%
#86540000000
0!
0%
#86545000000
1!
1%
#86550000000
0!
0%
#86555000000
1!
1%
#86560000000
0!
0%
#86565000000
1!
1%
#86570000000
0!
0%
#86575000000
1!
1%
#86580000000
0!
0%
#86585000000
1!
1%
#86590000000
0!
0%
#86595000000
1!
1%
#86600000000
0!
0%
#86605000000
1!
1%
#86610000000
0!
0%
#86615000000
1!
1%
#86620000000
0!
0%
#86625000000
1!
1%
#86630000000
0!
0%
#86635000000
1!
1%
#86640000000
0!
0%
#86645000000
1!
1%
#86650000000
0!
0%
#86655000000
1!
1%
#86660000000
0!
0%
#86665000000
1!
1%
#86670000000
0!
0%
#86675000000
1!
1%
#86680000000
0!
0%
#86685000000
1!
1%
#86690000000
0!
0%
#86695000000
1!
1%
#86700000000
0!
0%
#86705000000
1!
1%
#86710000000
0!
0%
#86715000000
1!
1%
#86720000000
0!
0%
#86725000000
1!
1%
#86730000000
0!
0%
#86735000000
1!
1%
#86740000000
0!
0%
#86745000000
1!
1%
#86750000000
0!
0%
#86755000000
1!
1%
#86760000000
0!
0%
#86765000000
1!
1%
#86770000000
0!
0%
#86775000000
1!
1%
#86780000000
0!
0%
#86785000000
1!
1%
#86790000000
0!
0%
#86795000000
1!
1%
#86800000000
0!
0%
#86805000000
1!
1%
#86810000000
0!
0%
#86815000000
1!
1%
#86820000000
0!
0%
#86825000000
1!
1%
#86830000000
0!
0%
#86835000000
1!
1%
#86840000000
0!
0%
#86845000000
1!
1%
#86850000000
0!
0%
#86855000000
1!
1%
#86860000000
0!
0%
#86865000000
1!
1%
#86870000000
0!
0%
#86875000000
1!
1%
#86880000000
0!
0%
#86885000000
1!
1%
#86890000000
0!
0%
#86895000000
1!
1%
#86900000000
0!
0%
#86905000000
1!
1%
#86910000000
0!
0%
#86915000000
1!
1%
#86920000000
0!
0%
#86925000000
1!
1%
#86930000000
0!
0%
#86935000000
1!
1%
#86940000000
0!
0%
#86945000000
1!
1%
#86950000000
0!
0%
#86955000000
1!
1%
#86960000000
0!
0%
#86965000000
1!
1%
#86970000000
0!
0%
#86975000000
1!
1%
#86980000000
0!
0%
#86985000000
1!
1%
#86990000000
0!
0%
#86995000000
1!
1%
#87000000000
0!
0%
#87005000000
1!
1%
#87010000000
0!
0%
#87015000000
1!
1%
#87020000000
0!
0%
#87025000000
1!
1%
#87030000000
0!
0%
#87035000000
1!
1%
#87040000000
0!
0%
#87045000000
1!
1%
#87050000000
0!
0%
#87055000000
1!
1%
#87060000000
0!
0%
#87065000000
1!
1%
#87070000000
0!
0%
#87075000000
1!
1%
#87080000000
0!
0%
#87085000000
1!
1%
#87090000000
0!
0%
#87095000000
1!
1%
#87100000000
0!
0%
#87105000000
1!
1%
#87110000000
0!
0%
#87115000000
1!
1%
#87120000000
0!
0%
#87125000000
1!
1%
#87130000000
0!
0%
#87135000000
1!
1%
#87140000000
0!
0%
#87145000000
1!
1%
#87150000000
0!
0%
#87155000000
1!
1%
#87160000000
0!
0%
#87165000000
1!
1%
#87170000000
0!
0%
#87175000000
1!
1%
#87180000000
0!
0%
#87185000000
1!
1%
#87190000000
0!
0%
#87195000000
1!
1%
#87200000000
0!
0%
#87205000000
1!
1%
#87210000000
0!
0%
#87215000000
1!
1%
#87220000000
0!
0%
#87225000000
1!
1%
#87230000000
0!
0%
#87235000000
1!
1%
#87240000000
0!
0%
#87245000000
1!
1%
#87250000000
0!
0%
#87255000000
1!
1%
#87260000000
0!
0%
#87265000000
1!
1%
#87270000000
0!
0%
#87275000000
1!
1%
#87280000000
0!
0%
#87285000000
1!
1%
#87290000000
0!
0%
#87295000000
1!
1%
#87300000000
0!
0%
#87305000000
1!
1%
#87310000000
0!
0%
#87315000000
1!
1%
#87320000000
0!
0%
#87325000000
1!
1%
#87330000000
0!
0%
#87335000000
1!
1%
#87340000000
0!
0%
#87345000000
1!
1%
#87350000000
0!
0%
#87355000000
1!
1%
#87360000000
0!
0%
#87365000000
1!
1%
#87370000000
0!
0%
#87375000000
1!
1%
#87380000000
0!
0%
#87385000000
1!
1%
#87390000000
0!
0%
#87395000000
1!
1%
#87400000000
0!
0%
#87405000000
1!
1%
#87410000000
0!
0%
#87415000000
1!
1%
#87420000000
0!
0%
#87425000000
1!
1%
#87430000000
0!
0%
#87435000000
1!
1%
#87440000000
0!
0%
#87445000000
1!
1%
#87450000000
0!
0%
#87455000000
1!
1%
#87460000000
0!
0%
#87465000000
1!
1%
#87470000000
0!
0%
#87475000000
1!
1%
#87480000000
0!
0%
#87485000000
1!
1%
#87490000000
0!
0%
#87495000000
1!
1%
#87500000000
0!
0%
#87505000000
1!
1%
#87510000000
0!
0%
#87515000000
1!
1%
#87520000000
0!
0%
#87525000000
1!
1%
#87530000000
0!
0%
#87535000000
1!
1%
#87540000000
0!
0%
#87545000000
1!
1%
#87550000000
0!
0%
#87555000000
1!
1%
#87560000000
0!
0%
#87565000000
1!
1%
#87570000000
0!
0%
#87575000000
1!
1%
#87580000000
0!
0%
#87585000000
1!
1%
#87590000000
0!
0%
#87595000000
1!
1%
#87600000000
0!
0%
#87605000000
1!
1%
#87610000000
0!
0%
#87615000000
1!
1%
#87620000000
0!
0%
#87625000000
1!
1%
#87630000000
0!
0%
#87635000000
1!
1%
#87640000000
0!
0%
#87645000000
1!
1%
#87650000000
0!
0%
#87655000000
1!
1%
#87660000000
0!
0%
#87665000000
1!
1%
#87670000000
0!
0%
#87675000000
1!
1%
#87680000000
0!
0%
#87685000000
1!
1%
#87690000000
0!
0%
#87695000000
1!
1%
#87700000000
0!
0%
#87705000000
1!
1%
#87710000000
0!
0%
#87715000000
1!
1%
#87720000000
0!
0%
#87725000000
1!
1%
#87730000000
0!
0%
#87735000000
1!
1%
#87740000000
0!
0%
#87745000000
1!
1%
#87750000000
0!
0%
#87755000000
1!
1%
#87760000000
0!
0%
#87765000000
1!
1%
#87770000000
0!
0%
#87775000000
1!
1%
#87780000000
0!
0%
#87785000000
1!
1%
#87790000000
0!
0%
#87795000000
1!
1%
#87800000000
0!
0%
#87805000000
1!
1%
#87810000000
0!
0%
#87815000000
1!
1%
#87820000000
0!
0%
#87825000000
1!
1%
#87830000000
0!
0%
#87835000000
1!
1%
#87840000000
0!
0%
#87845000000
1!
1%
#87850000000
0!
0%
#87855000000
1!
1%
#87860000000
0!
0%
#87865000000
1!
1%
#87870000000
0!
0%
#87875000000
1!
1%
#87880000000
0!
0%
#87885000000
1!
1%
#87890000000
0!
0%
#87895000000
1!
1%
#87900000000
0!
0%
#87905000000
1!
1%
#87910000000
0!
0%
#87915000000
1!
1%
#87920000000
0!
0%
#87925000000
1!
1%
#87930000000
0!
0%
#87935000000
1!
1%
#87940000000
0!
0%
#87945000000
1!
1%
#87950000000
0!
0%
#87955000000
1!
1%
#87960000000
0!
0%
#87965000000
1!
1%
#87970000000
0!
0%
#87975000000
1!
1%
#87980000000
0!
0%
#87985000000
1!
1%
#87990000000
0!
0%
#87995000000
1!
1%
#88000000000
0!
0%
#88005000000
1!
1%
#88010000000
0!
0%
#88015000000
1!
1%
#88020000000
0!
0%
#88025000000
1!
1%
#88030000000
0!
0%
#88035000000
1!
1%
#88040000000
0!
0%
#88045000000
1!
1%
#88050000000
0!
0%
#88055000000
1!
1%
#88060000000
0!
0%
#88065000000
1!
1%
#88070000000
0!
0%
#88075000000
1!
1%
#88080000000
0!
0%
#88085000000
1!
1%
#88090000000
0!
0%
#88095000000
1!
1%
#88100000000
0!
0%
#88105000000
1!
1%
#88110000000
0!
0%
#88115000000
1!
1%
#88120000000
0!
0%
#88125000000
1!
1%
#88130000000
0!
0%
#88135000000
1!
1%
#88140000000
0!
0%
#88145000000
1!
1%
#88150000000
0!
0%
#88155000000
1!
1%
#88160000000
0!
0%
#88165000000
1!
1%
#88170000000
0!
0%
#88175000000
1!
1%
#88180000000
0!
0%
#88185000000
1!
1%
#88190000000
0!
0%
#88195000000
1!
1%
#88200000000
0!
0%
#88205000000
1!
1%
#88210000000
0!
0%
#88215000000
1!
1%
#88220000000
0!
0%
#88225000000
1!
1%
#88230000000
0!
0%
#88235000000
1!
1%
#88240000000
0!
0%
#88245000000
1!
1%
#88250000000
0!
0%
#88255000000
1!
1%
#88260000000
0!
0%
#88265000000
1!
1%
#88270000000
0!
0%
#88275000000
1!
1%
#88280000000
0!
0%
#88285000000
1!
1%
#88290000000
0!
0%
#88295000000
1!
1%
#88300000000
0!
0%
#88305000000
1!
1%
#88310000000
0!
0%
#88315000000
1!
1%
#88320000000
0!
0%
#88325000000
1!
1%
#88330000000
0!
0%
#88335000000
1!
1%
#88340000000
0!
0%
#88345000000
1!
1%
#88350000000
0!
0%
#88355000000
1!
1%
#88360000000
0!
0%
#88365000000
1!
1%
#88370000000
0!
0%
#88375000000
1!
1%
#88380000000
0!
0%
#88385000000
1!
1%
#88390000000
0!
0%
#88395000000
1!
1%
#88400000000
0!
0%
#88405000000
1!
1%
#88410000000
0!
0%
#88415000000
1!
1%
#88420000000
0!
0%
#88425000000
1!
1%
#88430000000
0!
0%
#88435000000
1!
1%
#88440000000
0!
0%
#88445000000
1!
1%
#88450000000
0!
0%
#88455000000
1!
1%
#88460000000
0!
0%
#88465000000
1!
1%
#88470000000
0!
0%
#88475000000
1!
1%
#88480000000
0!
0%
#88485000000
1!
1%
#88490000000
0!
0%
#88495000000
1!
1%
#88500000000
0!
0%
#88505000000
1!
1%
#88510000000
0!
0%
#88515000000
1!
1%
#88520000000
0!
0%
#88525000000
1!
1%
#88530000000
0!
0%
#88535000000
1!
1%
#88540000000
0!
0%
#88545000000
1!
1%
#88550000000
0!
0%
#88555000000
1!
1%
#88560000000
0!
0%
#88565000000
1!
1%
#88570000000
0!
0%
#88575000000
1!
1%
#88580000000
0!
0%
#88585000000
1!
1%
#88590000000
0!
0%
#88595000000
1!
1%
#88600000000
0!
0%
#88605000000
1!
1%
#88610000000
0!
0%
#88615000000
1!
1%
#88620000000
0!
0%
#88625000000
1!
1%
#88630000000
0!
0%
#88635000000
1!
1%
#88640000000
0!
0%
#88645000000
1!
1%
#88650000000
0!
0%
#88655000000
1!
1%
#88660000000
0!
0%
#88665000000
1!
1%
#88670000000
0!
0%
#88675000000
1!
1%
#88680000000
0!
0%
#88685000000
1!
1%
#88690000000
0!
0%
#88695000000
1!
1%
#88700000000
0!
0%
#88705000000
1!
1%
#88710000000
0!
0%
#88715000000
1!
1%
#88720000000
0!
0%
#88725000000
1!
1%
#88730000000
0!
0%
#88735000000
1!
1%
#88740000000
0!
0%
#88745000000
1!
1%
#88750000000
0!
0%
#88755000000
1!
1%
#88760000000
0!
0%
#88765000000
1!
1%
#88770000000
0!
0%
#88775000000
1!
1%
#88780000000
0!
0%
#88785000000
1!
1%
#88790000000
0!
0%
#88795000000
1!
1%
#88800000000
0!
0%
#88805000000
1!
1%
#88810000000
0!
0%
#88815000000
1!
1%
#88820000000
0!
0%
#88825000000
1!
1%
#88830000000
0!
0%
#88835000000
1!
1%
#88840000000
0!
0%
#88845000000
1!
1%
#88850000000
0!
0%
#88855000000
1!
1%
#88860000000
0!
0%
#88865000000
1!
1%
#88870000000
0!
0%
#88875000000
1!
1%
#88880000000
0!
0%
#88885000000
1!
1%
#88890000000
0!
0%
#88895000000
1!
1%
#88900000000
0!
0%
#88905000000
1!
1%
#88910000000
0!
0%
#88915000000
1!
1%
#88920000000
0!
0%
#88925000000
1!
1%
#88930000000
0!
0%
#88935000000
1!
1%
#88940000000
0!
0%
#88945000000
1!
1%
#88950000000
0!
0%
#88955000000
1!
1%
#88960000000
0!
0%
#88965000000
1!
1%
#88970000000
0!
0%
#88975000000
1!
1%
#88980000000
0!
0%
#88985000000
1!
1%
#88990000000
0!
0%
#88995000000
1!
1%
#89000000000
0!
0%
#89005000000
1!
1%
#89010000000
0!
0%
#89015000000
1!
1%
#89020000000
0!
0%
#89025000000
1!
1%
#89030000000
0!
0%
#89035000000
1!
1%
#89040000000
0!
0%
#89045000000
1!
1%
#89050000000
0!
0%
#89055000000
1!
1%
#89060000000
0!
0%
#89065000000
1!
1%
#89070000000
0!
0%
#89075000000
1!
1%
#89080000000
0!
0%
#89085000000
1!
1%
#89090000000
0!
0%
#89095000000
1!
1%
#89100000000
0!
0%
#89105000000
1!
1%
#89110000000
0!
0%
#89115000000
1!
1%
#89120000000
0!
0%
#89125000000
1!
1%
#89130000000
0!
0%
#89135000000
1!
1%
#89140000000
0!
0%
#89145000000
1!
1%
#89150000000
0!
0%
#89155000000
1!
1%
#89160000000
0!
0%
#89165000000
1!
1%
#89170000000
0!
0%
#89175000000
1!
1%
#89180000000
0!
0%
#89185000000
1!
1%
#89190000000
0!
0%
#89195000000
1!
1%
#89200000000
0!
0%
#89205000000
1!
1%
#89210000000
0!
0%
#89215000000
1!
1%
#89220000000
0!
0%
#89225000000
1!
1%
#89230000000
0!
0%
#89235000000
1!
1%
#89240000000
0!
0%
#89245000000
1!
1%
#89250000000
0!
0%
#89255000000
1!
1%
#89260000000
0!
0%
#89265000000
1!
1%
#89270000000
0!
0%
#89275000000
1!
1%
#89280000000
0!
0%
#89285000000
1!
1%
#89290000000
0!
0%
#89295000000
1!
1%
#89300000000
0!
0%
#89305000000
1!
1%
#89310000000
0!
0%
#89315000000
1!
1%
#89320000000
0!
0%
#89325000000
1!
1%
#89330000000
0!
0%
#89335000000
1!
1%
#89340000000
0!
0%
#89345000000
1!
1%
#89350000000
0!
0%
#89355000000
1!
1%
#89360000000
0!
0%
#89365000000
1!
1%
#89370000000
0!
0%
#89375000000
1!
1%
#89380000000
0!
0%
#89385000000
1!
1%
#89390000000
0!
0%
#89395000000
1!
1%
#89400000000
0!
0%
#89405000000
1!
1%
#89410000000
0!
0%
#89415000000
1!
1%
#89420000000
0!
0%
#89425000000
1!
1%
#89430000000
0!
0%
#89435000000
1!
1%
#89440000000
0!
0%
#89445000000
1!
1%
#89450000000
0!
0%
#89455000000
1!
1%
#89460000000
0!
0%
#89465000000
1!
1%
#89470000000
0!
0%
#89475000000
1!
1%
#89480000000
0!
0%
#89485000000
1!
1%
#89490000000
0!
0%
#89495000000
1!
1%
#89500000000
0!
0%
#89505000000
1!
1%
#89510000000
0!
0%
#89515000000
1!
1%
#89520000000
0!
0%
#89525000000
1!
1%
#89530000000
0!
0%
#89535000000
1!
1%
#89540000000
0!
0%
#89545000000
1!
1%
#89550000000
0!
0%
#89555000000
1!
1%
#89560000000
0!
0%
#89565000000
1!
1%
#89570000000
0!
0%
#89575000000
1!
1%
#89580000000
0!
0%
#89585000000
1!
1%
#89590000000
0!
0%
#89595000000
1!
1%
#89600000000
0!
0%
#89605000000
1!
1%
#89610000000
0!
0%
#89615000000
1!
1%
#89620000000
0!
0%
#89625000000
1!
1%
#89630000000
0!
0%
#89635000000
1!
1%
#89640000000
0!
0%
#89645000000
1!
1%
#89650000000
0!
0%
#89655000000
1!
1%
#89660000000
0!
0%
#89665000000
1!
1%
#89670000000
0!
0%
#89675000000
1!
1%
#89680000000
0!
0%
#89685000000
1!
1%
#89690000000
0!
0%
#89695000000
1!
1%
#89700000000
0!
0%
#89705000000
1!
1%
#89710000000
0!
0%
#89715000000
1!
1%
#89720000000
0!
0%
#89725000000
1!
1%
#89730000000
0!
0%
#89735000000
1!
1%
#89740000000
0!
0%
#89745000000
1!
1%
#89750000000
0!
0%
#89755000000
1!
1%
#89760000000
0!
0%
#89765000000
1!
1%
#89770000000
0!
0%
#89775000000
1!
1%
#89780000000
0!
0%
#89785000000
1!
1%
#89790000000
0!
0%
#89795000000
1!
1%
#89800000000
0!
0%
#89805000000
1!
1%
#89810000000
0!
0%
#89815000000
1!
1%
#89820000000
0!
0%
#89825000000
1!
1%
#89830000000
0!
0%
#89835000000
1!
1%
#89840000000
0!
0%
#89845000000
1!
1%
#89850000000
0!
0%
#89855000000
1!
1%
#89860000000
0!
0%
#89865000000
1!
1%
#89870000000
0!
0%
#89875000000
1!
1%
#89880000000
0!
0%
#89885000000
1!
1%
#89890000000
0!
0%
#89895000000
1!
1%
#89900000000
0!
0%
#89905000000
1!
1%
#89910000000
0!
0%
#89915000000
1!
1%
#89920000000
0!
0%
#89925000000
1!
1%
#89930000000
0!
0%
#89935000000
1!
1%
#89940000000
0!
0%
#89945000000
1!
1%
#89950000000
0!
0%
#89955000000
1!
1%
#89960000000
0!
0%
#89965000000
1!
1%
#89970000000
0!
0%
#89975000000
1!
1%
#89980000000
0!
0%
#89985000000
1!
1%
#89990000000
0!
0%
#89995000000
1!
1%
#90000000000
0!
0%
#90005000000
1!
1%
#90010000000
0!
0%
#90015000000
1!
1%
#90020000000
0!
0%
#90025000000
1!
1%
#90030000000
0!
0%
#90035000000
1!
1%
#90040000000
0!
0%
#90045000000
1!
1%
#90050000000
0!
0%
#90055000000
1!
1%
#90060000000
0!
0%
#90065000000
1!
1%
#90070000000
0!
0%
#90075000000
1!
1%
#90080000000
0!
0%
#90085000000
1!
1%
#90090000000
0!
0%
#90095000000
1!
1%
#90100000000
0!
0%
#90105000000
1!
1%
#90110000000
0!
0%
#90115000000
1!
1%
#90120000000
0!
0%
#90125000000
1!
1%
#90130000000
0!
0%
#90135000000
1!
1%
#90140000000
0!
0%
#90145000000
1!
1%
#90150000000
0!
0%
#90155000000
1!
1%
#90160000000
0!
0%
#90165000000
1!
1%
#90170000000
0!
0%
#90175000000
1!
1%
#90180000000
0!
0%
#90185000000
1!
1%
#90190000000
0!
0%
#90195000000
1!
1%
#90200000000
0!
0%
#90205000000
1!
1%
#90210000000
0!
0%
#90215000000
1!
1%
#90220000000
0!
0%
#90225000000
1!
1%
#90230000000
0!
0%
#90235000000
1!
1%
#90240000000
0!
0%
#90245000000
1!
1%
#90250000000
0!
0%
#90255000000
1!
1%
#90260000000
0!
0%
#90265000000
1!
1%
#90270000000
0!
0%
#90275000000
1!
1%
#90280000000
0!
0%
#90285000000
1!
1%
#90290000000
0!
0%
#90295000000
1!
1%
#90300000000
0!
0%
#90305000000
1!
1%
#90310000000
0!
0%
#90315000000
1!
1%
#90320000000
0!
0%
#90325000000
1!
1%
#90330000000
0!
0%
#90335000000
1!
1%
#90340000000
0!
0%
#90345000000
1!
1%
#90350000000
0!
0%
#90355000000
1!
1%
#90360000000
0!
0%
#90365000000
1!
1%
#90370000000
0!
0%
#90375000000
1!
1%
#90380000000
0!
0%
#90385000000
1!
1%
#90390000000
0!
0%
#90395000000
1!
1%
#90400000000
0!
0%
#90405000000
1!
1%
#90410000000
0!
0%
#90415000000
1!
1%
#90420000000
0!
0%
#90425000000
1!
1%
#90430000000
0!
0%
#90435000000
1!
1%
#90440000000
0!
0%
#90445000000
1!
1%
#90450000000
0!
0%
#90455000000
1!
1%
#90460000000
0!
0%
#90465000000
1!
1%
#90470000000
0!
0%
#90475000000
1!
1%
#90480000000
0!
0%
#90485000000
1!
1%
#90490000000
0!
0%
#90495000000
1!
1%
#90500000000
0!
0%
#90505000000
1!
1%
#90510000000
0!
0%
#90515000000
1!
1%
#90520000000
0!
0%
#90525000000
1!
1%
#90530000000
0!
0%
#90535000000
1!
1%
#90540000000
0!
0%
#90545000000
1!
1%
#90550000000
0!
0%
#90555000000
1!
1%
#90560000000
0!
0%
#90565000000
1!
1%
#90570000000
0!
0%
#90575000000
1!
1%
#90580000000
0!
0%
#90585000000
1!
1%
#90590000000
0!
0%
#90595000000
1!
1%
#90600000000
0!
0%
#90605000000
1!
1%
#90610000000
0!
0%
#90615000000
1!
1%
#90620000000
0!
0%
#90625000000
1!
1%
#90630000000
0!
0%
#90635000000
1!
1%
#90640000000
0!
0%
#90645000000
1!
1%
#90650000000
0!
0%
#90655000000
1!
1%
#90660000000
0!
0%
#90665000000
1!
1%
#90670000000
0!
0%
#90675000000
1!
1%
#90680000000
0!
0%
#90685000000
1!
1%
#90690000000
0!
0%
#90695000000
1!
1%
#90700000000
0!
0%
#90705000000
1!
1%
#90710000000
0!
0%
#90715000000
1!
1%
#90720000000
0!
0%
#90725000000
1!
1%
#90730000000
0!
0%
#90735000000
1!
1%
#90740000000
0!
0%
#90745000000
1!
1%
#90750000000
0!
0%
#90755000000
1!
1%
#90760000000
0!
0%
#90765000000
1!
1%
#90770000000
0!
0%
#90775000000
1!
1%
#90780000000
0!
0%
#90785000000
1!
1%
#90790000000
0!
0%
#90795000000
1!
1%
#90800000000
0!
0%
#90805000000
1!
1%
#90810000000
0!
0%
#90815000000
1!
1%
#90820000000
0!
0%
#90825000000
1!
1%
#90830000000
0!
0%
#90835000000
1!
1%
#90840000000
0!
0%
#90845000000
1!
1%
#90850000000
0!
0%
#90855000000
1!
1%
#90860000000
0!
0%
#90865000000
1!
1%
#90870000000
0!
0%
#90875000000
1!
1%
#90880000000
0!
0%
#90885000000
1!
1%
#90890000000
0!
0%
#90895000000
1!
1%
#90900000000
0!
0%
#90905000000
1!
1%
#90910000000
0!
0%
#90915000000
1!
1%
#90920000000
0!
0%
#90925000000
1!
1%
#90930000000
0!
0%
#90935000000
1!
1%
#90940000000
0!
0%
#90945000000
1!
1%
#90950000000
0!
0%
#90955000000
1!
1%
#90960000000
0!
0%
#90965000000
1!
1%
#90970000000
0!
0%
#90975000000
1!
1%
#90980000000
0!
0%
#90985000000
1!
1%
#90990000000
0!
0%
#90995000000
1!
1%
#91000000000
0!
0%
#91005000000
1!
1%
#91010000000
0!
0%
#91015000000
1!
1%
#91020000000
0!
0%
#91025000000
1!
1%
#91030000000
0!
0%
#91035000000
1!
1%
#91040000000
0!
0%
#91045000000
1!
1%
#91050000000
0!
0%
#91055000000
1!
1%
#91060000000
0!
0%
#91065000000
1!
1%
#91070000000
0!
0%
#91075000000
1!
1%
#91080000000
0!
0%
#91085000000
1!
1%
#91090000000
0!
0%
#91095000000
1!
1%
#91100000000
0!
0%
#91105000000
1!
1%
#91110000000
0!
0%
#91115000000
1!
1%
#91120000000
0!
0%
#91125000000
1!
1%
#91130000000
0!
0%
#91135000000
1!
1%
#91140000000
0!
0%
#91145000000
1!
1%
#91150000000
0!
0%
#91155000000
1!
1%
#91160000000
0!
0%
#91165000000
1!
1%
#91170000000
0!
0%
#91175000000
1!
1%
#91180000000
0!
0%
#91185000000
1!
1%
#91190000000
0!
0%
#91195000000
1!
1%
#91200000000
0!
0%
#91205000000
1!
1%
#91210000000
0!
0%
#91215000000
1!
1%
#91220000000
0!
0%
#91225000000
1!
1%
#91230000000
0!
0%
#91235000000
1!
1%
#91240000000
0!
0%
#91245000000
1!
1%
#91250000000
0!
0%
#91255000000
1!
1%
#91260000000
0!
0%
#91265000000
1!
1%
#91270000000
0!
0%
#91275000000
1!
1%
#91280000000
0!
0%
#91285000000
1!
1%
#91290000000
0!
0%
#91295000000
1!
1%
#91300000000
0!
0%
#91305000000
1!
1%
#91310000000
0!
0%
#91315000000
1!
1%
#91320000000
0!
0%
#91325000000
1!
1%
#91330000000
0!
0%
#91335000000
1!
1%
#91340000000
0!
0%
#91345000000
1!
1%
#91350000000
0!
0%
#91355000000
1!
1%
#91360000000
0!
0%
#91365000000
1!
1%
#91370000000
0!
0%
#91375000000
1!
1%
#91380000000
0!
0%
#91385000000
1!
1%
#91390000000
0!
0%
#91395000000
1!
1%
#91400000000
0!
0%
#91405000000
1!
1%
#91410000000
0!
0%
#91415000000
1!
1%
#91420000000
0!
0%
#91425000000
1!
1%
#91430000000
0!
0%
#91435000000
1!
1%
#91440000000
0!
0%
#91445000000
1!
1%
#91450000000
0!
0%
#91455000000
1!
1%
#91460000000
0!
0%
#91465000000
1!
1%
#91470000000
0!
0%
#91475000000
1!
1%
#91480000000
0!
0%
#91485000000
1!
1%
#91490000000
0!
0%
#91495000000
1!
1%
#91500000000
0!
0%
#91505000000
1!
1%
#91510000000
0!
0%
#91515000000
1!
1%
#91520000000
0!
0%
#91525000000
1!
1%
#91530000000
0!
0%
#91535000000
1!
1%
#91540000000
0!
0%
#91545000000
1!
1%
#91550000000
0!
0%
#91555000000
1!
1%
#91560000000
0!
0%
#91565000000
1!
1%
#91570000000
0!
0%
#91575000000
1!
1%
#91580000000
0!
0%
#91585000000
1!
1%
#91590000000
0!
0%
#91595000000
1!
1%
#91600000000
0!
0%
#91605000000
1!
1%
#91610000000
0!
0%
#91615000000
1!
1%
#91620000000
0!
0%
#91625000000
1!
1%
#91630000000
0!
0%
#91635000000
1!
1%
#91640000000
0!
0%
#91645000000
1!
1%
#91650000000
0!
0%
#91655000000
1!
1%
#91660000000
0!
0%
#91665000000
1!
1%
#91670000000
0!
0%
#91675000000
1!
1%
#91680000000
0!
0%
#91685000000
1!
1%
#91690000000
0!
0%
#91695000000
1!
1%
#91700000000
0!
0%
#91705000000
1!
1%
#91710000000
0!
0%
#91715000000
1!
1%
#91720000000
0!
0%
#91725000000
1!
1%
#91730000000
0!
0%
#91735000000
1!
1%
#91740000000
0!
0%
#91745000000
1!
1%
#91750000000
0!
0%
#91755000000
1!
1%
#91760000000
0!
0%
#91765000000
1!
1%
#91770000000
0!
0%
#91775000000
1!
1%
#91780000000
0!
0%
#91785000000
1!
1%
#91790000000
0!
0%
#91795000000
1!
1%
#91800000000
0!
0%
#91805000000
1!
1%
#91810000000
0!
0%
#91815000000
1!
1%
#91820000000
0!
0%
#91825000000
1!
1%
#91830000000
0!
0%
#91835000000
1!
1%
#91840000000
0!
0%
#91845000000
1!
1%
#91850000000
0!
0%
#91855000000
1!
1%
#91860000000
0!
0%
#91865000000
1!
1%
#91870000000
0!
0%
#91875000000
1!
1%
#91880000000
0!
0%
#91885000000
1!
1%
#91890000000
0!
0%
#91895000000
1!
1%
#91900000000
0!
0%
#91905000000
1!
1%
#91910000000
0!
0%
#91915000000
1!
1%
#91920000000
0!
0%
#91925000000
1!
1%
#91930000000
0!
0%
#91935000000
1!
1%
#91940000000
0!
0%
#91945000000
1!
1%
#91950000000
0!
0%
#91955000000
1!
1%
#91960000000
0!
0%
#91965000000
1!
1%
#91970000000
0!
0%
#91975000000
1!
1%
#91980000000
0!
0%
#91985000000
1!
1%
#91990000000
0!
0%
#91995000000
1!
1%
#92000000000
0!
0%
#92005000000
1!
1%
#92010000000
0!
0%
#92015000000
1!
1%
#92020000000
0!
0%
#92025000000
1!
1%
#92030000000
0!
0%
#92035000000
1!
1%
#92040000000
0!
0%
#92045000000
1!
1%
#92050000000
0!
0%
#92055000000
1!
1%
#92060000000
0!
0%
#92065000000
1!
1%
#92070000000
0!
0%
#92075000000
1!
1%
#92080000000
0!
0%
#92085000000
1!
1%
#92090000000
0!
0%
#92095000000
1!
1%
#92100000000
0!
0%
#92105000000
1!
1%
#92110000000
0!
0%
#92115000000
1!
1%
#92120000000
0!
0%
#92125000000
1!
1%
#92130000000
0!
0%
#92135000000
1!
1%
#92140000000
0!
0%
#92145000000
1!
1%
#92150000000
0!
0%
#92155000000
1!
1%
#92160000000
0!
0%
#92165000000
1!
1%
#92170000000
0!
0%
#92175000000
1!
1%
#92180000000
0!
0%
#92185000000
1!
1%
#92190000000
0!
0%
#92195000000
1!
1%
#92200000000
0!
0%
#92205000000
1!
1%
#92210000000
0!
0%
#92215000000
1!
1%
#92220000000
0!
0%
#92225000000
1!
1%
#92230000000
0!
0%
#92235000000
1!
1%
#92240000000
0!
0%
#92245000000
1!
1%
#92250000000
0!
0%
#92255000000
1!
1%
#92260000000
0!
0%
#92265000000
1!
1%
#92270000000
0!
0%
#92275000000
1!
1%
#92280000000
0!
0%
#92285000000
1!
1%
#92290000000
0!
0%
#92295000000
1!
1%
#92300000000
0!
0%
#92305000000
1!
1%
#92310000000
0!
0%
#92315000000
1!
1%
#92320000000
0!
0%
#92325000000
1!
1%
#92330000000
0!
0%
#92335000000
1!
1%
#92340000000
0!
0%
#92345000000
1!
1%
#92350000000
0!
0%
#92355000000
1!
1%
#92360000000
0!
0%
#92365000000
1!
1%
#92370000000
0!
0%
#92375000000
1!
1%
#92380000000
0!
0%
#92385000000
1!
1%
#92390000000
0!
0%
#92395000000
1!
1%
#92400000000
0!
0%
#92405000000
1!
1%
#92410000000
0!
0%
#92415000000
1!
1%
#92420000000
0!
0%
#92425000000
1!
1%
#92430000000
0!
0%
#92435000000
1!
1%
#92440000000
0!
0%
#92445000000
1!
1%
#92450000000
0!
0%
#92455000000
1!
1%
#92460000000
0!
0%
#92465000000
1!
1%
#92470000000
0!
0%
#92475000000
1!
1%
#92480000000
0!
0%
#92485000000
1!
1%
#92490000000
0!
0%
#92495000000
1!
1%
#92500000000
0!
0%
#92505000000
1!
1%
#92510000000
0!
0%
#92515000000
1!
1%
#92520000000
0!
0%
#92525000000
1!
1%
#92530000000
0!
0%
#92535000000
1!
1%
#92540000000
0!
0%
#92545000000
1!
1%
#92550000000
0!
0%
#92555000000
1!
1%
#92560000000
0!
0%
#92565000000
1!
1%
#92570000000
0!
0%
#92575000000
1!
1%
#92580000000
0!
0%
#92585000000
1!
1%
#92590000000
0!
0%
#92595000000
1!
1%
#92600000000
0!
0%
#92605000000
1!
1%
#92610000000
0!
0%
#92615000000
1!
1%
#92620000000
0!
0%
#92625000000
1!
1%
#92630000000
0!
0%
#92635000000
1!
1%
#92640000000
0!
0%
#92645000000
1!
1%
#92650000000
0!
0%
#92655000000
1!
1%
#92660000000
0!
0%
#92665000000
1!
1%
#92670000000
0!
0%
#92675000000
1!
1%
#92680000000
0!
0%
#92685000000
1!
1%
#92690000000
0!
0%
#92695000000
1!
1%
#92700000000
0!
0%
#92705000000
1!
1%
#92710000000
0!
0%
#92715000000
1!
1%
#92720000000
0!
0%
#92725000000
1!
1%
#92730000000
0!
0%
#92735000000
1!
1%
#92740000000
0!
0%
#92745000000
1!
1%
#92750000000
0!
0%
#92755000000
1!
1%
#92760000000
0!
0%
#92765000000
1!
1%
#92770000000
0!
0%
#92775000000
1!
1%
#92780000000
0!
0%
#92785000000
1!
1%
#92790000000
0!
0%
#92795000000
1!
1%
#92800000000
0!
0%
#92805000000
1!
1%
#92810000000
0!
0%
#92815000000
1!
1%
#92820000000
0!
0%
#92825000000
1!
1%
#92830000000
0!
0%
#92835000000
1!
1%
#92840000000
0!
0%
#92845000000
1!
1%
#92850000000
0!
0%
#92855000000
1!
1%
#92860000000
0!
0%
#92865000000
1!
1%
#92870000000
0!
0%
#92875000000
1!
1%
#92880000000
0!
0%
#92885000000
1!
1%
#92890000000
0!
0%
#92895000000
1!
1%
#92900000000
0!
0%
#92905000000
1!
1%
#92910000000
0!
0%
#92915000000
1!
1%
#92920000000
0!
0%
#92925000000
1!
1%
#92930000000
0!
0%
#92935000000
1!
1%
#92940000000
0!
0%
#92945000000
1!
1%
#92950000000
0!
0%
#92955000000
1!
1%
#92960000000
0!
0%
#92965000000
1!
1%
#92970000000
0!
0%
#92975000000
1!
1%
#92980000000
0!
0%
#92985000000
1!
1%
#92990000000
0!
0%
#92995000000
1!
1%
#93000000000
0!
0%
#93005000000
1!
1%
#93010000000
0!
0%
#93015000000
1!
1%
#93020000000
0!
0%
#93025000000
1!
1%
#93030000000
0!
0%
#93035000000
1!
1%
#93040000000
0!
0%
#93045000000
1!
1%
#93050000000
0!
0%
#93055000000
1!
1%
#93060000000
0!
0%
#93065000000
1!
1%
#93070000000
0!
0%
#93075000000
1!
1%
#93080000000
0!
0%
#93085000000
1!
1%
#93090000000
0!
0%
#93095000000
1!
1%
#93100000000
0!
0%
#93105000000
1!
1%
#93110000000
0!
0%
#93115000000
1!
1%
#93120000000
0!
0%
#93125000000
1!
1%
#93130000000
0!
0%
#93135000000
1!
1%
#93140000000
0!
0%
#93145000000
1!
1%
#93150000000
0!
0%
#93155000000
1!
1%
#93160000000
0!
0%
#93165000000
1!
1%
#93170000000
0!
0%
#93175000000
1!
1%
#93180000000
0!
0%
#93185000000
1!
1%
#93190000000
0!
0%
#93195000000
1!
1%
#93200000000
0!
0%
#93205000000
1!
1%
#93210000000
0!
0%
#93215000000
1!
1%
#93220000000
0!
0%
#93225000000
1!
1%
#93230000000
0!
0%
#93235000000
1!
1%
#93240000000
0!
0%
#93245000000
1!
1%
#93250000000
0!
0%
#93255000000
1!
1%
#93260000000
0!
0%
#93265000000
1!
1%
#93270000000
0!
0%
#93275000000
1!
1%
#93280000000
0!
0%
#93285000000
1!
1%
#93290000000
0!
0%
#93295000000
1!
1%
#93300000000
0!
0%
#93305000000
1!
1%
#93310000000
0!
0%
#93315000000
1!
1%
#93320000000
0!
0%
#93325000000
1!
1%
#93330000000
0!
0%
#93335000000
1!
1%
#93340000000
0!
0%
#93345000000
1!
1%
#93350000000
0!
0%
#93355000000
1!
1%
#93360000000
0!
0%
#93365000000
1!
1%
#93370000000
0!
0%
#93375000000
1!
1%
#93380000000
0!
0%
#93385000000
1!
1%
#93390000000
0!
0%
#93395000000
1!
1%
#93400000000
0!
0%
#93405000000
1!
1%
#93410000000
0!
0%
#93415000000
1!
1%
#93420000000
0!
0%
#93425000000
1!
1%
#93430000000
0!
0%
#93435000000
1!
1%
#93440000000
0!
0%
#93445000000
1!
1%
#93450000000
0!
0%
#93455000000
1!
1%
#93460000000
0!
0%
#93465000000
1!
1%
#93470000000
0!
0%
#93475000000
1!
1%
#93480000000
0!
0%
#93485000000
1!
1%
#93490000000
0!
0%
#93495000000
1!
1%
#93500000000
0!
0%
#93505000000
1!
1%
#93510000000
0!
0%
#93515000000
1!
1%
#93520000000
0!
0%
#93525000000
1!
1%
#93530000000
0!
0%
#93535000000
1!
1%
#93540000000
0!
0%
#93545000000
1!
1%
#93550000000
0!
0%
#93555000000
1!
1%
#93560000000
0!
0%
#93565000000
1!
1%
#93570000000
0!
0%
#93575000000
1!
1%
#93580000000
0!
0%
#93585000000
1!
1%
#93590000000
0!
0%
#93595000000
1!
1%
#93600000000
0!
0%
#93605000000
1!
1%
#93610000000
0!
0%
#93615000000
1!
1%
#93620000000
0!
0%
#93625000000
1!
1%
#93630000000
0!
0%
#93635000000
1!
1%
#93640000000
0!
0%
#93645000000
1!
1%
#93650000000
0!
0%
#93655000000
1!
1%
#93660000000
0!
0%
#93665000000
1!
1%
#93670000000
0!
0%
#93675000000
1!
1%
#93680000000
0!
0%
#93685000000
1!
1%
#93690000000
0!
0%
#93695000000
1!
1%
#93700000000
0!
0%
#93705000000
1!
1%
#93710000000
0!
0%
#93715000000
1!
1%
#93720000000
0!
0%
#93725000000
1!
1%
#93730000000
0!
0%
#93735000000
1!
1%
#93740000000
0!
0%
#93745000000
1!
1%
#93750000000
0!
0%
#93755000000
1!
1%
#93760000000
0!
0%
#93765000000
1!
1%
#93770000000
0!
0%
#93775000000
1!
1%
#93780000000
0!
0%
#93785000000
1!
1%
#93790000000
0!
0%
#93795000000
1!
1%
#93800000000
0!
0%
#93805000000
1!
1%
#93810000000
0!
0%
#93815000000
1!
1%
#93820000000
0!
0%
#93825000000
1!
1%
#93830000000
0!
0%
#93835000000
1!
1%
#93840000000
0!
0%
#93845000000
1!
1%
#93850000000
0!
0%
#93855000000
1!
1%
#93860000000
0!
0%
#93865000000
1!
1%
#93870000000
0!
0%
#93875000000
1!
1%
#93880000000
0!
0%
#93885000000
1!
1%
#93890000000
0!
0%
#93895000000
1!
1%
#93900000000
0!
0%
#93905000000
1!
1%
#93910000000
0!
0%
#93915000000
1!
1%
#93920000000
0!
0%
#93925000000
1!
1%
#93930000000
0!
0%
#93935000000
1!
1%
#93940000000
0!
0%
#93945000000
1!
1%
#93950000000
0!
0%
#93955000000
1!
1%
#93960000000
0!
0%
#93965000000
1!
1%
#93970000000
0!
0%
#93975000000
1!
1%
#93980000000
0!
0%
#93985000000
1!
1%
#93990000000
0!
0%
#93995000000
1!
1%
#94000000000
0!
0%
#94005000000
1!
1%
#94010000000
0!
0%
#94015000000
1!
1%
#94020000000
0!
0%
#94025000000
1!
1%
#94030000000
0!
0%
#94035000000
1!
1%
#94040000000
0!
0%
#94045000000
1!
1%
#94050000000
0!
0%
#94055000000
1!
1%
#94060000000
0!
0%
#94065000000
1!
1%
#94070000000
0!
0%
#94075000000
1!
1%
#94080000000
0!
0%
#94085000000
1!
1%
#94090000000
0!
0%
#94095000000
1!
1%
#94100000000
0!
0%
#94105000000
1!
1%
#94110000000
0!
0%
#94115000000
1!
1%
#94120000000
0!
0%
#94125000000
1!
1%
#94130000000
0!
0%
#94135000000
1!
1%
#94140000000
0!
0%
#94145000000
1!
1%
#94150000000
0!
0%
#94155000000
1!
1%
#94160000000
0!
0%
#94165000000
1!
1%
#94170000000
0!
0%
#94175000000
1!
1%
#94180000000
0!
0%
#94185000000
1!
1%
#94190000000
0!
0%
#94195000000
1!
1%
#94200000000
0!
0%
#94205000000
1!
1%
#94210000000
0!
0%
#94215000000
1!
1%
#94220000000
0!
0%
#94225000000
1!
1%
#94230000000
0!
0%
#94235000000
1!
1%
#94240000000
0!
0%
#94245000000
1!
1%
#94250000000
0!
0%
#94255000000
1!
1%
#94260000000
0!
0%
#94265000000
1!
1%
#94270000000
0!
0%
#94275000000
1!
1%
#94280000000
0!
0%
#94285000000
1!
1%
#94290000000
0!
0%
#94295000000
1!
1%
#94300000000
0!
0%
#94305000000
1!
1%
#94310000000
0!
0%
#94315000000
1!
1%
#94320000000
0!
0%
#94325000000
1!
1%
#94330000000
0!
0%
#94335000000
1!
1%
#94340000000
0!
0%
#94345000000
1!
1%
#94350000000
0!
0%
#94355000000
1!
1%
#94360000000
0!
0%
#94365000000
1!
1%
#94370000000
0!
0%
#94375000000
1!
1%
#94380000000
0!
0%
#94385000000
1!
1%
#94390000000
0!
0%
#94395000000
1!
1%
#94400000000
0!
0%
#94405000000
1!
1%
#94410000000
0!
0%
#94415000000
1!
1%
#94420000000
0!
0%
#94425000000
1!
1%
#94430000000
0!
0%
#94435000000
1!
1%
#94440000000
0!
0%
#94445000000
1!
1%
#94450000000
0!
0%
#94455000000
1!
1%
#94460000000
0!
0%
#94465000000
1!
1%
#94470000000
0!
0%
#94475000000
1!
1%
#94480000000
0!
0%
#94485000000
1!
1%
#94490000000
0!
0%
#94495000000
1!
1%
#94500000000
0!
0%
#94505000000
1!
1%
#94510000000
0!
0%
#94515000000
1!
1%
#94520000000
0!
0%
#94525000000
1!
1%
#94530000000
0!
0%
#94535000000
1!
1%
#94540000000
0!
0%
#94545000000
1!
1%
#94550000000
0!
0%
#94555000000
1!
1%
#94560000000
0!
0%
#94565000000
1!
1%
#94570000000
0!
0%
#94575000000
1!
1%
#94580000000
0!
0%
#94585000000
1!
1%
#94590000000
0!
0%
#94595000000
1!
1%
#94600000000
0!
0%
#94605000000
1!
1%
#94610000000
0!
0%
#94615000000
1!
1%
#94620000000
0!
0%
#94625000000
1!
1%
#94630000000
0!
0%
#94635000000
1!
1%
#94640000000
0!
0%
#94645000000
1!
1%
#94650000000
0!
0%
#94655000000
1!
1%
#94660000000
0!
0%
#94665000000
1!
1%
#94670000000
0!
0%
#94675000000
1!
1%
#94680000000
0!
0%
#94685000000
1!
1%
#94690000000
0!
0%
#94695000000
1!
1%
#94700000000
0!
0%
#94705000000
1!
1%
#94710000000
0!
0%
#94715000000
1!
1%
#94720000000
0!
0%
#94725000000
1!
1%
#94730000000
0!
0%
#94735000000
1!
1%
#94740000000
0!
0%
#94745000000
1!
1%
#94750000000
0!
0%
#94755000000
1!
1%
#94760000000
0!
0%
#94765000000
1!
1%
#94770000000
0!
0%
#94775000000
1!
1%
#94780000000
0!
0%
#94785000000
1!
1%
#94790000000
0!
0%
#94795000000
1!
1%
#94800000000
0!
0%
#94805000000
1!
1%
#94810000000
0!
0%
#94815000000
1!
1%
#94820000000
0!
0%
#94825000000
1!
1%
#94830000000
0!
0%
#94835000000
1!
1%
#94840000000
0!
0%
#94845000000
1!
1%
#94850000000
0!
0%
#94855000000
1!
1%
#94860000000
0!
0%
#94865000000
1!
1%
#94870000000
0!
0%
#94875000000
1!
1%
#94880000000
0!
0%
#94885000000
1!
1%
#94890000000
0!
0%
#94895000000
1!
1%
#94900000000
0!
0%
#94905000000
1!
1%
#94910000000
0!
0%
#94915000000
1!
1%
#94920000000
0!
0%
#94925000000
1!
1%
#94930000000
0!
0%
#94935000000
1!
1%
#94940000000
0!
0%
#94945000000
1!
1%
#94950000000
0!
0%
#94955000000
1!
1%
#94960000000
0!
0%
#94965000000
1!
1%
#94970000000
0!
0%
#94975000000
1!
1%
#94980000000
0!
0%
#94985000000
1!
1%
#94990000000
0!
0%
#94995000000
1!
1%
#95000000000
0!
0%
#95005000000
1!
1%
#95010000000
0!
0%
#95015000000
1!
1%
#95020000000
0!
0%
#95025000000
1!
1%
#95030000000
0!
0%
#95035000000
1!
1%
#95040000000
0!
0%
#95045000000
1!
1%
#95050000000
0!
0%
#95055000000
1!
1%
#95060000000
0!
0%
#95065000000
1!
1%
#95070000000
0!
0%
#95075000000
1!
1%
#95080000000
0!
0%
#95085000000
1!
1%
#95090000000
0!
0%
#95095000000
1!
1%
#95100000000
0!
0%
#95105000000
1!
1%
#95110000000
0!
0%
#95115000000
1!
1%
#95120000000
0!
0%
#95125000000
1!
1%
#95130000000
0!
0%
#95135000000
1!
1%
#95140000000
0!
0%
#95145000000
1!
1%
#95150000000
0!
0%
#95155000000
1!
1%
#95160000000
0!
0%
#95165000000
1!
1%
#95170000000
0!
0%
#95175000000
1!
1%
#95180000000
0!
0%
#95185000000
1!
1%
#95190000000
0!
0%
#95195000000
1!
1%
#95200000000
0!
0%
#95205000000
1!
1%
#95210000000
0!
0%
#95215000000
1!
1%
#95220000000
0!
0%
#95225000000
1!
1%
#95230000000
0!
0%
#95235000000
1!
1%
#95240000000
0!
0%
#95245000000
1!
1%
#95250000000
0!
0%
#95255000000
1!
1%
#95260000000
0!
0%
#95265000000
1!
1%
#95270000000
0!
0%
#95275000000
1!
1%
#95280000000
0!
0%
#95285000000
1!
1%
#95290000000
0!
0%
#95295000000
1!
1%
#95300000000
0!
0%
#95305000000
1!
1%
#95310000000
0!
0%
#95315000000
1!
1%
#95320000000
0!
0%
#95325000000
1!
1%
#95330000000
0!
0%
#95335000000
1!
1%
#95340000000
0!
0%
#95345000000
1!
1%
#95350000000
0!
0%
#95355000000
1!
1%
#95360000000
0!
0%
#95365000000
1!
1%
#95370000000
0!
0%
#95375000000
1!
1%
#95380000000
0!
0%
#95385000000
1!
1%
#95390000000
0!
0%
#95395000000
1!
1%
#95400000000
0!
0%
#95405000000
1!
1%
#95410000000
0!
0%
#95415000000
1!
1%
#95420000000
0!
0%
#95425000000
1!
1%
#95430000000
0!
0%
#95435000000
1!
1%
#95440000000
0!
0%
#95445000000
1!
1%
#95450000000
0!
0%
#95455000000
1!
1%
#95460000000
0!
0%
#95465000000
1!
1%
#95470000000
0!
0%
#95475000000
1!
1%
#95480000000
0!
0%
#95485000000
1!
1%
#95490000000
0!
0%
#95495000000
1!
1%
#95500000000
0!
0%
#95505000000
1!
1%
#95510000000
0!
0%
#95515000000
1!
1%
#95520000000
0!
0%
#95525000000
1!
1%
#95530000000
0!
0%
#95535000000
1!
1%
#95540000000
0!
0%
#95545000000
1!
1%
#95550000000
0!
0%
#95555000000
1!
1%
#95560000000
0!
0%
#95565000000
1!
1%
#95570000000
0!
0%
#95575000000
1!
1%
#95580000000
0!
0%
#95585000000
1!
1%
#95590000000
0!
0%
#95595000000
1!
1%
#95600000000
0!
0%
#95605000000
1!
1%
#95610000000
0!
0%
#95615000000
1!
1%
#95620000000
0!
0%
#95625000000
1!
1%
#95630000000
0!
0%
#95635000000
1!
1%
#95640000000
0!
0%
#95645000000
1!
1%
#95650000000
0!
0%
#95655000000
1!
1%
#95660000000
0!
0%
#95665000000
1!
1%
#95670000000
0!
0%
#95675000000
1!
1%
#95680000000
0!
0%
#95685000000
1!
1%
#95690000000
0!
0%
#95695000000
1!
1%
#95700000000
0!
0%
#95705000000
1!
1%
#95710000000
0!
0%
#95715000000
1!
1%
#95720000000
0!
0%
#95725000000
1!
1%
#95730000000
0!
0%
#95735000000
1!
1%
#95740000000
0!
0%
#95745000000
1!
1%
#95750000000
0!
0%
#95755000000
1!
1%
#95760000000
0!
0%
#95765000000
1!
1%
#95770000000
0!
0%
#95775000000
1!
1%
#95780000000
0!
0%
#95785000000
1!
1%
#95790000000
0!
0%
#95795000000
1!
1%
#95800000000
0!
0%
#95805000000
1!
1%
#95810000000
0!
0%
#95815000000
1!
1%
#95820000000
0!
0%
#95825000000
1!
1%
#95830000000
0!
0%
#95835000000
1!
1%
#95840000000
0!
0%
#95845000000
1!
1%
#95850000000
0!
0%
#95855000000
1!
1%
#95860000000
0!
0%
#95865000000
1!
1%
#95870000000
0!
0%
#95875000000
1!
1%
#95880000000
0!
0%
#95885000000
1!
1%
#95890000000
0!
0%
#95895000000
1!
1%
#95900000000
0!
0%
#95905000000
1!
1%
#95910000000
0!
0%
#95915000000
1!
1%
#95920000000
0!
0%
#95925000000
1!
1%
#95930000000
0!
0%
#95935000000
1!
1%
#95940000000
0!
0%
#95945000000
1!
1%
#95950000000
0!
0%
#95955000000
1!
1%
#95960000000
0!
0%
#95965000000
1!
1%
#95970000000
0!
0%
#95975000000
1!
1%
#95980000000
0!
0%
#95985000000
1!
1%
#95990000000
0!
0%
#95995000000
1!
1%
#96000000000
0!
0%
#96005000000
1!
1%
#96010000000
0!
0%
#96015000000
1!
1%
#96020000000
0!
0%
#96025000000
1!
1%
#96030000000
0!
0%
#96035000000
1!
1%
#96040000000
0!
0%
#96045000000
1!
1%
#96050000000
0!
0%
#96055000000
1!
1%
#96060000000
0!
0%
#96065000000
1!
1%
#96070000000
0!
0%
#96075000000
1!
1%
#96080000000
0!
0%
#96085000000
1!
1%
#96090000000
0!
0%
#96095000000
1!
1%
#96100000000
0!
0%
#96105000000
1!
1%
#96110000000
0!
0%
#96115000000
1!
1%
#96120000000
0!
0%
#96125000000
1!
1%
#96130000000
0!
0%
#96135000000
1!
1%
#96140000000
0!
0%
#96145000000
1!
1%
#96150000000
0!
0%
#96155000000
1!
1%
#96160000000
0!
0%
#96165000000
1!
1%
#96170000000
0!
0%
#96175000000
1!
1%
#96180000000
0!
0%
#96185000000
1!
1%
#96190000000
0!
0%
#96195000000
1!
1%
#96200000000
0!
0%
#96205000000
1!
1%
#96210000000
0!
0%
#96215000000
1!
1%
#96220000000
0!
0%
#96225000000
1!
1%
#96230000000
0!
0%
#96235000000
1!
1%
#96240000000
0!
0%
#96245000000
1!
1%
#96250000000
0!
0%
#96255000000
1!
1%
#96260000000
0!
0%
#96265000000
1!
1%
#96270000000
0!
0%
#96275000000
1!
1%
#96280000000
0!
0%
#96285000000
1!
1%
#96290000000
0!
0%
#96295000000
1!
1%
#96300000000
0!
0%
#96305000000
1!
1%
#96310000000
0!
0%
#96315000000
1!
1%
#96320000000
0!
0%
#96325000000
1!
1%
#96330000000
0!
0%
#96335000000
1!
1%
#96340000000
0!
0%
#96345000000
1!
1%
#96350000000
0!
0%
#96355000000
1!
1%
#96360000000
0!
0%
#96365000000
1!
1%
#96370000000
0!
0%
#96375000000
1!
1%
#96380000000
0!
0%
#96385000000
1!
1%
#96390000000
0!
0%
#96395000000
1!
1%
#96400000000
0!
0%
#96405000000
1!
1%
#96410000000
0!
0%
#96415000000
1!
1%
#96420000000
0!
0%
#96425000000
1!
1%
#96430000000
0!
0%
#96435000000
1!
1%
#96440000000
0!
0%
#96445000000
1!
1%
#96450000000
0!
0%
#96455000000
1!
1%
#96460000000
0!
0%
#96465000000
1!
1%
#96470000000
0!
0%
#96475000000
1!
1%
#96480000000
0!
0%
#96485000000
1!
1%
#96490000000
0!
0%
#96495000000
1!
1%
#96500000000
0!
0%
#96505000000
1!
1%
#96510000000
0!
0%
#96515000000
1!
1%
#96520000000
0!
0%
#96525000000
1!
1%
#96530000000
0!
0%
#96535000000
1!
1%
#96540000000
0!
0%
#96545000000
1!
1%
#96550000000
0!
0%
#96555000000
1!
1%
#96560000000
0!
0%
#96565000000
1!
1%
#96570000000
0!
0%
#96575000000
1!
1%
#96580000000
0!
0%
#96585000000
1!
1%
#96590000000
0!
0%
#96595000000
1!
1%
#96600000000
0!
0%
#96605000000
1!
1%
#96610000000
0!
0%
#96615000000
1!
1%
#96620000000
0!
0%
#96625000000
1!
1%
#96630000000
0!
0%
#96635000000
1!
1%
#96640000000
0!
0%
#96645000000
1!
1%
#96650000000
0!
0%
#96655000000
1!
1%
#96660000000
0!
0%
#96665000000
1!
1%
#96670000000
0!
0%
#96675000000
1!
1%
#96680000000
0!
0%
#96685000000
1!
1%
#96690000000
0!
0%
#96695000000
1!
1%
#96700000000
0!
0%
#96705000000
1!
1%
#96710000000
0!
0%
#96715000000
1!
1%
#96720000000
0!
0%
#96725000000
1!
1%
#96730000000
0!
0%
#96735000000
1!
1%
#96740000000
0!
0%
#96745000000
1!
1%
#96750000000
0!
0%
#96755000000
1!
1%
#96760000000
0!
0%
#96765000000
1!
1%
#96770000000
0!
0%
#96775000000
1!
1%
#96780000000
0!
0%
#96785000000
1!
1%
#96790000000
0!
0%
#96795000000
1!
1%
#96800000000
0!
0%
#96805000000
1!
1%
#96810000000
0!
0%
#96815000000
1!
1%
#96820000000
0!
0%
#96825000000
1!
1%
#96830000000
0!
0%
#96835000000
1!
1%
#96840000000
0!
0%
#96845000000
1!
1%
#96850000000
0!
0%
#96855000000
1!
1%
#96860000000
0!
0%
#96865000000
1!
1%
#96870000000
0!
0%
#96875000000
1!
1%
#96880000000
0!
0%
#96885000000
1!
1%
#96890000000
0!
0%
#96895000000
1!
1%
#96900000000
0!
0%
#96905000000
1!
1%
#96910000000
0!
0%
#96915000000
1!
1%
#96920000000
0!
0%
#96925000000
1!
1%
#96930000000
0!
0%
#96935000000
1!
1%
#96940000000
0!
0%
#96945000000
1!
1%
#96950000000
0!
0%
#96955000000
1!
1%
#96960000000
0!
0%
#96965000000
1!
1%
#96970000000
0!
0%
#96975000000
1!
1%
#96980000000
0!
0%
#96985000000
1!
1%
#96990000000
0!
0%
#96995000000
1!
1%
#97000000000
0!
0%
#97005000000
1!
1%
#97010000000
0!
0%
#97015000000
1!
1%
#97020000000
0!
0%
#97025000000
1!
1%
#97030000000
0!
0%
#97035000000
1!
1%
#97040000000
0!
0%
#97045000000
1!
1%
#97050000000
0!
0%
#97055000000
1!
1%
#97060000000
0!
0%
#97065000000
1!
1%
#97070000000
0!
0%
#97075000000
1!
1%
#97080000000
0!
0%
#97085000000
1!
1%
#97090000000
0!
0%
#97095000000
1!
1%
#97100000000
0!
0%
#97105000000
1!
1%
#97110000000
0!
0%
#97115000000
1!
1%
#97120000000
0!
0%
#97125000000
1!
1%
#97130000000
0!
0%
#97135000000
1!
1%
#97140000000
0!
0%
#97145000000
1!
1%
#97150000000
0!
0%
#97155000000
1!
1%
#97160000000
0!
0%
#97165000000
1!
1%
#97170000000
0!
0%
#97175000000
1!
1%
#97180000000
0!
0%
#97185000000
1!
1%
#97190000000
0!
0%
#97195000000
1!
1%
#97200000000
0!
0%
#97205000000
1!
1%
#97210000000
0!
0%
#97215000000
1!
1%
#97220000000
0!
0%
#97225000000
1!
1%
#97230000000
0!
0%
#97235000000
1!
1%
#97240000000
0!
0%
#97245000000
1!
1%
#97250000000
0!
0%
#97255000000
1!
1%
#97260000000
0!
0%
#97265000000
1!
1%
#97270000000
0!
0%
#97275000000
1!
1%
#97280000000
0!
0%
#97285000000
1!
1%
#97290000000
0!
0%
#97295000000
1!
1%
#97300000000
0!
0%
#97305000000
1!
1%
#97310000000
0!
0%
#97315000000
1!
1%
#97320000000
0!
0%
#97325000000
1!
1%
#97330000000
0!
0%
#97335000000
1!
1%
#97340000000
0!
0%
#97345000000
1!
1%
#97350000000
0!
0%
#97355000000
1!
1%
#97360000000
0!
0%
#97365000000
1!
1%
#97370000000
0!
0%
#97375000000
1!
1%
#97380000000
0!
0%
#97385000000
1!
1%
#97390000000
0!
0%
#97395000000
1!
1%
#97400000000
0!
0%
#97405000000
1!
1%
#97410000000
0!
0%
#97415000000
1!
1%
#97420000000
0!
0%
#97425000000
1!
1%
#97430000000
0!
0%
#97435000000
1!
1%
#97440000000
0!
0%
#97445000000
1!
1%
#97450000000
0!
0%
#97455000000
1!
1%
#97460000000
0!
0%
#97465000000
1!
1%
#97470000000
0!
0%
#97475000000
1!
1%
#97480000000
0!
0%
#97485000000
1!
1%
#97490000000
0!
0%
#97495000000
1!
1%
#97500000000
0!
0%
#97505000000
1!
1%
#97510000000
0!
0%
#97515000000
1!
1%
#97520000000
0!
0%
#97525000000
1!
1%
#97530000000
0!
0%
#97535000000
1!
1%
#97540000000
0!
0%
#97545000000
1!
1%
#97550000000
0!
0%
#97555000000
1!
1%
#97560000000
0!
0%
#97565000000
1!
1%
#97570000000
0!
0%
#97575000000
1!
1%
#97580000000
0!
0%
#97585000000
1!
1%
#97590000000
0!
0%
#97595000000
1!
1%
#97600000000
0!
0%
#97605000000
1!
1%
#97610000000
0!
0%
#97615000000
1!
1%
#97620000000
0!
0%
#97625000000
1!
1%
#97630000000
0!
0%
#97635000000
1!
1%
#97640000000
0!
0%
#97645000000
1!
1%
#97650000000
0!
0%
#97655000000
1!
1%
#97660000000
0!
0%
#97665000000
1!
1%
#97670000000
0!
0%
#97675000000
1!
1%
#97680000000
0!
0%
#97685000000
1!
1%
#97690000000
0!
0%
#97695000000
1!
1%
#97700000000
0!
0%
#97705000000
1!
1%
#97710000000
0!
0%
#97715000000
1!
1%
#97720000000
0!
0%
#97725000000
1!
1%
#97730000000
0!
0%
#97735000000
1!
1%
#97740000000
0!
0%
#97745000000
1!
1%
#97750000000
0!
0%
#97755000000
1!
1%
#97760000000
0!
0%
#97765000000
1!
1%
#97770000000
0!
0%
#97775000000
1!
1%
#97780000000
0!
0%
#97785000000
1!
1%
#97790000000
0!
0%
#97795000000
1!
1%
#97800000000
0!
0%
#97805000000
1!
1%
#97810000000
0!
0%
#97815000000
1!
1%
#97820000000
0!
0%
#97825000000
1!
1%
#97830000000
0!
0%
#97835000000
1!
1%
#97840000000
0!
0%
#97845000000
1!
1%
#97850000000
0!
0%
#97855000000
1!
1%
#97860000000
0!
0%
#97865000000
1!
1%
#97870000000
0!
0%
#97875000000
1!
1%
#97880000000
0!
0%
#97885000000
1!
1%
#97890000000
0!
0%
#97895000000
1!
1%
#97900000000
0!
0%
#97905000000
1!
1%
#97910000000
0!
0%
#97915000000
1!
1%
#97920000000
0!
0%
#97925000000
1!
1%
#97930000000
0!
0%
#97935000000
1!
1%
#97940000000
0!
0%
#97945000000
1!
1%
#97950000000
0!
0%
#97955000000
1!
1%
#97960000000
0!
0%
#97965000000
1!
1%
#97970000000
0!
0%
#97975000000
1!
1%
#97980000000
0!
0%
#97985000000
1!
1%
#97990000000
0!
0%
#97995000000
1!
1%
#98000000000
0!
0%
#98005000000
1!
1%
#98010000000
0!
0%
#98015000000
1!
1%
#98020000000
0!
0%
#98025000000
1!
1%
#98030000000
0!
0%
#98035000000
1!
1%
#98040000000
0!
0%
#98045000000
1!
1%
#98050000000
0!
0%
#98055000000
1!
1%
#98060000000
0!
0%
#98065000000
1!
1%
#98070000000
0!
0%
#98075000000
1!
1%
#98080000000
0!
0%
#98085000000
1!
1%
#98090000000
0!
0%
#98095000000
1!
1%
#98100000000
0!
0%
#98105000000
1!
1%
#98110000000
0!
0%
#98115000000
1!
1%
#98120000000
0!
0%
#98125000000
1!
1%
#98130000000
0!
0%
#98135000000
1!
1%
#98140000000
0!
0%
#98145000000
1!
1%
#98150000000
0!
0%
#98155000000
1!
1%
#98160000000
0!
0%
#98165000000
1!
1%
#98170000000
0!
0%
#98175000000
1!
1%
#98180000000
0!
0%
#98185000000
1!
1%
#98190000000
0!
0%
#98195000000
1!
1%
#98200000000
0!
0%
#98205000000
1!
1%
#98210000000
0!
0%
#98215000000
1!
1%
#98220000000
0!
0%
#98225000000
1!
1%
#98230000000
0!
0%
#98235000000
1!
1%
#98240000000
0!
0%
#98245000000
1!
1%
#98250000000
0!
0%
#98255000000
1!
1%
#98260000000
0!
0%
#98265000000
1!
1%
#98270000000
0!
0%
#98275000000
1!
1%
#98280000000
0!
0%
#98285000000
1!
1%
#98290000000
0!
0%
#98295000000
1!
1%
#98300000000
0!
0%
#98305000000
1!
1%
#98310000000
0!
0%
#98315000000
1!
1%
#98320000000
0!
0%
#98325000000
1!
1%
#98330000000
0!
0%
#98335000000
1!
1%
#98340000000
0!
0%
#98345000000
1!
1%
#98350000000
0!
0%
#98355000000
1!
1%
#98360000000
0!
0%
#98365000000
1!
1%
#98370000000
0!
0%
#98375000000
1!
1%
#98380000000
0!
0%
#98385000000
1!
1%
#98390000000
0!
0%
#98395000000
1!
1%
#98400000000
0!
0%
#98405000000
1!
1%
#98410000000
0!
0%
#98415000000
1!
1%
#98420000000
0!
0%
#98425000000
1!
1%
#98430000000
0!
0%
#98435000000
1!
1%
#98440000000
0!
0%
#98445000000
1!
1%
#98450000000
0!
0%
#98455000000
1!
1%
#98460000000
0!
0%
#98465000000
1!
1%
#98470000000
0!
0%
#98475000000
1!
1%
#98480000000
0!
0%
#98485000000
1!
1%
#98490000000
0!
0%
#98495000000
1!
1%
#98500000000
0!
0%
#98505000000
1!
1%
#98510000000
0!
0%
#98515000000
1!
1%
#98520000000
0!
0%
#98525000000
1!
1%
#98530000000
0!
0%
#98535000000
1!
1%
#98540000000
0!
0%
#98545000000
1!
1%
#98550000000
0!
0%
#98555000000
1!
1%
#98560000000
0!
0%
#98565000000
1!
1%
#98570000000
0!
0%
#98575000000
1!
1%
#98580000000
0!
0%
#98585000000
1!
1%
#98590000000
0!
0%
#98595000000
1!
1%
#98600000000
0!
0%
#98605000000
1!
1%
#98610000000
0!
0%
#98615000000
1!
1%
#98620000000
0!
0%
#98625000000
1!
1%
#98630000000
0!
0%
#98635000000
1!
1%
#98640000000
0!
0%
#98645000000
1!
1%
#98650000000
0!
0%
#98655000000
1!
1%
#98660000000
0!
0%
#98665000000
1!
1%
#98670000000
0!
0%
#98675000000
1!
1%
#98680000000
0!
0%
#98685000000
1!
1%
#98690000000
0!
0%
#98695000000
1!
1%
#98700000000
0!
0%
#98705000000
1!
1%
#98710000000
0!
0%
#98715000000
1!
1%
#98720000000
0!
0%
#98725000000
1!
1%
#98730000000
0!
0%
#98735000000
1!
1%
#98740000000
0!
0%
#98745000000
1!
1%
#98750000000
0!
0%
#98755000000
1!
1%
#98760000000
0!
0%
#98765000000
1!
1%
#98770000000
0!
0%
#98775000000
1!
1%
#98780000000
0!
0%
#98785000000
1!
1%
#98790000000
0!
0%
#98795000000
1!
1%
#98800000000
0!
0%
#98805000000
1!
1%
#98810000000
0!
0%
#98815000000
1!
1%
#98820000000
0!
0%
#98825000000
1!
1%
#98830000000
0!
0%
#98835000000
1!
1%
#98840000000
0!
0%
#98845000000
1!
1%
#98850000000
0!
0%
#98855000000
1!
1%
#98860000000
0!
0%
#98865000000
1!
1%
#98870000000
0!
0%
#98875000000
1!
1%
#98880000000
0!
0%
#98885000000
1!
1%
#98890000000
0!
0%
#98895000000
1!
1%
#98900000000
0!
0%
#98905000000
1!
1%
#98910000000
0!
0%
#98915000000
1!
1%
#98920000000
0!
0%
#98925000000
1!
1%
#98930000000
0!
0%
#98935000000
1!
1%
#98940000000
0!
0%
#98945000000
1!
1%
#98950000000
0!
0%
#98955000000
1!
1%
#98960000000
0!
0%
#98965000000
1!
1%
#98970000000
0!
0%
#98975000000
1!
1%
#98980000000
0!
0%
#98985000000
1!
1%
#98990000000
0!
0%
#98995000000
1!
1%
#99000000000
0!
0%
#99005000000
1!
1%
#99010000000
0!
0%
#99015000000
1!
1%
#99020000000
0!
0%
#99025000000
1!
1%
#99030000000
0!
0%
#99035000000
1!
1%
#99040000000
0!
0%
#99045000000
1!
1%
#99050000000
0!
0%
#99055000000
1!
1%
#99060000000
0!
0%
#99065000000
1!
1%
#99070000000
0!
0%
#99075000000
1!
1%
#99080000000
0!
0%
#99085000000
1!
1%
#99090000000
0!
0%
#99095000000
1!
1%
#99100000000
0!
0%
#99105000000
1!
1%
#99110000000
0!
0%
#99115000000
1!
1%
#99120000000
0!
0%
#99125000000
1!
1%
#99130000000
0!
0%
#99135000000
1!
1%
#99140000000
0!
0%
#99145000000
1!
1%
#99150000000
0!
0%
#99155000000
1!
1%
#99160000000
0!
0%
#99165000000
1!
1%
#99170000000
0!
0%
#99175000000
1!
1%
#99180000000
0!
0%
#99185000000
1!
1%
#99190000000
0!
0%
#99195000000
1!
1%
#99200000000
0!
0%
#99205000000
1!
1%
#99210000000
0!
0%
#99215000000
1!
1%
#99220000000
0!
0%
#99225000000
1!
1%
#99230000000
0!
0%
#99235000000
1!
1%
#99240000000
0!
0%
#99245000000
1!
1%
#99250000000
0!
0%
#99255000000
1!
1%
#99260000000
0!
0%
#99265000000
1!
1%
#99270000000
0!
0%
#99275000000
1!
1%
#99280000000
0!
0%
#99285000000
1!
1%
#99290000000
0!
0%
#99295000000
1!
1%
#99300000000
0!
0%
#99305000000
1!
1%
#99310000000
0!
0%
#99315000000
1!
1%
#99320000000
0!
0%
#99325000000
1!
1%
#99330000000
0!
0%
#99335000000
1!
1%
#99340000000
0!
0%
#99345000000
1!
1%
#99350000000
0!
0%
#99355000000
1!
1%
#99360000000
0!
0%
#99365000000
1!
1%
#99370000000
0!
0%
#99375000000
1!
1%
#99380000000
0!
0%
#99385000000
1!
1%
#99390000000
0!
0%
#99395000000
1!
1%
#99400000000
0!
0%
#99405000000
1!
1%
#99410000000
0!
0%
#99415000000
1!
1%
#99420000000
0!
0%
#99425000000
1!
1%
#99430000000
0!
0%
#99435000000
1!
1%
#99440000000
0!
0%
#99445000000
1!
1%
#99450000000
0!
0%
#99455000000
1!
1%
#99460000000
0!
0%
#99465000000
1!
1%
#99470000000
0!
0%
#99475000000
1!
1%
#99480000000
0!
0%
#99485000000
1!
1%
#99490000000
0!
0%
#99495000000
1!
1%
#99500000000
0!
0%
#99505000000
1!
1%
#99510000000
0!
0%
#99515000000
1!
1%
#99520000000
0!
0%
#99525000000
1!
1%
#99530000000
0!
0%
#99535000000
1!
1%
#99540000000
0!
0%
#99545000000
1!
1%
#99550000000
0!
0%
#99555000000
1!
1%
#99560000000
0!
0%
#99565000000
1!
1%
#99570000000
0!
0%
#99575000000
1!
1%
#99580000000
0!
0%
#99585000000
1!
1%
#99590000000
0!
0%
#99595000000
1!
1%
#99600000000
0!
0%
#99605000000
1!
1%
#99610000000
0!
0%
#99615000000
1!
1%
#99620000000
0!
0%
#99625000000
1!
1%
#99630000000
0!
0%
#99635000000
1!
1%
#99640000000
0!
0%
#99645000000
1!
1%
#99650000000
0!
0%
#99655000000
1!
1%
#99660000000
0!
0%
#99665000000
1!
1%
#99670000000
0!
0%
#99675000000
1!
1%
#99680000000
0!
0%
#99685000000
1!
1%
#99690000000
0!
0%
#99695000000
1!
1%
#99700000000
0!
0%
#99705000000
1!
1%
#99710000000
0!
0%
#99715000000
1!
1%
#99720000000
0!
0%
#99725000000
1!
1%
#99730000000
0!
0%
#99735000000
1!
1%
#99740000000
0!
0%
#99745000000
1!
1%
#99750000000
0!
0%
#99755000000
1!
1%
#99760000000
0!
0%
#99765000000
1!
1%
#99770000000
0!
0%
#99775000000
1!
1%
#99780000000
0!
0%
#99785000000
1!
1%
#99790000000
0!
0%
#99795000000
1!
1%
#99800000000
0!
0%
#99805000000
1!
1%
#99810000000
0!
0%
#99815000000
1!
1%
#99820000000
0!
0%
#99825000000
1!
1%
#99830000000
0!
0%
#99835000000
1!
1%
#99840000000
0!
0%
#99845000000
1!
1%
#99850000000
0!
0%
#99855000000
1!
1%
#99860000000
0!
0%
#99865000000
1!
1%
#99870000000
0!
0%
#99875000000
1!
1%
#99880000000
0!
0%
#99885000000
1!
1%
#99890000000
0!
0%
#99895000000
1!
1%
#99900000000
0!
0%
#99905000000
1!
1%
#99910000000
0!
0%
#99915000000
1!
1%
#99920000000
0!
0%
#99925000000
1!
1%
#99930000000
0!
0%
#99935000000
1!
1%
#99940000000
0!
0%
#99945000000
1!
1%
#99950000000
0!
0%
#99955000000
1!
1%
#99960000000
0!
0%
#99965000000
1!
1%
#99970000000
0!
0%
#99975000000
1!
1%
#99980000000
0!
0%
#99985000000
1!
1%
#99990000000
0!
0%
#99995000000
1!
1%
#100000000000
0!
0%
#100005000000
1!
1%
#100010000000
0!
0%
#100015000000
1!
1%
#100020000000
0!
0%
#100025000000
1!
1%
#100030000000
0!
0%
#100035000000
1!
1%
#100040000000
0!
0%
#100045000000
1!
1%
#100050000000
0!
0%
#100055000000
1!
1%
#100060000000
0!
0%
#100065000000
1!
1%
#100070000000
0!
0%
#100075000000
1!
1%
#100080000000
0!
0%
#100085000000
1!
1%
#100090000000
0!
0%
#100095000000
1!
1%
#100100000000
0!
0%
#100105000000
1!
1%
#100110000000
0!
0%
#100115000000
1!
1%
#100120000000
0!
0%
#100125000000
1!
1%
#100130000000
0!
0%
#100135000000
1!
1%
#100140000000
0!
0%
#100145000000
1!
1%
#100150000000
0!
0%
#100155000000
1!
1%
#100160000000
0!
0%
#100165000000
1!
1%
#100170000000
0!
0%
#100175000000
1!
1%
#100180000000
0!
0%
#100185000000
1!
1%
#100190000000
0!
0%
#100195000000
1!
1%
#100200000000
0!
0%
#100205000000
1!
1%
#100210000000
0!
0%
#100215000000
1!
1%
#100220000000
0!
0%
#100225000000
1!
1%
#100230000000
0!
0%
#100235000000
1!
1%
#100240000000
0!
0%
#100245000000
1!
1%
#100250000000
0!
0%
#100255000000
1!
1%
#100260000000
0!
0%
#100265000000
1!
1%
#100270000000
0!
0%
#100275000000
1!
1%
#100280000000
0!
0%
#100285000000
1!
1%
#100290000000
0!
0%
#100295000000
1!
1%
#100300000000
0!
0%
#100305000000
1!
1%
#100310000000
0!
0%
#100315000000
1!
1%
#100320000000
0!
0%
#100325000000
1!
1%
#100330000000
0!
0%
#100335000000
1!
1%
#100340000000
0!
0%
#100345000000
1!
1%
#100350000000
0!
0%
#100355000000
1!
1%
#100360000000
0!
0%
#100365000000
1!
1%
#100370000000
0!
0%
#100375000000
1!
1%
#100380000000
0!
0%
#100385000000
1!
1%
#100390000000
0!
0%
#100395000000
1!
1%
#100400000000
0!
0%
#100405000000
1!
1%
#100410000000
0!
0%
#100415000000
1!
1%
#100420000000
0!
0%
#100425000000
1!
1%
#100430000000
0!
0%
#100435000000
1!
1%
#100440000000
0!
0%
#100445000000
1!
1%
#100450000000
0!
0%
#100455000000
1!
1%
#100460000000
0!
0%
#100465000000
1!
1%
#100470000000
0!
0%
#100475000000
1!
1%
#100480000000
0!
0%
#100485000000
1!
1%
#100490000000
0!
0%
#100495000000
1!
1%
#100500000000
0!
0%
#100505000000
1!
1%
#100510000000
0!
0%
#100515000000
1!
1%
#100520000000
0!
0%
#100525000000
1!
1%
#100530000000
0!
0%
#100535000000
1!
1%
#100540000000
0!
0%
#100545000000
1!
1%
#100550000000
0!
0%
#100555000000
1!
1%
#100560000000
0!
0%
#100565000000
1!
1%
#100570000000
0!
0%
#100575000000
1!
1%
#100580000000
0!
0%
#100585000000
1!
1%
#100590000000
0!
0%
#100595000000
1!
1%
#100600000000
0!
0%
#100605000000
1!
1%
#100610000000
0!
0%
#100615000000
1!
1%
#100620000000
0!
0%
#100625000000
1!
1%
#100630000000
0!
0%
#100635000000
1!
1%
#100640000000
0!
0%
#100645000000
1!
1%
#100650000000
0!
0%
#100655000000
1!
1%
#100660000000
0!
0%
#100665000000
1!
1%
#100670000000
0!
0%
#100675000000
1!
1%
#100680000000
0!
0%
#100685000000
1!
1%
#100690000000
0!
0%
#100695000000
1!
1%
#100700000000
0!
0%
#100705000000
1!
1%
#100710000000
0!
0%
#100715000000
1!
1%
#100720000000
0!
0%
#100725000000
1!
1%
#100730000000
0!
0%
#100735000000
1!
1%
#100740000000
0!
0%
#100745000000
1!
1%
#100750000000
0!
0%
#100755000000
1!
1%
#100760000000
0!
0%
#100765000000
1!
1%
#100770000000
0!
0%
#100775000000
1!
1%
#100780000000
0!
0%
#100785000000
1!
1%
#100790000000
0!
0%
#100795000000
1!
1%
#100800000000
0!
0%
#100805000000
1!
1%
#100810000000
0!
0%
#100815000000
1!
1%
#100820000000
0!
0%
#100825000000
1!
1%
#100830000000
0!
0%
#100835000000
1!
1%
#100840000000
0!
0%
#100845000000
1!
1%
#100850000000
0!
0%
#100855000000
1!
1%
#100860000000
0!
0%
#100865000000
1!
1%
#100870000000
0!
0%
#100875000000
1!
1%
#100880000000
0!
0%
#100885000000
1!
1%
#100890000000
0!
0%
#100895000000
1!
1%
#100900000000
0!
0%
#100905000000
1!
1%
#100910000000
0!
0%
#100915000000
1!
1%
#100920000000
0!
0%
#100925000000
1!
1%
#100930000000
0!
0%
#100935000000
1!
1%
#100940000000
0!
0%
#100945000000
1!
1%
#100950000000
0!
0%
#100955000000
1!
1%
#100960000000
0!
0%
#100965000000
1!
1%
#100970000000
0!
0%
#100975000000
1!
1%
#100980000000
0!
0%
#100985000000
1!
1%
#100990000000
0!
0%
#100995000000
1!
1%
#101000000000
0!
0%
#101005000000
1!
1%
#101010000000
0!
0%
#101015000000
1!
1%
#101020000000
0!
0%
#101025000000
1!
1%
#101030000000
0!
0%
#101035000000
1!
1%
#101040000000
0!
0%
#101045000000
1!
1%
#101050000000
0!
0%
#101055000000
1!
1%
#101060000000
0!
0%
#101065000000
1!
1%
#101070000000
0!
0%
#101075000000
1!
1%
#101080000000
0!
0%
#101085000000
1!
1%
#101090000000
0!
0%
#101095000000
1!
1%
#101100000000
0!
0%
#101105000000
1!
1%
#101110000000
0!
0%
#101115000000
1!
1%
#101120000000
0!
0%
#101125000000
1!
1%
#101130000000
0!
0%
#101135000000
1!
1%
#101140000000
0!
0%
#101145000000
1!
1%
#101150000000
0!
0%
#101155000000
1!
1%
#101160000000
0!
0%
#101165000000
1!
1%
#101170000000
0!
0%
#101175000000
1!
1%
#101180000000
0!
0%
#101185000000
1!
1%
#101190000000
0!
0%
#101195000000
1!
1%
#101200000000
0!
0%
#101205000000
1!
1%
#101210000000
0!
0%
#101215000000
1!
1%
#101220000000
0!
0%
#101225000000
1!
1%
#101230000000
0!
0%
#101235000000
1!
1%
#101240000000
0!
0%
#101245000000
1!
1%
#101250000000
0!
0%
#101255000000
1!
1%
#101260000000
0!
0%
#101265000000
1!
1%
#101270000000
0!
0%
#101275000000
1!
1%
#101280000000
0!
0%
#101285000000
1!
1%
#101290000000
0!
0%
#101295000000
1!
1%
#101300000000
0!
0%
#101305000000
1!
1%
#101310000000
0!
0%
#101315000000
1!
1%
#101320000000
0!
0%
#101325000000
1!
1%
#101330000000
0!
0%
#101335000000
1!
1%
#101340000000
0!
0%
#101345000000
1!
1%
#101350000000
0!
0%
#101355000000
1!
1%
#101360000000
0!
0%
#101365000000
1!
1%
#101370000000
0!
0%
#101375000000
1!
1%
#101380000000
0!
0%
#101385000000
1!
1%
#101390000000
0!
0%
#101395000000
1!
1%
#101400000000
0!
0%
#101405000000
1!
1%
#101410000000
0!
0%
#101415000000
1!
1%
#101420000000
0!
0%
#101425000000
1!
1%
#101430000000
0!
0%
#101435000000
1!
1%
#101440000000
0!
0%
#101445000000
1!
1%
#101450000000
0!
0%
#101455000000
1!
1%
#101460000000
0!
0%
#101465000000
1!
1%
#101470000000
0!
0%
#101475000000
1!
1%
#101480000000
0!
0%
#101485000000
1!
1%
#101490000000
0!
0%
#101495000000
1!
1%
#101500000000
0!
0%
#101505000000
1!
1%
#101510000000
0!
0%
#101515000000
1!
1%
#101520000000
0!
0%
#101525000000
1!
1%
#101530000000
0!
0%
#101535000000
1!
1%
#101540000000
0!
0%
#101545000000
1!
1%
#101550000000
0!
0%
#101555000000
1!
1%
#101560000000
0!
0%
#101565000000
1!
1%
#101570000000
0!
0%
#101575000000
1!
1%
#101580000000
0!
0%
#101585000000
1!
1%
#101590000000
0!
0%
#101595000000
1!
1%
#101600000000
0!
0%
#101605000000
1!
1%
#101610000000
0!
0%
#101615000000
1!
1%
#101620000000
0!
0%
#101625000000
1!
1%
#101630000000
0!
0%
#101635000000
1!
1%
#101640000000
0!
0%
#101645000000
1!
1%
#101650000000
0!
0%
#101655000000
1!
1%
#101660000000
0!
0%
#101665000000
1!
1%
#101670000000
0!
0%
#101675000000
1!
1%
#101680000000
0!
0%
#101685000000
1!
1%
#101690000000
0!
0%
#101695000000
1!
1%
#101700000000
0!
0%
#101705000000
1!
1%
#101710000000
0!
0%
#101715000000
1!
1%
#101720000000
0!
0%
#101725000000
1!
1%
#101730000000
0!
0%
#101735000000
1!
1%
#101740000000
0!
0%
#101745000000
1!
1%
#101750000000
0!
0%
#101755000000
1!
1%
#101760000000
0!
0%
#101765000000
1!
1%
#101770000000
0!
0%
#101775000000
1!
1%
#101780000000
0!
0%
#101785000000
1!
1%
#101790000000
0!
0%
#101795000000
1!
1%
#101800000000
0!
0%
#101805000000
1!
1%
#101810000000
0!
0%
#101815000000
1!
1%
#101820000000
0!
0%
#101825000000
1!
1%
#101830000000
0!
0%
#101835000000
1!
1%
#101840000000
0!
0%
#101845000000
1!
1%
#101850000000
0!
0%
#101855000000
1!
1%
#101860000000
0!
0%
#101865000000
1!
1%
#101870000000
0!
0%
#101875000000
1!
1%
#101880000000
0!
0%
#101885000000
1!
1%
#101890000000
0!
0%
#101895000000
1!
1%
#101900000000
0!
0%
#101905000000
1!
1%
#101910000000
0!
0%
#101915000000
1!
1%
#101920000000
0!
0%
#101925000000
1!
1%
#101930000000
0!
0%
#101935000000
1!
1%
#101940000000
0!
0%
#101945000000
1!
1%
#101950000000
0!
0%
#101955000000
1!
1%
#101960000000
0!
0%
#101965000000
1!
1%
#101970000000
0!
0%
#101975000000
1!
1%
#101980000000
0!
0%
#101985000000
1!
1%
#101990000000
0!
0%
#101995000000
1!
1%
#102000000000
0!
0%
#102005000000
1!
1%
#102010000000
0!
0%
#102015000000
1!
1%
#102020000000
0!
0%
#102025000000
1!
1%
#102030000000
0!
0%
#102035000000
1!
1%
#102040000000
0!
0%
#102045000000
1!
1%
#102050000000
0!
0%
#102055000000
1!
1%
#102060000000
0!
0%
#102065000000
1!
1%
#102070000000
0!
0%
#102075000000
1!
1%
#102080000000
0!
0%
#102085000000
1!
1%
#102090000000
0!
0%
#102095000000
1!
1%
#102100000000
0!
0%
#102105000000
1!
1%
#102110000000
0!
0%
#102115000000
1!
1%
#102120000000
0!
0%
#102125000000
1!
1%
#102130000000
0!
0%
#102135000000
1!
1%
#102140000000
0!
0%
#102145000000
1!
1%
#102150000000
0!
0%
#102155000000
1!
1%
#102160000000
0!
0%
#102165000000
1!
1%
#102170000000
0!
0%
#102175000000
1!
1%
#102180000000
0!
0%
#102185000000
1!
1%
#102190000000
0!
0%
#102195000000
1!
1%
#102200000000
0!
0%
#102205000000
1!
1%
#102210000000
0!
0%
#102215000000
1!
1%
#102220000000
0!
0%
#102225000000
1!
1%
#102230000000
0!
0%
#102235000000
1!
1%
#102240000000
0!
0%
#102245000000
1!
1%
#102250000000
0!
0%
#102255000000
1!
1%
#102260000000
0!
0%
#102265000000
1!
1%
#102270000000
0!
0%
#102275000000
1!
1%
#102280000000
0!
0%
#102285000000
1!
1%
#102290000000
0!
0%
#102295000000
1!
1%
#102300000000
0!
0%
#102305000000
1!
1%
#102310000000
0!
0%
#102315000000
1!
1%
#102320000000
0!
0%
#102325000000
1!
1%
#102330000000
0!
0%
#102335000000
1!
1%
#102340000000
0!
0%
#102345000000
1!
1%
#102350000000
0!
0%
#102355000000
1!
1%
#102360000000
0!
0%
#102365000000
1!
1%
#102370000000
0!
0%
#102375000000
1!
1%
#102380000000
0!
0%
#102385000000
1!
1%
#102390000000
0!
0%
#102395000000
1!
1%
#102400000000
0!
0%
#102405000000
1!
1%
#102410000000
0!
0%
#102415000000
1!
1%
#102420000000
0!
0%
#102425000000
1!
1%
#102430000000
0!
0%
#102435000000
1!
1%
#102440000000
0!
0%
#102445000000
1!
1%
#102450000000
0!
0%
#102455000000
1!
1%
#102460000000
0!
0%
#102465000000
1!
1%
#102470000000
0!
0%
#102475000000
1!
1%
#102480000000
0!
0%
#102485000000
1!
1%
#102490000000
0!
0%
#102495000000
1!
1%
#102500000000
0!
0%
#102505000000
1!
1%
#102510000000
0!
0%
#102515000000
1!
1%
#102520000000
0!
0%
#102525000000
1!
1%
#102530000000
0!
0%
#102535000000
1!
1%
#102540000000
0!
0%
#102545000000
1!
1%
#102550000000
0!
0%
#102555000000
1!
1%
#102560000000
0!
0%
#102565000000
1!
1%
#102570000000
0!
0%
#102575000000
1!
1%
#102580000000
0!
0%
#102585000000
1!
1%
#102590000000
0!
0%
#102595000000
1!
1%
#102600000000
0!
0%
#102605000000
1!
1%
#102610000000
0!
0%
#102615000000
1!
1%
#102620000000
0!
0%
#102625000000
1!
1%
#102630000000
0!
0%
#102635000000
1!
1%
#102640000000
0!
0%
#102645000000
1!
1%
#102650000000
0!
0%
#102655000000
1!
1%
#102660000000
0!
0%
#102665000000
1!
1%
#102670000000
0!
0%
#102675000000
1!
1%
#102680000000
0!
0%
#102685000000
1!
1%
#102690000000
0!
0%
#102695000000
1!
1%
#102700000000
0!
0%
#102705000000
1!
1%
#102710000000
0!
0%
#102715000000
1!
1%
#102720000000
0!
0%
#102725000000
1!
1%
#102730000000
0!
0%
#102735000000
1!
1%
#102740000000
0!
0%
#102745000000
1!
1%
#102750000000
0!
0%
#102755000000
1!
1%
#102760000000
0!
0%
#102765000000
1!
1%
#102770000000
0!
0%
#102775000000
1!
1%
#102780000000
0!
0%
#102785000000
1!
1%
#102790000000
0!
0%
#102795000000
1!
1%
#102800000000
0!
0%
#102805000000
1!
1%
#102810000000
0!
0%
#102815000000
1!
1%
#102820000000
0!
0%
#102825000000
1!
1%
#102830000000
0!
0%
#102835000000
1!
1%
#102840000000
0!
0%
#102845000000
1!
1%
#102850000000
0!
0%
#102855000000
1!
1%
#102860000000
0!
0%
#102865000000
1!
1%
#102870000000
0!
0%
#102875000000
1!
1%
#102880000000
0!
0%
#102885000000
1!
1%
#102890000000
0!
0%
#102895000000
1!
1%
#102900000000
0!
0%
#102905000000
1!
1%
#102910000000
0!
0%
#102915000000
1!
1%
#102920000000
0!
0%
#102925000000
1!
1%
#102930000000
0!
0%
#102935000000
1!
1%
#102940000000
0!
0%
#102945000000
1!
1%
#102950000000
0!
0%
#102955000000
1!
1%
#102960000000
0!
0%
#102965000000
1!
1%
#102970000000
0!
0%
#102975000000
1!
1%
#102980000000
0!
0%
#102985000000
1!
1%
#102990000000
0!
0%
#102995000000
1!
1%
#103000000000
0!
0%
#103005000000
1!
1%
#103010000000
0!
0%
#103015000000
1!
1%
#103020000000
0!
0%
#103025000000
1!
1%
#103030000000
0!
0%
#103035000000
1!
1%
#103040000000
0!
0%
#103045000000
1!
1%
#103050000000
0!
0%
#103055000000
1!
1%
#103060000000
0!
0%
#103065000000
1!
1%
#103070000000
0!
0%
#103075000000
1!
1%
#103080000000
0!
0%
#103085000000
1!
1%
#103090000000
0!
0%
#103095000000
1!
1%
#103100000000
0!
0%
#103105000000
1!
1%
#103110000000
0!
0%
#103115000000
1!
1%
#103120000000
0!
0%
#103125000000
1!
1%
#103130000000
0!
0%
#103135000000
1!
1%
#103140000000
0!
0%
#103145000000
1!
1%
#103150000000
0!
0%
#103155000000
1!
1%
#103160000000
0!
0%
#103165000000
1!
1%
#103170000000
0!
0%
#103175000000
1!
1%
#103180000000
0!
0%
#103185000000
1!
1%
#103190000000
0!
0%
#103195000000
1!
1%
#103200000000
0!
0%
#103205000000
1!
1%
#103210000000
0!
0%
#103215000000
1!
1%
#103220000000
0!
0%
#103225000000
1!
1%
#103230000000
0!
0%
#103235000000
1!
1%
#103240000000
0!
0%
#103245000000
1!
1%
#103250000000
0!
0%
#103255000000
1!
1%
#103260000000
0!
0%
#103265000000
1!
1%
#103270000000
0!
0%
#103275000000
1!
1%
#103280000000
0!
0%
#103285000000
1!
1%
#103290000000
0!
0%
#103295000000
1!
1%
#103300000000
0!
0%
#103305000000
1!
1%
#103310000000
0!
0%
#103315000000
1!
1%
#103320000000
0!
0%
#103325000000
1!
1%
#103330000000
0!
0%
#103335000000
1!
1%
#103340000000
0!
0%
#103345000000
1!
1%
#103350000000
0!
0%
#103355000000
1!
1%
#103360000000
0!
0%
#103365000000
1!
1%
#103370000000
0!
0%
#103375000000
1!
1%
#103380000000
0!
0%
#103385000000
1!
1%
#103390000000
0!
0%
#103395000000
1!
1%
#103400000000
0!
0%
#103405000000
1!
1%
#103410000000
0!
0%
#103415000000
1!
1%
#103420000000
0!
0%
#103425000000
1!
1%
#103430000000
0!
0%
#103435000000
1!
1%
#103440000000
0!
0%
#103445000000
1!
1%
#103450000000
0!
0%
#103455000000
1!
1%
#103460000000
0!
0%
#103465000000
1!
1%
#103470000000
0!
0%
#103475000000
1!
1%
#103480000000
0!
0%
#103485000000
1!
1%
#103490000000
0!
0%
#103495000000
1!
1%
#103500000000
0!
0%
#103505000000
1!
1%
#103510000000
0!
0%
#103515000000
1!
1%
#103520000000
0!
0%
#103525000000
1!
1%
#103530000000
0!
0%
#103535000000
1!
1%
#103540000000
0!
0%
#103545000000
1!
1%
#103550000000
0!
0%
#103555000000
1!
1%
#103560000000
0!
0%
#103565000000
1!
1%
#103570000000
0!
0%
#103575000000
1!
1%
#103580000000
0!
0%
#103585000000
1!
1%
#103590000000
0!
0%
#103595000000
1!
1%
#103600000000
0!
0%
#103605000000
1!
1%
#103610000000
0!
0%
#103615000000
1!
1%
#103620000000
0!
0%
#103625000000
1!
1%
#103630000000
0!
0%
#103635000000
1!
1%
#103640000000
0!
0%
#103645000000
1!
1%
#103650000000
0!
0%
#103655000000
1!
1%
#103660000000
0!
0%
#103665000000
1!
1%
#103670000000
0!
0%
#103675000000
1!
1%
#103680000000
0!
0%
#103685000000
1!
1%
#103690000000
0!
0%
#103695000000
1!
1%
#103700000000
0!
0%
#103705000000
1!
1%
#103710000000
0!
0%
#103715000000
1!
1%
#103720000000
0!
0%
#103725000000
1!
1%
#103730000000
0!
0%
#103735000000
1!
1%
#103740000000
0!
0%
#103745000000
1!
1%
#103750000000
0!
0%
#103755000000
1!
1%
#103760000000
0!
0%
#103765000000
1!
1%
#103770000000
0!
0%
#103775000000
1!
1%
#103780000000
0!
0%
#103785000000
1!
1%
#103790000000
0!
0%
#103795000000
1!
1%
#103800000000
0!
0%
#103805000000
1!
1%
#103810000000
0!
0%
#103815000000
1!
1%
#103820000000
0!
0%
#103825000000
1!
1%
#103830000000
0!
0%
#103835000000
1!
1%
#103840000000
0!
0%
#103845000000
1!
1%
#103850000000
0!
0%
#103855000000
1!
1%
#103860000000
0!
0%
#103865000000
1!
1%
#103870000000
0!
0%
#103875000000
1!
1%
#103880000000
0!
0%
#103885000000
1!
1%
#103890000000
0!
0%
#103895000000
1!
1%
#103900000000
0!
0%
#103905000000
1!
1%
#103910000000
0!
0%
#103915000000
1!
1%
#103920000000
0!
0%
#103925000000
1!
1%
#103930000000
0!
0%
#103935000000
1!
1%
#103940000000
0!
0%
#103945000000
1!
1%
#103950000000
0!
0%
#103955000000
1!
1%
#103960000000
0!
0%
#103965000000
1!
1%
#103970000000
0!
0%
#103975000000
1!
1%
#103980000000
0!
0%
#103985000000
1!
1%
#103990000000
0!
0%
#103995000000
1!
1%
#104000000000
0!
0%
#104005000000
1!
1%
#104010000000
0!
0%
#104015000000
1!
1%
#104020000000
0!
0%
#104025000000
1!
1%
#104030000000
0!
0%
#104035000000
1!
1%
#104040000000
0!
0%
#104045000000
1!
1%
#104050000000
0!
0%
#104055000000
1!
1%
#104060000000
0!
0%
#104065000000
1!
1%
#104070000000
0!
0%
#104075000000
1!
1%
#104080000000
0!
0%
#104085000000
1!
1%
#104090000000
0!
0%
#104095000000
1!
1%
#104100000000
0!
0%
#104105000000
1!
1%
#104110000000
0!
0%
#104115000000
1!
1%
#104120000000
0!
0%
#104125000000
1!
1%
#104130000000
0!
0%
#104135000000
1!
1%
#104140000000
0!
0%
#104145000000
1!
1%
#104150000000
0!
0%
#104155000000
1!
1%
#104160000000
0!
0%
#104165000000
1!
1%
#104170000000
0!
0%
#104175000000
1!
1%
#104180000000
0!
0%
#104185000000
1!
1%
#104190000000
0!
0%
#104195000000
1!
1%
#104200000000
0!
0%
#104205000000
1!
1%
#104210000000
0!
0%
#104215000000
1!
1%
#104220000000
0!
0%
#104225000000
1!
1%
#104230000000
0!
0%
#104235000000
1!
1%
#104240000000
0!
0%
#104245000000
1!
1%
#104250000000
0!
0%
#104255000000
1!
1%
#104260000000
0!
0%
#104265000000
1!
1%
#104270000000
0!
0%
#104275000000
1!
1%
#104280000000
0!
0%
#104285000000
1!
1%
#104290000000
0!
0%
#104295000000
1!
1%
#104300000000
0!
0%
#104305000000
1!
1%
#104310000000
0!
0%
#104315000000
1!
1%
#104320000000
0!
0%
#104325000000
1!
1%
#104330000000
0!
0%
#104335000000
1!
1%
#104340000000
0!
0%
#104345000000
1!
1%
#104350000000
0!
0%
#104355000000
1!
1%
#104360000000
0!
0%
#104365000000
1!
1%
#104370000000
0!
0%
#104375000000
1!
1%
#104380000000
0!
0%
#104385000000
1!
1%
#104390000000
0!
0%
#104395000000
1!
1%
#104400000000
0!
0%
#104405000000
1!
1%
#104410000000
0!
0%
#104415000000
1!
1%
#104420000000
0!
0%
#104425000000
1!
1%
#104430000000
0!
0%
#104435000000
1!
1%
#104440000000
0!
0%
#104445000000
1!
1%
#104450000000
0!
0%
#104455000000
1!
1%
#104460000000
0!
0%
#104465000000
1!
1%
#104470000000
0!
0%
#104475000000
1!
1%
#104480000000
0!
0%
#104485000000
1!
1%
#104490000000
0!
0%
#104495000000
1!
1%
#104500000000
0!
0%
#104505000000
1!
1%
#104510000000
0!
0%
#104515000000
1!
1%
#104520000000
0!
0%
#104525000000
1!
1%
#104530000000
0!
0%
#104535000000
1!
1%
#104540000000
0!
0%
#104545000000
1!
1%
#104550000000
0!
0%
#104555000000
1!
1%
#104560000000
0!
0%
#104565000000
1!
1%
#104570000000
0!
0%
#104575000000
1!
1%
#104580000000
0!
0%
#104585000000
1!
1%
#104590000000
0!
0%
#104595000000
1!
1%
#104600000000
0!
0%
#104605000000
1!
1%
#104610000000
0!
0%
#104615000000
1!
1%
#104620000000
0!
0%
#104625000000
1!
1%
#104630000000
0!
0%
#104635000000
1!
1%
#104640000000
0!
0%
#104645000000
1!
1%
#104650000000
0!
0%
#104655000000
1!
1%
#104660000000
0!
0%
#104665000000
1!
1%
#104670000000
0!
0%
#104675000000
1!
1%
#104680000000
0!
0%
#104685000000
1!
1%
#104690000000
0!
0%
#104695000000
1!
1%
#104700000000
0!
0%
#104705000000
1!
1%
#104710000000
0!
0%
#104715000000
1!
1%
#104720000000
0!
0%
#104725000000
1!
1%
#104730000000
0!
0%
#104735000000
1!
1%
#104740000000
0!
0%
#104745000000
1!
1%
#104750000000
0!
0%
#104755000000
1!
1%
#104760000000
0!
0%
#104765000000
1!
1%
#104770000000
0!
0%
#104775000000
1!
1%
#104780000000
0!
0%
#104785000000
1!
1%
#104790000000
0!
0%
#104795000000
1!
1%
#104800000000
0!
0%
#104805000000
1!
1%
#104810000000
0!
0%
#104815000000
1!
1%
#104820000000
0!
0%
#104825000000
1!
1%
#104830000000
0!
0%
#104835000000
1!
1%
#104840000000
0!
0%
#104845000000
1!
1%
#104850000000
0!
0%
#104855000000
1!
1%
#104860000000
0!
0%
#104865000000
1!
1%
#104870000000
0!
0%
#104875000000
1!
1%
#104880000000
0!
0%
#104885000000
1!
1%
#104890000000
0!
0%
#104895000000
1!
1%
#104900000000
0!
0%
#104905000000
1!
1%
#104910000000
0!
0%
#104915000000
1!
1%
#104920000000
0!
0%
#104925000000
1!
1%
#104930000000
0!
0%
#104935000000
1!
1%
#104940000000
0!
0%
#104945000000
1!
1%
#104950000000
0!
0%
#104955000000
1!
1%
#104960000000
0!
0%
#104965000000
1!
1%
#104970000000
0!
0%
#104975000000
1!
1%
#104980000000
0!
0%
#104985000000
1!
1%
#104990000000
0!
0%
#104995000000
1!
1%
#105000000000
0!
0%
#105005000000
1!
1%
#105010000000
0!
0%
#105015000000
1!
1%
#105020000000
0!
0%
#105025000000
1!
1%
#105030000000
0!
0%
#105035000000
1!
1%
#105040000000
0!
0%
#105045000000
1!
1%
#105050000000
0!
0%
#105055000000
1!
1%
#105060000000
0!
0%
#105065000000
1!
1%
#105070000000
0!
0%
#105075000000
1!
1%
#105080000000
0!
0%
#105085000000
1!
1%
#105090000000
0!
0%
#105095000000
1!
1%
#105100000000
0!
0%
#105105000000
1!
1%
#105110000000
0!
0%
#105115000000
1!
1%
#105120000000
0!
0%
#105125000000
1!
1%
#105130000000
0!
0%
#105135000000
1!
1%
#105140000000
0!
0%
#105145000000
1!
1%
#105150000000
0!
0%
#105155000000
1!
1%
#105160000000
0!
0%
#105165000000
1!
1%
#105170000000
0!
0%
#105175000000
1!
1%
#105180000000
0!
0%
#105185000000
1!
1%
#105190000000
0!
0%
#105195000000
1!
1%
#105200000000
0!
0%
#105205000000
1!
1%
#105210000000
0!
0%
#105215000000
1!
1%
#105220000000
0!
0%
#105225000000
1!
1%
#105230000000
0!
0%
#105235000000
1!
1%
#105240000000
0!
0%
#105245000000
1!
1%
#105250000000
0!
0%
#105255000000
1!
1%
#105260000000
0!
0%
#105265000000
1!
1%
#105270000000
0!
0%
#105275000000
1!
1%
#105280000000
0!
0%
#105285000000
1!
1%
#105290000000
0!
0%
#105295000000
1!
1%
#105300000000
0!
0%
#105305000000
1!
1%
#105310000000
0!
0%
#105315000000
1!
1%
#105320000000
0!
0%
#105325000000
1!
1%
#105330000000
0!
0%
#105335000000
1!
1%
#105340000000
0!
0%
#105345000000
1!
1%
#105350000000
0!
0%
#105355000000
1!
1%
#105360000000
0!
0%
#105365000000
1!
1%
#105370000000
0!
0%
#105375000000
1!
1%
#105380000000
0!
0%
#105385000000
1!
1%
#105390000000
0!
0%
#105395000000
1!
1%
#105400000000
0!
0%
#105405000000
1!
1%
#105410000000
0!
0%
#105415000000
1!
1%
#105420000000
0!
0%
#105425000000
1!
1%
#105430000000
0!
0%
#105435000000
1!
1%
#105440000000
0!
0%
#105445000000
1!
1%
#105450000000
0!
0%
#105455000000
1!
1%
#105460000000
0!
0%
#105465000000
1!
1%
#105470000000
0!
0%
#105475000000
1!
1%
#105480000000
0!
0%
#105485000000
1!
1%
#105490000000
0!
0%
#105495000000
1!
1%
#105500000000
0!
0%
#105505000000
1!
1%
#105510000000
0!
0%
#105515000000
1!
1%
#105520000000
0!
0%
#105525000000
1!
1%
#105530000000
0!
0%
#105535000000
1!
1%
#105540000000
0!
0%
#105545000000
1!
1%
#105550000000
0!
0%
#105555000000
1!
1%
#105560000000
0!
0%
#105565000000
1!
1%
#105570000000
0!
0%
#105575000000
1!
1%
#105580000000
0!
0%
#105585000000
1!
1%
#105590000000
0!
0%
#105595000000
1!
1%
#105600000000
0!
0%
#105605000000
1!
1%
#105610000000
0!
0%
#105615000000
1!
1%
#105620000000
0!
0%
#105625000000
1!
1%
#105630000000
0!
0%
#105635000000
1!
1%
#105640000000
0!
0%
#105645000000
1!
1%
#105650000000
0!
0%
#105655000000
1!
1%
#105660000000
0!
0%
#105665000000
1!
1%
#105670000000
0!
0%
#105675000000
1!
1%
#105680000000
0!
0%
#105685000000
1!
1%
#105690000000
0!
0%
#105695000000
1!
1%
#105700000000
0!
0%
#105705000000
1!
1%
#105710000000
0!
0%
#105715000000
1!
1%
#105720000000
0!
0%
#105725000000
1!
1%
#105730000000
0!
0%
#105735000000
1!
1%
#105740000000
0!
0%
#105745000000
1!
1%
#105750000000
0!
0%
#105755000000
1!
1%
#105760000000
0!
0%
#105765000000
1!
1%
#105770000000
0!
0%
#105775000000
1!
1%
#105780000000
0!
0%
#105785000000
1!
1%
#105790000000
0!
0%
#105795000000
1!
1%
#105800000000
0!
0%
#105805000000
1!
1%
#105810000000
0!
0%
#105815000000
1!
1%
#105820000000
0!
0%
#105825000000
1!
1%
#105830000000
0!
0%
#105835000000
1!
1%
#105840000000
0!
0%
#105845000000
1!
1%
#105850000000
0!
0%
#105855000000
1!
1%
#105860000000
0!
0%
#105865000000
1!
1%
#105870000000
0!
0%
#105875000000
1!
1%
#105880000000
0!
0%
#105885000000
1!
1%
#105890000000
0!
0%
#105895000000
1!
1%
#105900000000
0!
0%
#105905000000
1!
1%
#105910000000
0!
0%
#105915000000
1!
1%
#105920000000
0!
0%
#105925000000
1!
1%
#105930000000
0!
0%
#105935000000
1!
1%
#105940000000
0!
0%
#105945000000
1!
1%
#105950000000
0!
0%
#105955000000
1!
1%
#105960000000
0!
0%
#105965000000
1!
1%
#105970000000
0!
0%
#105975000000
1!
1%
#105980000000
0!
0%
#105985000000
1!
1%
#105990000000
0!
0%
#105995000000
1!
1%
#106000000000
0!
0%
#106005000000
1!
1%
#106010000000
0!
0%
#106015000000
1!
1%
#106020000000
0!
0%
#106025000000
1!
1%
#106030000000
0!
0%
#106035000000
1!
1%
#106040000000
0!
0%
#106045000000
1!
1%
#106050000000
0!
0%
#106055000000
1!
1%
#106060000000
0!
0%
#106065000000
1!
1%
#106070000000
0!
0%
#106075000000
1!
1%
#106080000000
0!
0%
#106085000000
1!
1%
#106090000000
0!
0%
#106095000000
1!
1%
#106100000000
0!
0%
#106105000000
1!
1%
#106110000000
0!
0%
#106115000000
1!
1%
#106120000000
0!
0%
#106125000000
1!
1%
#106130000000
0!
0%
#106135000000
1!
1%
#106140000000
0!
0%
#106145000000
1!
1%
#106150000000
0!
0%
#106155000000
1!
1%
#106160000000
0!
0%
#106165000000
1!
1%
#106170000000
0!
0%
#106175000000
1!
1%
#106180000000
0!
0%
#106185000000
1!
1%
#106190000000
0!
0%
#106195000000
1!
1%
#106200000000
0!
0%
#106205000000
1!
1%
#106210000000
0!
0%
#106215000000
1!
1%
#106220000000
0!
0%
#106225000000
1!
1%
#106230000000
0!
0%
#106235000000
1!
1%
#106240000000
0!
0%
#106245000000
1!
1%
#106250000000
0!
0%
#106255000000
1!
1%
#106260000000
0!
0%
#106265000000
1!
1%
#106270000000
0!
0%
#106275000000
1!
1%
#106280000000
0!
0%
#106285000000
1!
1%
#106290000000
0!
0%
#106295000000
1!
1%
#106300000000
0!
0%
#106305000000
1!
1%
#106310000000
0!
0%
#106315000000
1!
1%
#106320000000
0!
0%
#106325000000
1!
1%
#106330000000
0!
0%
#106335000000
1!
1%
#106340000000
0!
0%
#106345000000
1!
1%
#106350000000
0!
0%
#106355000000
1!
1%
#106360000000
0!
0%
#106365000000
1!
1%
#106370000000
0!
0%
#106375000000
1!
1%
#106380000000
0!
0%
#106385000000
1!
1%
#106390000000
0!
0%
#106395000000
1!
1%
#106400000000
0!
0%
#106405000000
1!
1%
#106410000000
0!
0%
#106415000000
1!
1%
#106420000000
0!
0%
#106425000000
1!
1%
#106430000000
0!
0%
#106435000000
1!
1%
#106440000000
0!
0%
#106445000000
1!
1%
#106450000000
0!
0%
#106455000000
1!
1%
#106460000000
0!
0%
#106465000000
1!
1%
#106470000000
0!
0%
#106475000000
1!
1%
#106480000000
0!
0%
#106485000000
1!
1%
#106490000000
0!
0%
#106495000000
1!
1%
#106500000000
0!
0%
#106505000000
1!
1%
#106510000000
0!
0%
#106515000000
1!
1%
#106520000000
0!
0%
#106525000000
1!
1%
#106530000000
0!
0%
#106535000000
1!
1%
#106540000000
0!
0%
#106545000000
1!
1%
#106550000000
0!
0%
#106555000000
1!
1%
#106560000000
0!
0%
#106565000000
1!
1%
#106570000000
0!
0%
#106575000000
1!
1%
#106580000000
0!
0%
#106585000000
1!
1%
#106590000000
0!
0%
#106595000000
1!
1%
#106600000000
0!
0%
#106605000000
1!
1%
#106610000000
0!
0%
#106615000000
1!
1%
#106620000000
0!
0%
#106625000000
1!
1%
#106630000000
0!
0%
#106635000000
1!
1%
#106640000000
0!
0%
#106645000000
1!
1%
#106650000000
0!
0%
#106655000000
1!
1%
#106660000000
0!
0%
#106665000000
1!
1%
#106670000000
0!
0%
#106675000000
1!
1%
#106680000000
0!
0%
#106685000000
1!
1%
#106690000000
0!
0%
#106695000000
1!
1%
#106700000000
0!
0%
#106705000000
1!
1%
#106710000000
0!
0%
#106715000000
1!
1%
#106720000000
0!
0%
#106725000000
1!
1%
#106730000000
0!
0%
#106735000000
1!
1%
#106740000000
0!
0%
#106745000000
1!
1%
#106750000000
0!
0%
#106755000000
1!
1%
#106760000000
0!
0%
#106765000000
1!
1%
#106770000000
0!
0%
#106775000000
1!
1%
#106780000000
0!
0%
#106785000000
1!
1%
#106790000000
0!
0%
#106795000000
1!
1%
#106800000000
0!
0%
#106805000000
1!
1%
#106810000000
0!
0%
#106815000000
1!
1%
#106820000000
0!
0%
#106825000000
1!
1%
#106830000000
0!
0%
#106835000000
1!
1%
#106840000000
0!
0%
#106845000000
1!
1%
#106850000000
0!
0%
#106855000000
1!
1%
#106860000000
0!
0%
#106865000000
1!
1%
#106870000000
0!
0%
#106875000000
1!
1%
#106880000000
0!
0%
#106885000000
1!
1%
#106890000000
0!
0%
#106895000000
1!
1%
#106900000000
0!
0%
#106905000000
1!
1%
#106910000000
0!
0%
#106915000000
1!
1%
#106920000000
0!
0%
#106925000000
1!
1%
#106930000000
0!
0%
#106935000000
1!
1%
#106940000000
0!
0%
#106945000000
1!
1%
#106950000000
0!
0%
#106955000000
1!
1%
#106960000000
0!
0%
#106965000000
1!
1%
#106970000000
0!
0%
#106975000000
1!
1%
#106980000000
0!
0%
#106985000000
1!
1%
#106990000000
0!
0%
#106995000000
1!
1%
#107000000000
0!
0%
#107005000000
1!
1%
#107010000000
0!
0%
#107015000000
1!
1%
#107020000000
0!
0%
#107025000000
1!
1%
#107030000000
0!
0%
#107035000000
1!
1%
#107040000000
0!
0%
#107045000000
1!
1%
#107050000000
0!
0%
#107055000000
1!
1%
#107060000000
0!
0%
#107065000000
1!
1%
#107070000000
0!
0%
#107075000000
1!
1%
#107080000000
0!
0%
#107085000000
1!
1%
#107090000000
0!
0%
#107095000000
1!
1%
#107100000000
0!
0%
#107105000000
1!
1%
#107110000000
0!
0%
#107115000000
1!
1%
#107120000000
0!
0%
#107125000000
1!
1%
#107130000000
0!
0%
#107135000000
1!
1%
#107140000000
0!
0%
#107145000000
1!
1%
#107150000000
0!
0%
#107155000000
1!
1%
#107160000000
0!
0%
#107165000000
1!
1%
#107170000000
0!
0%
#107175000000
1!
1%
#107180000000
0!
0%
#107185000000
1!
1%
#107190000000
0!
0%
#107195000000
1!
1%
#107200000000
0!
0%
#107205000000
1!
1%
#107210000000
0!
0%
#107215000000
1!
1%
#107220000000
0!
0%
#107225000000
1!
1%
#107230000000
0!
0%
#107235000000
1!
1%
#107240000000
0!
0%
#107245000000
1!
1%
#107250000000
0!
0%
#107255000000
1!
1%
#107260000000
0!
0%
#107265000000
1!
1%
#107270000000
0!
0%
#107275000000
1!
1%
#107280000000
0!
0%
#107285000000
1!
1%
#107290000000
0!
0%
#107295000000
1!
1%
#107300000000
0!
0%
#107305000000
1!
1%
#107310000000
0!
0%
#107315000000
1!
1%
#107320000000
0!
0%
#107325000000
1!
1%
#107330000000
0!
0%
#107335000000
1!
1%
#107340000000
0!
0%
#107345000000
1!
1%
#107350000000
0!
0%
#107355000000
1!
1%
#107360000000
0!
0%
#107365000000
1!
1%
#107370000000
0!
0%
#107375000000
1!
1%
#107380000000
0!
0%
#107385000000
1!
1%
#107390000000
0!
0%
#107395000000
1!
1%
#107400000000
0!
0%
#107405000000
1!
1%
#107410000000
0!
0%
#107415000000
1!
1%
#107420000000
0!
0%
#107425000000
1!
1%
#107430000000
0!
0%
#107435000000
1!
1%
#107440000000
0!
0%
#107445000000
1!
1%
#107450000000
0!
0%
#107455000000
1!
1%
#107460000000
0!
0%
#107465000000
1!
1%
#107470000000
0!
0%
#107475000000
1!
1%
#107480000000
0!
0%
#107485000000
1!
1%
#107490000000
0!
0%
#107495000000
1!
1%
#107500000000
0!
0%
#107505000000
1!
1%
#107510000000
0!
0%
#107515000000
1!
1%
#107520000000
0!
0%
#107525000000
1!
1%
#107530000000
0!
0%
#107535000000
1!
1%
#107540000000
0!
0%
#107545000000
1!
1%
#107550000000
0!
0%
#107555000000
1!
1%
#107560000000
0!
0%
#107565000000
1!
1%
#107570000000
0!
0%
#107575000000
1!
1%
#107580000000
0!
0%
#107585000000
1!
1%
#107590000000
0!
0%
#107595000000
1!
1%
#107600000000
0!
0%
#107605000000
1!
1%
#107610000000
0!
0%
#107615000000
1!
1%
#107620000000
0!
0%
#107625000000
1!
1%
#107630000000
0!
0%
#107635000000
1!
1%
#107640000000
0!
0%
#107645000000
1!
1%
#107650000000
0!
0%
#107655000000
1!
1%
#107660000000
0!
0%
#107665000000
1!
1%
#107670000000
0!
0%
#107675000000
1!
1%
#107680000000
0!
0%
#107685000000
1!
1%
#107690000000
0!
0%
#107695000000
1!
1%
#107700000000
0!
0%
#107705000000
1!
1%
#107710000000
0!
0%
#107715000000
1!
1%
#107720000000
0!
0%
#107725000000
1!
1%
#107730000000
0!
0%
#107735000000
1!
1%
#107740000000
0!
0%
#107745000000
1!
1%
#107750000000
0!
0%
#107755000000
1!
1%
#107760000000
0!
0%
#107765000000
1!
1%
#107770000000
0!
0%
#107775000000
1!
1%
#107780000000
0!
0%
#107785000000
1!
1%
#107790000000
0!
0%
#107795000000
1!
1%
#107800000000
0!
0%
#107805000000
1!
1%
#107810000000
0!
0%
#107815000000
1!
1%
#107820000000
0!
0%
#107825000000
1!
1%
#107830000000
0!
0%
#107835000000
1!
1%
#107840000000
0!
0%
#107845000000
1!
1%
#107850000000
0!
0%
#107855000000
1!
1%
#107860000000
0!
0%
#107865000000
1!
1%
#107870000000
0!
0%
#107875000000
1!
1%
#107880000000
0!
0%
#107885000000
1!
1%
#107890000000
0!
0%
#107895000000
1!
1%
#107900000000
0!
0%
#107905000000
1!
1%
#107910000000
0!
0%
#107915000000
1!
1%
#107920000000
0!
0%
#107925000000
1!
1%
#107930000000
0!
0%
#107935000000
1!
1%
#107940000000
0!
0%
#107945000000
1!
1%
#107950000000
0!
0%
#107955000000
1!
1%
#107960000000
0!
0%
#107965000000
1!
1%
#107970000000
0!
0%
#107975000000
1!
1%
#107980000000
0!
0%
#107985000000
1!
1%
#107990000000
0!
0%
#107995000000
1!
1%
#108000000000
0!
0%
#108005000000
1!
1%
#108010000000
0!
0%
#108015000000
1!
1%
#108020000000
0!
0%
#108025000000
1!
1%
#108030000000
0!
0%
#108035000000
1!
1%
#108040000000
0!
0%
#108045000000
1!
1%
#108050000000
0!
0%
#108055000000
1!
1%
#108060000000
0!
0%
#108065000000
1!
1%
#108070000000
0!
0%
#108075000000
1!
1%
#108080000000
0!
0%
#108085000000
1!
1%
#108090000000
0!
0%
#108095000000
1!
1%
#108100000000
0!
0%
#108105000000
1!
1%
#108110000000
0!
0%
#108115000000
1!
1%
#108120000000
0!
0%
#108125000000
1!
1%
#108130000000
0!
0%
#108135000000
1!
1%
#108140000000
0!
0%
#108145000000
1!
1%
#108150000000
0!
0%
#108155000000
1!
1%
#108160000000
0!
0%
#108165000000
1!
1%
#108170000000
0!
0%
#108175000000
1!
1%
#108180000000
0!
0%
#108185000000
1!
1%
#108190000000
0!
0%
#108195000000
1!
1%
#108200000000
0!
0%
#108205000000
1!
1%
#108210000000
0!
0%
#108215000000
1!
1%
#108220000000
0!
0%
#108225000000
1!
1%
#108230000000
0!
0%
#108235000000
1!
1%
#108240000000
0!
0%
#108245000000
1!
1%
#108250000000
0!
0%
#108255000000
1!
1%
#108260000000
0!
0%
#108265000000
1!
1%
#108270000000
0!
0%
#108275000000
1!
1%
#108280000000
0!
0%
#108285000000
1!
1%
#108290000000
0!
0%
#108295000000
1!
1%
#108300000000
0!
0%
#108305000000
1!
1%
#108310000000
0!
0%
#108315000000
1!
1%
#108320000000
0!
0%
#108325000000
1!
1%
#108330000000
0!
0%
#108335000000
1!
1%
#108340000000
0!
0%
#108345000000
1!
1%
#108350000000
0!
0%
#108355000000
1!
1%
#108360000000
0!
0%
#108365000000
1!
1%
#108370000000
0!
0%
#108375000000
1!
1%
#108380000000
0!
0%
#108385000000
1!
1%
#108390000000
0!
0%
#108395000000
1!
1%
#108400000000
0!
0%
#108405000000
1!
1%
#108410000000
0!
0%
#108415000000
1!
1%
#108420000000
0!
0%
#108425000000
1!
1%
#108430000000
0!
0%
#108435000000
1!
1%
#108440000000
0!
0%
#108445000000
1!
1%
#108450000000
0!
0%
#108455000000
1!
1%
#108460000000
0!
0%
#108465000000
1!
1%
#108470000000
0!
0%
#108475000000
1!
1%
#108480000000
0!
0%
#108485000000
1!
1%
#108490000000
0!
0%
#108495000000
1!
1%
#108500000000
0!
0%
#108505000000
1!
1%
#108510000000
0!
0%
#108515000000
1!
1%
#108520000000
0!
0%
#108525000000
1!
1%
#108530000000
0!
0%
#108535000000
1!
1%
#108540000000
0!
0%
#108545000000
1!
1%
#108550000000
0!
0%
#108555000000
1!
1%
#108560000000
0!
0%
#108565000000
1!
1%
#108570000000
0!
0%
#108575000000
1!
1%
#108580000000
0!
0%
#108585000000
1!
1%
#108590000000
0!
0%
#108595000000
1!
1%
#108600000000
0!
0%
#108605000000
1!
1%
#108610000000
0!
0%
#108615000000
1!
1%
#108620000000
0!
0%
#108625000000
1!
1%
#108630000000
0!
0%
#108635000000
1!
1%
#108640000000
0!
0%
#108645000000
1!
1%
#108650000000
0!
0%
#108655000000
1!
1%
#108660000000
0!
0%
#108665000000
1!
1%
#108670000000
0!
0%
#108675000000
1!
1%
#108680000000
0!
0%
#108685000000
1!
1%
#108690000000
0!
0%
#108695000000
1!
1%
#108700000000
0!
0%
#108705000000
1!
1%
#108710000000
0!
0%
#108715000000
1!
1%
#108720000000
0!
0%
#108725000000
1!
1%
#108730000000
0!
0%
#108735000000
1!
1%
#108740000000
0!
0%
#108745000000
1!
1%
#108750000000
0!
0%
#108755000000
1!
1%
#108760000000
0!
0%
#108765000000
1!
1%
#108770000000
0!
0%
#108775000000
1!
1%
#108780000000
0!
0%
#108785000000
1!
1%
#108790000000
0!
0%
#108795000000
1!
1%
#108800000000
0!
0%
#108805000000
1!
1%
#108810000000
0!
0%
#108815000000
1!
1%
#108820000000
0!
0%
#108825000000
1!
1%
#108830000000
0!
0%
#108835000000
1!
1%
#108840000000
0!
0%
#108845000000
1!
1%
#108850000000
0!
0%
#108855000000
1!
1%
#108860000000
0!
0%
#108865000000
1!
1%
#108870000000
0!
0%
#108875000000
1!
1%
#108880000000
0!
0%
#108885000000
1!
1%
#108890000000
0!
0%
#108895000000
1!
1%
#108900000000
0!
0%
#108905000000
1!
1%
#108910000000
0!
0%
#108915000000
1!
1%
#108920000000
0!
0%
#108925000000
1!
1%
#108930000000
0!
0%
#108935000000
1!
1%
#108940000000
0!
0%
#108945000000
1!
1%
#108950000000
0!
0%
#108955000000
1!
1%
#108960000000
0!
0%
#108965000000
1!
1%
#108970000000
0!
0%
#108975000000
1!
1%
#108980000000
0!
0%
#108985000000
1!
1%
#108990000000
0!
0%
#108995000000
1!
1%
#109000000000
0!
0%
#109005000000
1!
1%
#109010000000
0!
0%
#109015000000
1!
1%
#109020000000
0!
0%
#109025000000
1!
1%
#109030000000
0!
0%
#109035000000
1!
1%
#109040000000
0!
0%
#109045000000
1!
1%
#109050000000
0!
0%
#109055000000
1!
1%
#109060000000
0!
0%
#109065000000
1!
1%
#109070000000
0!
0%
#109075000000
1!
1%
#109080000000
0!
0%
#109085000000
1!
1%
#109090000000
0!
0%
#109095000000
1!
1%
#109100000000
0!
0%
#109105000000
1!
1%
#109110000000
0!
0%
#109115000000
1!
1%
#109120000000
0!
0%
#109125000000
1!
1%
#109130000000
0!
0%
#109135000000
1!
1%
#109140000000
0!
0%
#109145000000
1!
1%
#109150000000
0!
0%
#109155000000
1!
1%
#109160000000
0!
0%
#109165000000
1!
1%
#109170000000
0!
0%
#109175000000
1!
1%
#109180000000
0!
0%
#109185000000
1!
1%
#109190000000
0!
0%
#109195000000
1!
1%
#109200000000
0!
0%
#109205000000
1!
1%
#109210000000
0!
0%
#109215000000
1!
1%
#109220000000
0!
0%
#109225000000
1!
1%
#109230000000
0!
0%
#109235000000
1!
1%
#109240000000
0!
0%
#109245000000
1!
1%
#109250000000
0!
0%
#109255000000
1!
1%
#109260000000
0!
0%
#109265000000
1!
1%
#109270000000
0!
0%
#109275000000
1!
1%
#109280000000
0!
0%
#109285000000
1!
1%
#109290000000
0!
0%
#109295000000
1!
1%
#109300000000
0!
0%
#109305000000
1!
1%
#109310000000
0!
0%
#109315000000
1!
1%
#109320000000
0!
0%
#109325000000
1!
1%
#109330000000
0!
0%
#109335000000
1!
1%
#109340000000
0!
0%
#109345000000
1!
1%
#109350000000
0!
0%
#109355000000
1!
1%
#109360000000
0!
0%
#109365000000
1!
1%
#109370000000
0!
0%
#109375000000
1!
1%
#109380000000
0!
0%
#109385000000
1!
1%
#109390000000
0!
0%
#109395000000
1!
1%
#109400000000
0!
0%
#109405000000
1!
1%
#109410000000
0!
0%
#109415000000
1!
1%
#109420000000
0!
0%
#109425000000
1!
1%
#109430000000
0!
0%
#109435000000
1!
1%
#109440000000
0!
0%
#109445000000
1!
1%
#109450000000
0!
0%
#109455000000
1!
1%
#109460000000
0!
0%
#109465000000
1!
1%
#109470000000
0!
0%
#109475000000
1!
1%
#109480000000
0!
0%
#109485000000
1!
1%
#109490000000
0!
0%
#109495000000
1!
1%
#109500000000
0!
0%
#109505000000
1!
1%
#109510000000
0!
0%
#109515000000
1!
1%
#109520000000
0!
0%
#109525000000
1!
1%
#109530000000
0!
0%
#109535000000
1!
1%
#109540000000
0!
0%
#109545000000
1!
1%
#109550000000
0!
0%
#109555000000
1!
1%
#109560000000
0!
0%
#109565000000
1!
1%
#109570000000
0!
0%
#109575000000
1!
1%
#109580000000
0!
0%
#109585000000
1!
1%
#109590000000
0!
0%
#109595000000
1!
1%
#109600000000
0!
0%
#109605000000
1!
1%
#109610000000
0!
0%
#109615000000
1!
1%
#109620000000
0!
0%
#109625000000
1!
1%
#109630000000
0!
0%
#109635000000
1!
1%
#109640000000
0!
0%
#109645000000
1!
1%
#109650000000
0!
0%
#109655000000
1!
1%
#109660000000
0!
0%
#109665000000
1!
1%
#109670000000
0!
0%
#109675000000
1!
1%
#109680000000
0!
0%
#109685000000
1!
1%
#109690000000
0!
0%
#109695000000
1!
1%
#109700000000
0!
0%
#109705000000
1!
1%
#109710000000
0!
0%
#109715000000
1!
1%
#109720000000
0!
0%
#109725000000
1!
1%
#109730000000
0!
0%
#109735000000
1!
1%
#109740000000
0!
0%
#109745000000
1!
1%
#109750000000
0!
0%
#109755000000
1!
1%
#109760000000
0!
0%
#109765000000
1!
1%
#109770000000
0!
0%
#109775000000
1!
1%
#109780000000
0!
0%
#109785000000
1!
1%
#109790000000
0!
0%
#109795000000
1!
1%
#109800000000
0!
0%
#109805000000
1!
1%
#109810000000
0!
0%
#109815000000
1!
1%
#109820000000
0!
0%
#109825000000
1!
1%
#109830000000
0!
0%
#109835000000
1!
1%
#109840000000
0!
0%
#109845000000
1!
1%
#109850000000
0!
0%
#109855000000
1!
1%
#109860000000
0!
0%
#109865000000
1!
1%
#109870000000
0!
0%
#109875000000
1!
1%
#109880000000
0!
0%
#109885000000
1!
1%
#109890000000
0!
0%
#109895000000
1!
1%
#109900000000
0!
0%
#109905000000
1!
1%
#109910000000
0!
0%
#109915000000
1!
1%
#109920000000
0!
0%
#109925000000
1!
1%
#109930000000
0!
0%
#109935000000
1!
1%
#109940000000
0!
0%
#109945000000
1!
1%
#109950000000
0!
0%
#109955000000
1!
1%
#109960000000
0!
0%
#109965000000
1!
1%
#109970000000
0!
0%
#109975000000
1!
1%
#109980000000
0!
0%
#109985000000
1!
1%
#109990000000
0!
0%
#109995000000
1!
1%
#110000000000
0!
0%
#110005000000
1!
1%
#110010000000
0!
0%
#110015000000
1!
1%
#110020000000
0!
0%
#110025000000
1!
1%
#110030000000
0!
0%
#110035000000
1!
1%
#110040000000
0!
0%
#110045000000
1!
1%
#110050000000
0!
0%
#110055000000
1!
1%
#110060000000
0!
0%
#110065000000
1!
1%
#110070000000
0!
0%
#110075000000
1!
1%
#110080000000
0!
0%
#110085000000
1!
1%
#110090000000
0!
0%
#110095000000
1!
1%
#110100000000
0!
0%
#110105000000
1!
1%
#110110000000
0!
0%
#110115000000
1!
1%
#110120000000
0!
0%
#110125000000
1!
1%
#110130000000
0!
0%
#110135000000
1!
1%
#110140000000
0!
0%
#110145000000
1!
1%
#110150000000
0!
0%
#110155000000
1!
1%
#110160000000
0!
0%
#110165000000
1!
1%
#110170000000
0!
0%
#110175000000
1!
1%
#110180000000
0!
0%
#110185000000
1!
1%
#110190000000
0!
0%
#110195000000
1!
1%
#110200000000
0!
0%
#110205000000
1!
1%
#110210000000
0!
0%
#110215000000
1!
1%
#110220000000
0!
0%
#110225000000
1!
1%
#110230000000
0!
0%
#110235000000
1!
1%
#110240000000
0!
0%
#110245000000
1!
1%
#110250000000
0!
0%
#110255000000
1!
1%
#110260000000
0!
0%
#110265000000
1!
1%
#110270000000
0!
0%
#110275000000
1!
1%
#110280000000
0!
0%
#110285000000
1!
1%
#110290000000
0!
0%
#110295000000
1!
1%
#110300000000
0!
0%
#110305000000
1!
1%
#110310000000
0!
0%
#110315000000
1!
1%
#110320000000
0!
0%
#110325000000
1!
1%
#110330000000
0!
0%
#110335000000
1!
1%
#110340000000
0!
0%
#110345000000
1!
1%
#110350000000
0!
0%
#110355000000
1!
1%
#110360000000
0!
0%
#110365000000
1!
1%
#110370000000
0!
0%
#110375000000
1!
1%
#110380000000
0!
0%
#110385000000
1!
1%
#110390000000
0!
0%
#110395000000
1!
1%
#110400000000
0!
0%
#110405000000
1!
1%
#110410000000
0!
0%
#110415000000
1!
1%
#110420000000
0!
0%
#110425000000
1!
1%
#110430000000
0!
0%
#110435000000
1!
1%
#110440000000
0!
0%
#110445000000
1!
1%
#110450000000
0!
0%
#110455000000
1!
1%
#110460000000
0!
0%
#110465000000
1!
1%
#110470000000
0!
0%
#110475000000
1!
1%
#110480000000
0!
0%
#110485000000
1!
1%
#110490000000
0!
0%
#110495000000
1!
1%
#110500000000
0!
0%
#110505000000
1!
1%
#110510000000
0!
0%
#110515000000
1!
1%
#110520000000
0!
0%
#110525000000
1!
1%
#110530000000
0!
0%
#110535000000
1!
1%
#110540000000
0!
0%
#110545000000
1!
1%
#110550000000
0!
0%
#110555000000
1!
1%
#110560000000
0!
0%
#110565000000
1!
1%
#110570000000
0!
0%
#110575000000
1!
1%
#110580000000
0!
0%
#110585000000
1!
1%
#110590000000
0!
0%
#110595000000
1!
1%
#110600000000
0!
0%
#110605000000
1!
1%
#110610000000
0!
0%
#110615000000
1!
1%
#110620000000
0!
0%
#110625000000
1!
1%
#110630000000
0!
0%
#110635000000
1!
1%
#110640000000
0!
0%
#110645000000
1!
1%
#110650000000
0!
0%
#110655000000
1!
1%
#110660000000
0!
0%
#110665000000
1!
1%
#110670000000
0!
0%
#110675000000
1!
1%
#110680000000
0!
0%
#110685000000
1!
1%
#110690000000
0!
0%
#110695000000
1!
1%
#110700000000
0!
0%
#110705000000
1!
1%
#110710000000
0!
0%
#110715000000
1!
1%
#110720000000
0!
0%
#110725000000
1!
1%
#110730000000
0!
0%
#110735000000
1!
1%
#110740000000
0!
0%
#110745000000
1!
1%
#110750000000
0!
0%
#110755000000
1!
1%
#110760000000
0!
0%
#110765000000
1!
1%
#110770000000
0!
0%
#110775000000
1!
1%
#110780000000
0!
0%
#110785000000
1!
1%
#110790000000
0!
0%
#110795000000
1!
1%
#110800000000
0!
0%
#110805000000
1!
1%
#110810000000
0!
0%
#110815000000
1!
1%
#110820000000
0!
0%
#110825000000
1!
1%
#110830000000
0!
0%
#110835000000
1!
1%
#110840000000
0!
0%
#110845000000
1!
1%
#110850000000
0!
0%
#110855000000
1!
1%
#110860000000
0!
0%
#110865000000
1!
1%
#110870000000
0!
0%
#110875000000
1!
1%
#110880000000
0!
0%
#110885000000
1!
1%
#110890000000
0!
0%
#110895000000
1!
1%
#110900000000
0!
0%
#110905000000
1!
1%
#110910000000
0!
0%
#110915000000
1!
1%
#110920000000
0!
0%
#110925000000
1!
1%
#110930000000
0!
0%
#110935000000
1!
1%
#110940000000
0!
0%
#110945000000
1!
1%
#110950000000
0!
0%
#110955000000
1!
1%
#110960000000
0!
0%
#110965000000
1!
1%
#110970000000
0!
0%
#110975000000
1!
1%
#110980000000
0!
0%
#110985000000
1!
1%
#110990000000
0!
0%
#110995000000
1!
1%
#111000000000
0!
0%
#111005000000
1!
1%
#111010000000
0!
0%
#111015000000
1!
1%
#111020000000
0!
0%
#111025000000
1!
1%
#111030000000
0!
0%
#111035000000
1!
1%
#111040000000
0!
0%
#111045000000
1!
1%
#111050000000
0!
0%
#111055000000
1!
1%
#111060000000
0!
0%
#111065000000
1!
1%
#111070000000
0!
0%
#111075000000
1!
1%
#111080000000
0!
0%
#111085000000
1!
1%
#111090000000
0!
0%
#111095000000
1!
1%
#111100000000
0!
0%
#111105000000
1!
1%
#111110000000
0!
0%
#111115000000
1!
1%
#111120000000
0!
0%
#111125000000
1!
1%
#111130000000
0!
0%
#111135000000
1!
1%
#111140000000
0!
0%
#111145000000
1!
1%
#111150000000
0!
0%
#111155000000
1!
1%
#111160000000
0!
0%
#111165000000
1!
1%
#111170000000
0!
0%
#111175000000
1!
1%
#111180000000
0!
0%
#111185000000
1!
1%
#111190000000
0!
0%
#111195000000
1!
1%
#111200000000
0!
0%
#111205000000
1!
1%
#111210000000
0!
0%
#111215000000
1!
1%
#111220000000
0!
0%
#111225000000
1!
1%
#111230000000
0!
0%
#111235000000
1!
1%
#111240000000
0!
0%
#111245000000
1!
1%
#111250000000
0!
0%
#111255000000
1!
1%
#111260000000
0!
0%
#111265000000
1!
1%
#111270000000
0!
0%
#111275000000
1!
1%
#111280000000
0!
0%
#111285000000
1!
1%
#111290000000
0!
0%
#111295000000
1!
1%
#111300000000
0!
0%
#111305000000
1!
1%
#111310000000
0!
0%
#111315000000
1!
1%
#111320000000
0!
0%
#111325000000
1!
1%
#111330000000
0!
0%
#111335000000
1!
1%
#111340000000
0!
0%
#111345000000
1!
1%
#111350000000
0!
0%
#111355000000
1!
1%
#111360000000
0!
0%
#111365000000
1!
1%
#111370000000
0!
0%
#111375000000
1!
1%
#111380000000
0!
0%
#111385000000
1!
1%
#111390000000
0!
0%
#111395000000
1!
1%
#111400000000
0!
0%
#111405000000
1!
1%
#111410000000
0!
0%
#111415000000
1!
1%
#111420000000
0!
0%
#111425000000
1!
1%
#111430000000
0!
0%
#111435000000
1!
1%
#111440000000
0!
0%
#111445000000
1!
1%
#111450000000
0!
0%
#111455000000
1!
1%
#111460000000
0!
0%
#111465000000
1!
1%
#111470000000
0!
0%
#111475000000
1!
1%
#111480000000
0!
0%
#111485000000
1!
1%
#111490000000
0!
0%
#111495000000
1!
1%
#111500000000
0!
0%
#111505000000
1!
1%
#111510000000
0!
0%
#111515000000
1!
1%
#111520000000
0!
0%
#111525000000
1!
1%
#111530000000
0!
0%
#111535000000
1!
1%
#111540000000
0!
0%
#111545000000
1!
1%
#111550000000
0!
0%
#111555000000
1!
1%
#111560000000
0!
0%
#111565000000
1!
1%
#111570000000
0!
0%
#111575000000
1!
1%
#111580000000
0!
0%
#111585000000
1!
1%
#111590000000
0!
0%
#111595000000
1!
1%
#111600000000
0!
0%
#111605000000
1!
1%
#111610000000
0!
0%
#111615000000
1!
1%
#111620000000
0!
0%
#111625000000
1!
1%
#111630000000
0!
0%
#111635000000
1!
1%
#111640000000
0!
0%
#111645000000
1!
1%
#111650000000
0!
0%
#111655000000
1!
1%
#111660000000
0!
0%
#111665000000
1!
1%
#111670000000
0!
0%
#111675000000
1!
1%
#111680000000
0!
0%
#111685000000
1!
1%
#111690000000
0!
0%
#111695000000
1!
1%
#111700000000
0!
0%
#111705000000
1!
1%
#111710000000
0!
0%
#111715000000
1!
1%
#111720000000
0!
0%
#111725000000
1!
1%
#111730000000
0!
0%
#111735000000
1!
1%
#111740000000
0!
0%
#111745000000
1!
1%
#111750000000
0!
0%
#111755000000
1!
1%
#111760000000
0!
0%
#111765000000
1!
1%
#111770000000
0!
0%
#111775000000
1!
1%
#111780000000
0!
0%
#111785000000
1!
1%
#111790000000
0!
0%
#111795000000
1!
1%
#111800000000
0!
0%
#111805000000
1!
1%
#111810000000
0!
0%
#111815000000
1!
1%
#111820000000
0!
0%
#111825000000
1!
1%
#111830000000
0!
0%
#111835000000
1!
1%
#111840000000
0!
0%
#111845000000
1!
1%
#111850000000
0!
0%
#111855000000
1!
1%
#111860000000
0!
0%
#111865000000
1!
1%
#111870000000
0!
0%
#111875000000
1!
1%
#111880000000
0!
0%
#111885000000
1!
1%
#111890000000
0!
0%
#111895000000
1!
1%
#111900000000
0!
0%
#111905000000
1!
1%
#111910000000
0!
0%
#111915000000
1!
1%
#111920000000
0!
0%
#111925000000
1!
1%
#111930000000
0!
0%
#111935000000
1!
1%
#111940000000
0!
0%
#111945000000
1!
1%
#111950000000
0!
0%
#111955000000
1!
1%
#111960000000
0!
0%
#111965000000
1!
1%
#111970000000
0!
0%
#111975000000
1!
1%
#111980000000
0!
0%
#111985000000
1!
1%
#111990000000
0!
0%
#111995000000
1!
1%
#112000000000
0!
0%
#112005000000
1!
1%
#112010000000
0!
0%
#112015000000
1!
1%
#112020000000
0!
0%
#112025000000
1!
1%
#112030000000
0!
0%
#112035000000
1!
1%
#112040000000
0!
0%
#112045000000
1!
1%
#112050000000
0!
0%
#112055000000
1!
1%
#112060000000
0!
0%
#112065000000
1!
1%
#112070000000
0!
0%
#112075000000
1!
1%
#112080000000
0!
0%
#112085000000
1!
1%
#112090000000
0!
0%
#112095000000
1!
1%
#112100000000
0!
0%
#112105000000
1!
1%
#112110000000
0!
0%
#112115000000
1!
1%
#112120000000
0!
0%
#112125000000
1!
1%
#112130000000
0!
0%
#112135000000
1!
1%
#112140000000
0!
0%
#112145000000
1!
1%
#112150000000
0!
0%
#112155000000
1!
1%
#112160000000
0!
0%
#112165000000
1!
1%
#112170000000
0!
0%
#112175000000
1!
1%
#112180000000
0!
0%
#112185000000
1!
1%
#112190000000
0!
0%
#112195000000
1!
1%
#112200000000
0!
0%
#112205000000
1!
1%
#112210000000
0!
0%
#112215000000
1!
1%
#112220000000
0!
0%
#112225000000
1!
1%
#112230000000
0!
0%
#112235000000
1!
1%
#112240000000
0!
0%
#112245000000
1!
1%
#112250000000
0!
0%
#112255000000
1!
1%
#112260000000
0!
0%
#112265000000
1!
1%
#112270000000
0!
0%
#112275000000
1!
1%
#112280000000
0!
0%
#112285000000
1!
1%
#112290000000
0!
0%
#112295000000
1!
1%
#112300000000
0!
0%
#112305000000
1!
1%
#112310000000
0!
0%
#112315000000
1!
1%
#112320000000
0!
0%
#112325000000
1!
1%
#112330000000
0!
0%
#112335000000
1!
1%
#112340000000
0!
0%
#112345000000
1!
1%
#112350000000
0!
0%
#112355000000
1!
1%
#112360000000
0!
0%
#112365000000
1!
1%
#112370000000
0!
0%
#112375000000
1!
1%
#112380000000
0!
0%
#112385000000
1!
1%
#112390000000
0!
0%
#112395000000
1!
1%
#112400000000
0!
0%
#112405000000
1!
1%
#112410000000
0!
0%
#112415000000
1!
1%
#112420000000
0!
0%
#112425000000
1!
1%
#112430000000
0!
0%
#112435000000
1!
1%
#112440000000
0!
0%
#112445000000
1!
1%
#112450000000
0!
0%
#112455000000
1!
1%
#112460000000
0!
0%
#112465000000
1!
1%
#112470000000
0!
0%
#112475000000
1!
1%
#112480000000
0!
0%
#112485000000
1!
1%
#112490000000
0!
0%
#112495000000
1!
1%
#112500000000
0!
0%
#112505000000
1!
1%
#112510000000
0!
0%
#112515000000
1!
1%
#112520000000
0!
0%
#112525000000
1!
1%
#112530000000
0!
0%
#112535000000
1!
1%
#112540000000
0!
0%
#112545000000
1!
1%
#112550000000
0!
0%
#112555000000
1!
1%
#112560000000
0!
0%
#112565000000
1!
1%
#112570000000
0!
0%
#112575000000
1!
1%
#112580000000
0!
0%
#112585000000
1!
1%
#112590000000
0!
0%
#112595000000
1!
1%
#112600000000
0!
0%
#112605000000
1!
1%
#112610000000
0!
0%
#112615000000
1!
1%
#112620000000
0!
0%
#112625000000
1!
1%
#112630000000
0!
0%
#112635000000
1!
1%
#112640000000
0!
0%
#112645000000
1!
1%
#112650000000
0!
0%
#112655000000
1!
1%
#112660000000
0!
0%
#112665000000
1!
1%
#112670000000
0!
0%
#112675000000
1!
1%
#112680000000
0!
0%
#112685000000
1!
1%
#112690000000
0!
0%
#112695000000
1!
1%
#112700000000
0!
0%
#112705000000
1!
1%
#112710000000
0!
0%
#112715000000
1!
1%
#112720000000
0!
0%
#112725000000
1!
1%
#112730000000
0!
0%
#112735000000
1!
1%
#112740000000
0!
0%
#112745000000
1!
1%
#112750000000
0!
0%
#112755000000
1!
1%
#112760000000
0!
0%
#112765000000
1!
1%
#112770000000
0!
0%
#112775000000
1!
1%
#112780000000
0!
0%
#112785000000
1!
1%
#112790000000
0!
0%
#112795000000
1!
1%
#112800000000
0!
0%
#112805000000
1!
1%
#112810000000
0!
0%
#112815000000
1!
1%
#112820000000
0!
0%
#112825000000
1!
1%
#112830000000
0!
0%
#112835000000
1!
1%
#112840000000
0!
0%
#112845000000
1!
1%
#112850000000
0!
0%
#112855000000
1!
1%
#112860000000
0!
0%
#112865000000
1!
1%
#112870000000
0!
0%
#112875000000
1!
1%
#112880000000
0!
0%
#112885000000
1!
1%
#112890000000
0!
0%
#112895000000
1!
1%
#112900000000
0!
0%
#112905000000
1!
1%
#112910000000
0!
0%
#112915000000
1!
1%
#112920000000
0!
0%
#112925000000
1!
1%
#112930000000
0!
0%
#112935000000
1!
1%
#112940000000
0!
0%
#112945000000
1!
1%
#112950000000
0!
0%
#112955000000
1!
1%
#112960000000
0!
0%
#112965000000
1!
1%
#112970000000
0!
0%
#112975000000
1!
1%
#112980000000
0!
0%
#112985000000
1!
1%
#112990000000
0!
0%
#112995000000
1!
1%
#113000000000
0!
0%
#113005000000
1!
1%
#113010000000
0!
0%
#113015000000
1!
1%
#113020000000
0!
0%
#113025000000
1!
1%
#113030000000
0!
0%
#113035000000
1!
1%
#113040000000
0!
0%
#113045000000
1!
1%
#113050000000
0!
0%
#113055000000
1!
1%
#113060000000
0!
0%
#113065000000
1!
1%
#113070000000
0!
0%
#113075000000
1!
1%
#113080000000
0!
0%
#113085000000
1!
1%
#113090000000
0!
0%
#113095000000
1!
1%
#113100000000
0!
0%
#113105000000
1!
1%
#113110000000
0!
0%
#113115000000
1!
1%
#113120000000
0!
0%
#113125000000
1!
1%
#113130000000
0!
0%
#113135000000
1!
1%
#113140000000
0!
0%
#113145000000
1!
1%
#113150000000
0!
0%
#113155000000
1!
1%
#113160000000
0!
0%
#113165000000
1!
1%
#113170000000
0!
0%
#113175000000
1!
1%
#113180000000
0!
0%
#113185000000
1!
1%
#113190000000
0!
0%
#113195000000
1!
1%
#113200000000
0!
0%
#113205000000
1!
1%
#113210000000
0!
0%
#113215000000
1!
1%
#113220000000
0!
0%
#113225000000
1!
1%
#113230000000
0!
0%
#113235000000
1!
1%
#113240000000
0!
0%
#113245000000
1!
1%
#113250000000
0!
0%
#113255000000
1!
1%
#113260000000
0!
0%
#113265000000
1!
1%
#113270000000
0!
0%
#113275000000
1!
1%
#113280000000
0!
0%
#113285000000
1!
1%
#113290000000
0!
0%
#113295000000
1!
1%
#113300000000
0!
0%
#113305000000
1!
1%
#113310000000
0!
0%
#113315000000
1!
1%
#113320000000
0!
0%
#113325000000
1!
1%
#113330000000
0!
0%
#113335000000
1!
1%
#113340000000
0!
0%
#113345000000
1!
1%
#113350000000
0!
0%
#113355000000
1!
1%
#113360000000
0!
0%
#113365000000
1!
1%
#113370000000
0!
0%
#113375000000
1!
1%
#113380000000
0!
0%
#113385000000
1!
1%
#113390000000
0!
0%
#113395000000
1!
1%
#113400000000
0!
0%
#113405000000
1!
1%
#113410000000
0!
0%
#113415000000
1!
1%
#113420000000
0!
0%
#113425000000
1!
1%
#113430000000
0!
0%
#113435000000
1!
1%
#113440000000
0!
0%
#113445000000
1!
1%
#113450000000
0!
0%
#113455000000
1!
1%
#113460000000
0!
0%
#113465000000
1!
1%
#113470000000
0!
0%
#113475000000
1!
1%
#113480000000
0!
0%
#113485000000
1!
1%
#113490000000
0!
0%
#113495000000
1!
1%
#113500000000
0!
0%
#113505000000
1!
1%
#113510000000
0!
0%
#113515000000
1!
1%
#113520000000
0!
0%
#113525000000
1!
1%
#113530000000
0!
0%
#113535000000
1!
1%
#113540000000
0!
0%
#113545000000
1!
1%
#113550000000
0!
0%
#113555000000
1!
1%
#113560000000
0!
0%
#113565000000
1!
1%
#113570000000
0!
0%
#113575000000
1!
1%
#113580000000
0!
0%
#113585000000
1!
1%
#113590000000
0!
0%
#113595000000
1!
1%
#113600000000
0!
0%
#113605000000
1!
1%
#113610000000
0!
0%
#113615000000
1!
1%
#113620000000
0!
0%
#113625000000
1!
1%
#113630000000
0!
0%
#113635000000
1!
1%
#113640000000
0!
0%
#113645000000
1!
1%
#113650000000
0!
0%
#113655000000
1!
1%
#113660000000
0!
0%
#113665000000
1!
1%
#113670000000
0!
0%
#113675000000
1!
1%
#113680000000
0!
0%
#113685000000
1!
1%
#113690000000
0!
0%
#113695000000
1!
1%
#113700000000
0!
0%
#113705000000
1!
1%
#113710000000
0!
0%
#113715000000
1!
1%
#113720000000
0!
0%
#113725000000
1!
1%
#113730000000
0!
0%
#113735000000
1!
1%
#113740000000
0!
0%
#113745000000
1!
1%
#113750000000
0!
0%
#113755000000
1!
1%
#113760000000
0!
0%
#113765000000
1!
1%
#113770000000
0!
0%
#113775000000
1!
1%
#113780000000
0!
0%
#113785000000
1!
1%
#113790000000
0!
0%
#113795000000
1!
1%
#113800000000
0!
0%
#113805000000
1!
1%
#113810000000
0!
0%
#113815000000
1!
1%
#113820000000
0!
0%
#113825000000
1!
1%
#113830000000
0!
0%
#113835000000
1!
1%
#113840000000
0!
0%
#113845000000
1!
1%
#113850000000
0!
0%
#113855000000
1!
1%
#113860000000
0!
0%
#113865000000
1!
1%
#113870000000
0!
0%
#113875000000
1!
1%
#113880000000
0!
0%
#113885000000
1!
1%
#113890000000
0!
0%
#113895000000
1!
1%
#113900000000
0!
0%
#113905000000
1!
1%
#113910000000
0!
0%
#113915000000
1!
1%
#113920000000
0!
0%
#113925000000
1!
1%
#113930000000
0!
0%
#113935000000
1!
1%
#113940000000
0!
0%
#113945000000
1!
1%
#113950000000
0!
0%
#113955000000
1!
1%
#113960000000
0!
0%
#113965000000
1!
1%
#113970000000
0!
0%
#113975000000
1!
1%
#113980000000
0!
0%
#113985000000
1!
1%
#113990000000
0!
0%
#113995000000
1!
1%
#114000000000
0!
0%
#114005000000
1!
1%
#114010000000
0!
0%
#114015000000
1!
1%
#114020000000
0!
0%
#114025000000
1!
1%
#114030000000
0!
0%
#114035000000
1!
1%
#114040000000
0!
0%
#114045000000
1!
1%
#114050000000
0!
0%
#114055000000
1!
1%
#114060000000
0!
0%
#114065000000
1!
1%
#114070000000
0!
0%
#114075000000
1!
1%
#114080000000
0!
0%
#114085000000
1!
1%
#114090000000
0!
0%
#114095000000
1!
1%
#114100000000
0!
0%
#114105000000
1!
1%
#114110000000
0!
0%
#114115000000
1!
1%
#114120000000
0!
0%
#114125000000
1!
1%
#114130000000
0!
0%
#114135000000
1!
1%
#114140000000
0!
0%
#114145000000
1!
1%
#114150000000
0!
0%
#114155000000
1!
1%
#114160000000
0!
0%
#114165000000
1!
1%
#114170000000
0!
0%
#114175000000
1!
1%
#114180000000
0!
0%
#114185000000
1!
1%
#114190000000
0!
0%
#114195000000
1!
1%
#114200000000
0!
0%
#114205000000
1!
1%
#114210000000
0!
0%
#114215000000
1!
1%
#114220000000
0!
0%
#114225000000
1!
1%
#114230000000
0!
0%
#114235000000
1!
1%
#114240000000
0!
0%
#114245000000
1!
1%
#114250000000
0!
0%
#114255000000
1!
1%
#114260000000
0!
0%
#114265000000
1!
1%
#114270000000
0!
0%
#114275000000
1!
1%
#114280000000
0!
0%
#114285000000
1!
1%
#114290000000
0!
0%
#114295000000
1!
1%
#114300000000
0!
0%
#114305000000
1!
1%
#114310000000
0!
0%
#114315000000
1!
1%
#114320000000
0!
0%
#114325000000
1!
1%
#114330000000
0!
0%
#114335000000
1!
1%
#114340000000
0!
0%
#114345000000
1!
1%
#114350000000
0!
0%
#114355000000
1!
1%
#114360000000
0!
0%
#114365000000
1!
1%
#114370000000
0!
0%
#114375000000
1!
1%
#114380000000
0!
0%
#114385000000
1!
1%
#114390000000
0!
0%
#114395000000
1!
1%
#114400000000
0!
0%
#114405000000
1!
1%
#114410000000
0!
0%
#114415000000
1!
1%
#114420000000
0!
0%
#114425000000
1!
1%
#114430000000
0!
0%
#114435000000
1!
1%
#114440000000
0!
0%
#114445000000
1!
1%
#114450000000
0!
0%
#114455000000
1!
1%
#114460000000
0!
0%
#114465000000
1!
1%
#114470000000
0!
0%
#114475000000
1!
1%
#114480000000
0!
0%
#114485000000
1!
1%
#114490000000
0!
0%
#114495000000
1!
1%
#114500000000
0!
0%
#114505000000
1!
1%
#114510000000
0!
0%
#114515000000
1!
1%
#114520000000
0!
0%
#114525000000
1!
1%
#114530000000
0!
0%
#114535000000
1!
1%
#114540000000
0!
0%
#114545000000
1!
1%
#114550000000
0!
0%
#114555000000
1!
1%
#114560000000
0!
0%
#114565000000
1!
1%
#114570000000
0!
0%
#114575000000
1!
1%
#114580000000
0!
0%
#114585000000
1!
1%
#114590000000
0!
0%
#114595000000
1!
1%
#114600000000
0!
0%
#114605000000
1!
1%
#114610000000
0!
0%
#114615000000
1!
1%
#114620000000
0!
0%
#114625000000
1!
1%
#114630000000
0!
0%
#114635000000
1!
1%
#114640000000
0!
0%
#114645000000
1!
1%
#114650000000
0!
0%
#114655000000
1!
1%
#114660000000
0!
0%
#114665000000
1!
1%
#114670000000
0!
0%
#114675000000
1!
1%
#114680000000
0!
0%
#114685000000
1!
1%
#114690000000
0!
0%
#114695000000
1!
1%
#114700000000
0!
0%
#114705000000
1!
1%
#114710000000
0!
0%
#114715000000
1!
1%
#114720000000
0!
0%
#114725000000
1!
1%
#114730000000
0!
0%
#114735000000
1!
1%
#114740000000
0!
0%
#114745000000
1!
1%
#114750000000
0!
0%
#114755000000
1!
1%
#114760000000
0!
0%
#114765000000
1!
1%
#114770000000
0!
0%
#114775000000
1!
1%
#114780000000
0!
0%
#114785000000
1!
1%
#114790000000
0!
0%
#114795000000
1!
1%
#114800000000
0!
0%
#114805000000
1!
1%
#114810000000
0!
0%
#114815000000
1!
1%
#114820000000
0!
0%
#114825000000
1!
1%
#114830000000
0!
0%
#114835000000
1!
1%
#114840000000
0!
0%
#114845000000
1!
1%
#114850000000
0!
0%
#114855000000
1!
1%
#114860000000
0!
0%
#114865000000
1!
1%
#114870000000
0!
0%
#114875000000
1!
1%
#114880000000
0!
0%
#114885000000
1!
1%
#114890000000
0!
0%
#114895000000
1!
1%
#114900000000
0!
0%
#114905000000
1!
1%
#114910000000
0!
0%
#114915000000
1!
1%
#114920000000
0!
0%
#114925000000
1!
1%
#114930000000
0!
0%
#114935000000
1!
1%
#114940000000
0!
0%
#114945000000
1!
1%
#114950000000
0!
0%
#114955000000
1!
1%
#114960000000
0!
0%
#114965000000
1!
1%
#114970000000
0!
0%
#114975000000
1!
1%
#114980000000
0!
0%
#114985000000
1!
1%
#114990000000
0!
0%
#114995000000
1!
1%
#115000000000
0!
0%
#115005000000
1!
1%
#115010000000
0!
0%
#115015000000
1!
1%
#115020000000
0!
0%
#115025000000
1!
1%
#115030000000
0!
0%
#115035000000
1!
1%
#115040000000
0!
0%
#115045000000
1!
1%
#115050000000
0!
0%
#115055000000
1!
1%
#115060000000
0!
0%
#115065000000
1!
1%
#115070000000
0!
0%
#115075000000
1!
1%
#115080000000
0!
0%
#115085000000
1!
1%
#115090000000
0!
0%
#115095000000
1!
1%
#115100000000
0!
0%
#115105000000
1!
1%
#115110000000
0!
0%
#115115000000
1!
1%
#115120000000
0!
0%
#115125000000
1!
1%
#115130000000
0!
0%
#115135000000
1!
1%
#115140000000
0!
0%
#115145000000
1!
1%
#115150000000
0!
0%
#115155000000
1!
1%
#115160000000
0!
0%
#115165000000
1!
1%
#115170000000
0!
0%
#115175000000
1!
1%
#115180000000
0!
0%
#115185000000
1!
1%
#115190000000
0!
0%
#115195000000
1!
1%
#115200000000
0!
0%
#115205000000
1!
1%
#115210000000
0!
0%
#115215000000
1!
1%
#115220000000
0!
0%
#115225000000
1!
1%
#115230000000
0!
0%
#115235000000
1!
1%
#115240000000
0!
0%
#115245000000
1!
1%
#115250000000
0!
0%
#115255000000
1!
1%
#115260000000
0!
0%
#115265000000
1!
1%
#115270000000
0!
0%
#115275000000
1!
1%
#115280000000
0!
0%
#115285000000
1!
1%
#115290000000
0!
0%
#115295000000
1!
1%
#115300000000
0!
0%
#115305000000
1!
1%
#115310000000
0!
0%
#115315000000
1!
1%
#115320000000
0!
0%
#115325000000
1!
1%
#115330000000
0!
0%
#115335000000
1!
1%
#115340000000
0!
0%
#115345000000
1!
1%
#115350000000
0!
0%
#115355000000
1!
1%
#115360000000
0!
0%
#115365000000
1!
1%
#115370000000
0!
0%
#115375000000
1!
1%
#115380000000
0!
0%
#115385000000
1!
1%
#115390000000
0!
0%
#115395000000
1!
1%
#115400000000
0!
0%
#115405000000
1!
1%
#115410000000
0!
0%
#115415000000
1!
1%
#115420000000
0!
0%
#115425000000
1!
1%
#115430000000
0!
0%
#115435000000
1!
1%
#115440000000
0!
0%
#115445000000
1!
1%
#115450000000
0!
0%
#115455000000
1!
1%
#115460000000
0!
0%
#115465000000
1!
1%
#115470000000
0!
0%
#115475000000
1!
1%
#115480000000
0!
0%
#115485000000
1!
1%
#115490000000
0!
0%
#115495000000
1!
1%
#115500000000
0!
0%
#115505000000
1!
1%
#115510000000
0!
0%
#115515000000
1!
1%
#115520000000
0!
0%
#115525000000
1!
1%
#115530000000
0!
0%
#115535000000
1!
1%
#115540000000
0!
0%
#115545000000
1!
1%
#115550000000
0!
0%
#115555000000
1!
1%
#115560000000
0!
0%
#115565000000
1!
1%
#115570000000
0!
0%
#115575000000
1!
1%
#115580000000
0!
0%
#115585000000
1!
1%
#115590000000
0!
0%
#115595000000
1!
1%
#115600000000
0!
0%
#115605000000
1!
1%
#115610000000
0!
0%
#115615000000
1!
1%
#115620000000
0!
0%
#115625000000
1!
1%
#115630000000
0!
0%
#115635000000
1!
1%
#115640000000
0!
0%
#115645000000
1!
1%
#115650000000
0!
0%
#115655000000
1!
1%
#115660000000
0!
0%
#115665000000
1!
1%
#115670000000
0!
0%
#115675000000
1!
1%
#115680000000
0!
0%
#115685000000
1!
1%
#115690000000
0!
0%
#115695000000
1!
1%
#115700000000
0!
0%
#115705000000
1!
1%
#115710000000
0!
0%
#115715000000
1!
1%
#115720000000
0!
0%
#115725000000
1!
1%
#115730000000
0!
0%
#115735000000
1!
1%
#115740000000
0!
0%
#115745000000
1!
1%
#115750000000
0!
0%
#115755000000
1!
1%
#115760000000
0!
0%
#115765000000
1!
1%
#115770000000
0!
0%
#115775000000
1!
1%
#115780000000
0!
0%
#115785000000
1!
1%
#115790000000
0!
0%
#115795000000
1!
1%
#115800000000
0!
0%
#115805000000
1!
1%
#115810000000
0!
0%
#115815000000
1!
1%
#115820000000
0!
0%
#115825000000
1!
1%
#115830000000
0!
0%
#115835000000
1!
1%
#115840000000
0!
0%
#115845000000
1!
1%
#115850000000
0!
0%
#115855000000
1!
1%
#115860000000
0!
0%
#115865000000
1!
1%
#115870000000
0!
0%
#115875000000
1!
1%
#115880000000
0!
0%
#115885000000
1!
1%
#115890000000
0!
0%
#115895000000
1!
1%
#115900000000
0!
0%
#115905000000
1!
1%
#115910000000
0!
0%
#115915000000
1!
1%
#115920000000
0!
0%
#115925000000
1!
1%
#115930000000
0!
0%
#115935000000
1!
1%
#115940000000
0!
0%
#115945000000
1!
1%
#115950000000
0!
0%
#115955000000
1!
1%
#115960000000
0!
0%
#115965000000
1!
1%
#115970000000
0!
0%
#115975000000
1!
1%
#115980000000
0!
0%
#115985000000
1!
1%
#115990000000
0!
0%
#115995000000
1!
1%
#116000000000
0!
0%
#116005000000
1!
1%
#116010000000
0!
0%
#116015000000
1!
1%
#116020000000
0!
0%
#116025000000
1!
1%
#116030000000
0!
0%
#116035000000
1!
1%
#116040000000
0!
0%
#116045000000
1!
1%
#116050000000
0!
0%
#116055000000
1!
1%
#116060000000
0!
0%
#116065000000
1!
1%
#116070000000
0!
0%
#116075000000
1!
1%
#116080000000
0!
0%
#116085000000
1!
1%
#116090000000
0!
0%
#116095000000
1!
1%
#116100000000
0!
0%
#116105000000
1!
1%
#116110000000
0!
0%
#116115000000
1!
1%
#116120000000
0!
0%
#116125000000
1!
1%
#116130000000
0!
0%
#116135000000
1!
1%
#116140000000
0!
0%
#116145000000
1!
1%
#116150000000
0!
0%
#116155000000
1!
1%
#116160000000
0!
0%
#116165000000
1!
1%
#116170000000
0!
0%
#116175000000
1!
1%
#116180000000
0!
0%
#116185000000
1!
1%
#116190000000
0!
0%
#116195000000
1!
1%
#116200000000
0!
0%
#116205000000
1!
1%
#116210000000
0!
0%
#116215000000
1!
1%
#116220000000
0!
0%
#116225000000
1!
1%
#116230000000
0!
0%
#116235000000
1!
1%
#116240000000
0!
0%
#116245000000
1!
1%
#116250000000
0!
0%
#116255000000
1!
1%
#116260000000
0!
0%
#116265000000
1!
1%
#116270000000
0!
0%
#116275000000
1!
1%
#116280000000
0!
0%
#116285000000
1!
1%
#116290000000
0!
0%
#116295000000
1!
1%
#116300000000
0!
0%
#116305000000
1!
1%
#116310000000
0!
0%
#116315000000
1!
1%
#116320000000
0!
0%
#116325000000
1!
1%
#116330000000
0!
0%
#116335000000
1!
1%
#116340000000
0!
0%
#116345000000
1!
1%
#116350000000
0!
0%
#116355000000
1!
1%
#116360000000
0!
0%
#116365000000
1!
1%
#116370000000
0!
0%
#116375000000
1!
1%
#116380000000
0!
0%
#116385000000
1!
1%
#116390000000
0!
0%
#116395000000
1!
1%
#116400000000
0!
0%
#116405000000
1!
1%
#116410000000
0!
0%
#116415000000
1!
1%
#116420000000
0!
0%
#116425000000
1!
1%
#116430000000
0!
0%
#116435000000
1!
1%
#116440000000
0!
0%
#116445000000
1!
1%
#116450000000
0!
0%
#116455000000
1!
1%
#116460000000
0!
0%
#116465000000
1!
1%
#116470000000
0!
0%
#116475000000
1!
1%
#116480000000
0!
0%
#116485000000
1!
1%
#116490000000
0!
0%
#116495000000
1!
1%
#116500000000
0!
0%
#116505000000
1!
1%
#116510000000
0!
0%
#116515000000
1!
1%
#116520000000
0!
0%
#116525000000
1!
1%
#116530000000
0!
0%
#116535000000
1!
1%
#116540000000
0!
0%
#116545000000
1!
1%
#116550000000
0!
0%
#116555000000
1!
1%
#116560000000
0!
0%
#116565000000
1!
1%
#116570000000
0!
0%
#116575000000
1!
1%
#116580000000
0!
0%
#116585000000
1!
1%
#116590000000
0!
0%
#116595000000
1!
1%
#116600000000
0!
0%
#116605000000
1!
1%
#116610000000
0!
0%
#116615000000
1!
1%
#116620000000
0!
0%
#116625000000
1!
1%
#116630000000
0!
0%
#116635000000
1!
1%
#116640000000
0!
0%
#116645000000
1!
1%
#116650000000
0!
0%
#116655000000
1!
1%
#116660000000
0!
0%
#116665000000
1!
1%
#116670000000
0!
0%
#116675000000
1!
1%
#116680000000
0!
0%
#116685000000
1!
1%
#116690000000
0!
0%
#116695000000
1!
1%
#116700000000
0!
0%
#116705000000
1!
1%
#116710000000
0!
0%
#116715000000
1!
1%
#116720000000
0!
0%
#116725000000
1!
1%
#116730000000
0!
0%
#116735000000
1!
1%
#116740000000
0!
0%
#116745000000
1!
1%
#116750000000
0!
0%
#116755000000
1!
1%
#116760000000
0!
0%
#116765000000
1!
1%
#116770000000
0!
0%
#116775000000
1!
1%
#116780000000
0!
0%
#116785000000
1!
1%
#116790000000
0!
0%
#116795000000
1!
1%
#116800000000
0!
0%
#116805000000
1!
1%
#116810000000
0!
0%
#116815000000
1!
1%
#116820000000
0!
0%
#116825000000
1!
1%
#116830000000
0!
0%
#116835000000
1!
1%
#116840000000
0!
0%
#116845000000
1!
1%
#116850000000
0!
0%
#116855000000
1!
1%
#116860000000
0!
0%
#116865000000
1!
1%
#116870000000
0!
0%
#116875000000
1!
1%
#116880000000
0!
0%
#116885000000
1!
1%
#116890000000
0!
0%
#116895000000
1!
1%
#116900000000
0!
0%
#116905000000
1!
1%
#116910000000
0!
0%
#116915000000
1!
1%
#116920000000
0!
0%
#116925000000
1!
1%
#116930000000
0!
0%
#116935000000
1!
1%
#116940000000
0!
0%
#116945000000
1!
1%
#116950000000
0!
0%
#116955000000
1!
1%
#116960000000
0!
0%
#116965000000
1!
1%
#116970000000
0!
0%
#116975000000
1!
1%
#116980000000
0!
0%
#116985000000
1!
1%
#116990000000
0!
0%
#116995000000
1!
1%
#117000000000
0!
0%
#117005000000
1!
1%
#117010000000
0!
0%
#117015000000
1!
1%
#117020000000
0!
0%
#117025000000
1!
1%
#117030000000
0!
0%
#117035000000
1!
1%
#117040000000
0!
0%
#117045000000
1!
1%
#117050000000
0!
0%
#117055000000
1!
1%
#117060000000
0!
0%
#117065000000
1!
1%
#117070000000
0!
0%
#117075000000
1!
1%
#117080000000
0!
0%
#117085000000
1!
1%
#117090000000
0!
0%
#117095000000
1!
1%
#117100000000
0!
0%
#117105000000
1!
1%
#117110000000
0!
0%
#117115000000
1!
1%
#117120000000
0!
0%
#117125000000
1!
1%
#117130000000
0!
0%
#117135000000
1!
1%
#117140000000
0!
0%
#117145000000
1!
1%
#117150000000
0!
0%
#117155000000
1!
1%
#117160000000
0!
0%
#117165000000
1!
1%
#117170000000
0!
0%
#117175000000
1!
1%
#117180000000
0!
0%
#117185000000
1!
1%
#117190000000
0!
0%
#117195000000
1!
1%
#117200000000
0!
0%
#117205000000
1!
1%
#117210000000
0!
0%
#117215000000
1!
1%
#117220000000
0!
0%
#117225000000
1!
1%
#117230000000
0!
0%
#117235000000
1!
1%
#117240000000
0!
0%
#117245000000
1!
1%
#117250000000
0!
0%
#117255000000
1!
1%
#117260000000
0!
0%
#117265000000
1!
1%
#117270000000
0!
0%
#117275000000
1!
1%
#117280000000
0!
0%
#117285000000
1!
1%
#117290000000
0!
0%
#117295000000
1!
1%
#117300000000
0!
0%
#117305000000
1!
1%
#117310000000
0!
0%
#117315000000
1!
1%
#117320000000
0!
0%
#117325000000
1!
1%
#117330000000
0!
0%
#117335000000
1!
1%
#117340000000
0!
0%
#117345000000
1!
1%
#117350000000
0!
0%
#117355000000
1!
1%
#117360000000
0!
0%
#117365000000
1!
1%
#117370000000
0!
0%
#117375000000
1!
1%
#117380000000
0!
0%
#117385000000
1!
1%
#117390000000
0!
0%
#117395000000
1!
1%
#117400000000
0!
0%
#117405000000
1!
1%
#117410000000
0!
0%
#117415000000
1!
1%
#117420000000
0!
0%
#117425000000
1!
1%
#117430000000
0!
0%
#117435000000
1!
1%
#117440000000
0!
0%
#117445000000
1!
1%
#117450000000
0!
0%
#117455000000
1!
1%
#117460000000
0!
0%
#117465000000
1!
1%
#117470000000
0!
0%
#117475000000
1!
1%
#117480000000
0!
0%
#117485000000
1!
1%
#117490000000
0!
0%
#117495000000
1!
1%
#117500000000
0!
0%
#117505000000
1!
1%
#117510000000
0!
0%
#117515000000
1!
1%
#117520000000
0!
0%
#117525000000
1!
1%
#117530000000
0!
0%
#117535000000
1!
1%
#117540000000
0!
0%
#117545000000
1!
1%
#117550000000
0!
0%
#117555000000
1!
1%
#117560000000
0!
0%
#117565000000
1!
1%
#117570000000
0!
0%
#117575000000
1!
1%
#117580000000
0!
0%
#117585000000
1!
1%
#117590000000
0!
0%
#117595000000
1!
1%
#117600000000
0!
0%
#117605000000
1!
1%
#117610000000
0!
0%
#117615000000
1!
1%
#117620000000
0!
0%
#117625000000
1!
1%
#117630000000
0!
0%
#117635000000
1!
1%
#117640000000
0!
0%
#117645000000
1!
1%
#117650000000
0!
0%
#117655000000
1!
1%
#117660000000
0!
0%
#117665000000
1!
1%
#117670000000
0!
0%
#117675000000
1!
1%
#117680000000
0!
0%
#117685000000
1!
1%
#117690000000
0!
0%
#117695000000
1!
1%
#117700000000
0!
0%
#117705000000
1!
1%
#117710000000
0!
0%
#117715000000
1!
1%
#117720000000
0!
0%
#117725000000
1!
1%
#117730000000
0!
0%
#117735000000
1!
1%
#117740000000
0!
0%
#117745000000
1!
1%
#117750000000
0!
0%
#117755000000
1!
1%
#117760000000
0!
0%
#117765000000
1!
1%
#117770000000
0!
0%
#117775000000
1!
1%
#117780000000
0!
0%
#117785000000
1!
1%
#117790000000
0!
0%
#117795000000
1!
1%
#117800000000
0!
0%
#117805000000
1!
1%
#117810000000
0!
0%
#117815000000
1!
1%
#117820000000
0!
0%
#117825000000
1!
1%
#117830000000
0!
0%
#117835000000
1!
1%
#117840000000
0!
0%
#117845000000
1!
1%
#117850000000
0!
0%
#117855000000
1!
1%
#117860000000
0!
0%
#117865000000
1!
1%
#117870000000
0!
0%
#117875000000
1!
1%
#117880000000
0!
0%
#117885000000
1!
1%
#117890000000
0!
0%
#117895000000
1!
1%
#117900000000
0!
0%
#117905000000
1!
1%
#117910000000
0!
0%
#117915000000
1!
1%
#117920000000
0!
0%
#117925000000
1!
1%
#117930000000
0!
0%
#117935000000
1!
1%
#117940000000
0!
0%
#117945000000
1!
1%
#117950000000
0!
0%
#117955000000
1!
1%
#117960000000
0!
0%
#117965000000
1!
1%
#117970000000
0!
0%
#117975000000
1!
1%
#117980000000
0!
0%
#117985000000
1!
1%
#117990000000
0!
0%
#117995000000
1!
1%
#118000000000
0!
0%
#118005000000
1!
1%
#118010000000
0!
0%
#118015000000
1!
1%
#118020000000
0!
0%
#118025000000
1!
1%
#118030000000
0!
0%
#118035000000
1!
1%
#118040000000
0!
0%
#118045000000
1!
1%
#118050000000
0!
0%
#118055000000
1!
1%
#118060000000
0!
0%
#118065000000
1!
1%
#118070000000
0!
0%
#118075000000
1!
1%
#118080000000
0!
0%
#118085000000
1!
1%
#118090000000
0!
0%
#118095000000
1!
1%
#118100000000
0!
0%
#118105000000
1!
1%
#118110000000
0!
0%
#118115000000
1!
1%
#118120000000
0!
0%
#118125000000
1!
1%
#118130000000
0!
0%
#118135000000
1!
1%
#118140000000
0!
0%
#118145000000
1!
1%
#118150000000
0!
0%
#118155000000
1!
1%
#118160000000
0!
0%
#118165000000
1!
1%
#118170000000
0!
0%
#118175000000
1!
1%
#118180000000
0!
0%
#118185000000
1!
1%
#118190000000
0!
0%
#118195000000
1!
1%
#118200000000
0!
0%
#118205000000
1!
1%
#118210000000
0!
0%
#118215000000
1!
1%
#118220000000
0!
0%
#118225000000
1!
1%
#118230000000
0!
0%
#118235000000
1!
1%
#118240000000
0!
0%
#118245000000
1!
1%
#118250000000
0!
0%
#118255000000
1!
1%
#118260000000
0!
0%
#118265000000
1!
1%
#118270000000
0!
0%
#118275000000
1!
1%
#118280000000
0!
0%
#118285000000
1!
1%
#118290000000
0!
0%
#118295000000
1!
1%
#118300000000
0!
0%
#118305000000
1!
1%
#118310000000
0!
0%
#118315000000
1!
1%
#118320000000
0!
0%
#118325000000
1!
1%
#118330000000
0!
0%
#118335000000
1!
1%
#118340000000
0!
0%
#118345000000
1!
1%
#118350000000
0!
0%
#118355000000
1!
1%
#118360000000
0!
0%
#118365000000
1!
1%
#118370000000
0!
0%
#118375000000
1!
1%
#118380000000
0!
0%
#118385000000
1!
1%
#118390000000
0!
0%
#118395000000
1!
1%
#118400000000
0!
0%
#118405000000
1!
1%
#118410000000
0!
0%
#118415000000
1!
1%
#118420000000
0!
0%
#118425000000
1!
1%
#118430000000
0!
0%
#118435000000
1!
1%
#118440000000
0!
0%
#118445000000
1!
1%
#118450000000
0!
0%
#118455000000
1!
1%
#118460000000
0!
0%
#118465000000
1!
1%
#118470000000
0!
0%
#118475000000
1!
1%
#118480000000
0!
0%
#118485000000
1!
1%
#118490000000
0!
0%
#118495000000
1!
1%
#118500000000
0!
0%
#118505000000
1!
1%
#118510000000
0!
0%
#118515000000
1!
1%
#118520000000
0!
0%
#118525000000
1!
1%
#118530000000
0!
0%
#118535000000
1!
1%
#118540000000
0!
0%
#118545000000
1!
1%
#118550000000
0!
0%
#118555000000
1!
1%
#118560000000
0!
0%
#118565000000
1!
1%
#118570000000
0!
0%
#118575000000
1!
1%
#118580000000
0!
0%
#118585000000
1!
1%
#118590000000
0!
0%
#118595000000
1!
1%
#118600000000
0!
0%
#118605000000
1!
1%
#118610000000
0!
0%
#118615000000
1!
1%
#118620000000
0!
0%
#118625000000
1!
1%
#118630000000
0!
0%
#118635000000
1!
1%
#118640000000
0!
0%
#118645000000
1!
1%
#118650000000
0!
0%
#118655000000
1!
1%
#118660000000
0!
0%
#118665000000
1!
1%
#118670000000
0!
0%
#118675000000
1!
1%
#118680000000
0!
0%
#118685000000
1!
1%
#118690000000
0!
0%
#118695000000
1!
1%
#118700000000
0!
0%
#118705000000
1!
1%
#118710000000
0!
0%
#118715000000
1!
1%
#118720000000
0!
0%
#118725000000
1!
1%
#118730000000
0!
0%
#118735000000
1!
1%
#118740000000
0!
0%
#118745000000
1!
1%
#118750000000
0!
0%
#118755000000
1!
1%
#118760000000
0!
0%
#118765000000
1!
1%
#118770000000
0!
0%
#118775000000
1!
1%
#118780000000
0!
0%
#118785000000
1!
1%
#118790000000
0!
0%
#118795000000
1!
1%
#118800000000
0!
0%
#118805000000
1!
1%
#118810000000
0!
0%
#118815000000
1!
1%
#118820000000
0!
0%
#118825000000
1!
1%
#118830000000
0!
0%
#118835000000
1!
1%
#118840000000
0!
0%
#118845000000
1!
1%
#118850000000
0!
0%
#118855000000
1!
1%
#118860000000
0!
0%
#118865000000
1!
1%
#118870000000
0!
0%
#118875000000
1!
1%
#118880000000
0!
0%
#118885000000
1!
1%
#118890000000
0!
0%
#118895000000
1!
1%
#118900000000
0!
0%
#118905000000
1!
1%
#118910000000
0!
0%
#118915000000
1!
1%
#118920000000
0!
0%
#118925000000
1!
1%
#118930000000
0!
0%
#118935000000
1!
1%
#118940000000
0!
0%
#118945000000
1!
1%
#118950000000
0!
0%
#118955000000
1!
1%
#118960000000
0!
0%
#118965000000
1!
1%
#118970000000
0!
0%
#118975000000
1!
1%
#118980000000
0!
0%
#118985000000
1!
1%
#118990000000
0!
0%
#118995000000
1!
1%
#119000000000
0!
0%
#119005000000
1!
1%
#119010000000
0!
0%
#119015000000
1!
1%
#119020000000
0!
0%
#119025000000
1!
1%
#119030000000
0!
0%
#119035000000
1!
1%
#119040000000
0!
0%
#119045000000
1!
1%
#119050000000
0!
0%
#119055000000
1!
1%
#119060000000
0!
0%
#119065000000
1!
1%
#119070000000
0!
0%
#119075000000
1!
1%
#119080000000
0!
0%
#119085000000
1!
1%
#119090000000
0!
0%
#119095000000
1!
1%
#119100000000
0!
0%
#119105000000
1!
1%
#119110000000
0!
0%
#119115000000
1!
1%
#119120000000
0!
0%
#119125000000
1!
1%
#119130000000
0!
0%
#119135000000
1!
1%
#119140000000
0!
0%
#119145000000
1!
1%
#119150000000
0!
0%
#119155000000
1!
1%
#119160000000
0!
0%
#119165000000
1!
1%
#119170000000
0!
0%
#119175000000
1!
1%
#119180000000
0!
0%
#119185000000
1!
1%
#119190000000
0!
0%
#119195000000
1!
1%
#119200000000
0!
0%
#119205000000
1!
1%
#119210000000
0!
0%
#119215000000
1!
1%
#119220000000
0!
0%
#119225000000
1!
1%
#119230000000
0!
0%
#119235000000
1!
1%
#119240000000
0!
0%
#119245000000
1!
1%
#119250000000
0!
0%
#119255000000
1!
1%
#119260000000
0!
0%
#119265000000
1!
1%
#119270000000
0!
0%
#119275000000
1!
1%
#119280000000
0!
0%
#119285000000
1!
1%
#119290000000
0!
0%
#119295000000
1!
1%
#119300000000
0!
0%
#119305000000
1!
1%
#119310000000
0!
0%
#119315000000
1!
1%
#119320000000
0!
0%
#119325000000
1!
1%
#119330000000
0!
0%
#119335000000
1!
1%
#119340000000
0!
0%
#119345000000
1!
1%
#119350000000
0!
0%
#119355000000
1!
1%
#119360000000
0!
0%
#119365000000
1!
1%
#119370000000
0!
0%
#119375000000
1!
1%
#119380000000
0!
0%
#119385000000
1!
1%
#119390000000
0!
0%
#119395000000
1!
1%
#119400000000
0!
0%
#119405000000
1!
1%
#119410000000
0!
0%
#119415000000
1!
1%
#119420000000
0!
0%
#119425000000
1!
1%
#119430000000
0!
0%
#119435000000
1!
1%
#119440000000
0!
0%
#119445000000
1!
1%
#119450000000
0!
0%
#119455000000
1!
1%
#119460000000
0!
0%
#119465000000
1!
1%
#119470000000
0!
0%
#119475000000
1!
1%
#119480000000
0!
0%
#119485000000
1!
1%
#119490000000
0!
0%
#119495000000
1!
1%
#119500000000
0!
0%
#119505000000
1!
1%
#119510000000
0!
0%
#119515000000
1!
1%
#119520000000
0!
0%
#119525000000
1!
1%
#119530000000
0!
0%
#119535000000
1!
1%
#119540000000
0!
0%
#119545000000
1!
1%
#119550000000
0!
0%
#119555000000
1!
1%
#119560000000
0!
0%
#119565000000
1!
1%
#119570000000
0!
0%
#119575000000
1!
1%
#119580000000
0!
0%
#119585000000
1!
1%
#119590000000
0!
0%
#119595000000
1!
1%
#119600000000
0!
0%
#119605000000
1!
1%
#119610000000
0!
0%
#119615000000
1!
1%
#119620000000
0!
0%
#119625000000
1!
1%
#119630000000
0!
0%
#119635000000
1!
1%
#119640000000
0!
0%
#119645000000
1!
1%
#119650000000
0!
0%
#119655000000
1!
1%
#119660000000
0!
0%
#119665000000
1!
1%
#119670000000
0!
0%
#119675000000
1!
1%
#119680000000
0!
0%
#119685000000
1!
1%
#119690000000
0!
0%
#119695000000
1!
1%
#119700000000
0!
0%
#119705000000
1!
1%
#119710000000
0!
0%
#119715000000
1!
1%
#119720000000
0!
0%
#119725000000
1!
1%
#119730000000
0!
0%
#119735000000
1!
1%
#119740000000
0!
0%
#119745000000
1!
1%
#119750000000
0!
0%
#119755000000
1!
1%
#119760000000
0!
0%
#119765000000
1!
1%
#119770000000
0!
0%
#119775000000
1!
1%
#119780000000
0!
0%
#119785000000
1!
1%
#119790000000
0!
0%
#119795000000
1!
1%
#119800000000
0!
0%
#119805000000
1!
1%
#119810000000
0!
0%
#119815000000
1!
1%
#119820000000
0!
0%
#119825000000
1!
1%
#119830000000
0!
0%
#119835000000
1!
1%
#119840000000
0!
0%
#119845000000
1!
1%
#119850000000
0!
0%
#119855000000
1!
1%
#119860000000
0!
0%
#119865000000
1!
1%
#119870000000
0!
0%
#119875000000
1!
1%
#119880000000
0!
0%
#119885000000
1!
1%
#119890000000
0!
0%
#119895000000
1!
1%
#119900000000
0!
0%
#119905000000
1!
1%
#119910000000
0!
0%
#119915000000
1!
1%
#119920000000
0!
0%
#119925000000
1!
1%
#119930000000
0!
0%
#119935000000
1!
1%
#119940000000
0!
0%
#119945000000
1!
1%
#119950000000
0!
0%
#119955000000
1!
1%
#119960000000
0!
0%
#119965000000
1!
1%
#119970000000
0!
0%
#119975000000
1!
1%
#119980000000
0!
0%
#119985000000
1!
1%
#119990000000
0!
0%
#119995000000
1!
1%
#120000000000
0!
0%
#120005000000
1!
1%
#120010000000
0!
0%
#120015000000
1!
1%
#120020000000
0!
0%
#120025000000
1!
1%
#120030000000
0!
0%
#120035000000
1!
1%
#120040000000
0!
0%
#120045000000
1!
1%
#120050000000
0!
0%
#120055000000
1!
1%
#120060000000
0!
0%
#120065000000
1!
1%
#120070000000
0!
0%
#120075000000
1!
1%
#120080000000
0!
0%
#120085000000
1!
1%
#120090000000
0!
0%
#120095000000
1!
1%
#120100000000
0!
0%
#120105000000
1!
1%
#120110000000
0!
0%
#120115000000
1!
1%
#120120000000
0!
0%
#120125000000
1!
1%
#120130000000
0!
0%
#120135000000
1!
1%
#120140000000
0!
0%
#120145000000
1!
1%
#120150000000
0!
0%
#120155000000
1!
1%
#120160000000
0!
0%
#120165000000
1!
1%
#120170000000
0!
0%
#120175000000
1!
1%
#120180000000
0!
0%
#120185000000
1!
1%
#120190000000
0!
0%
#120195000000
1!
1%
#120200000000
0!
0%
#120205000000
1!
1%
#120210000000
0!
0%
#120215000000
1!
1%
#120220000000
0!
0%
#120225000000
1!
1%
#120230000000
0!
0%
#120235000000
1!
1%
#120240000000
0!
0%
#120245000000
1!
1%
#120250000000
0!
0%
#120255000000
1!
1%
#120260000000
0!
0%
#120265000000
1!
1%
#120270000000
0!
0%
#120275000000
1!
1%
#120280000000
0!
0%
#120285000000
1!
1%
#120290000000
0!
0%
#120295000000
1!
1%
#120300000000
0!
0%
#120305000000
1!
1%
#120310000000
0!
0%
#120315000000
1!
1%
#120320000000
0!
0%
#120325000000
1!
1%
#120330000000
0!
0%
#120335000000
1!
1%
#120340000000
0!
0%
#120345000000
1!
1%
#120350000000
0!
0%
#120355000000
1!
1%
#120360000000
0!
0%
#120365000000
1!
1%
#120370000000
0!
0%
#120375000000
1!
1%
#120380000000
0!
0%
#120385000000
1!
1%
#120390000000
0!
0%
#120395000000
1!
1%
#120400000000
0!
0%
#120405000000
1!
1%
#120410000000
0!
0%
#120415000000
1!
1%
#120420000000
0!
0%
#120425000000
1!
1%
#120430000000
0!
0%
#120435000000
1!
1%
#120440000000
0!
0%
#120445000000
1!
1%
#120450000000
0!
0%
#120455000000
1!
1%
#120460000000
0!
0%
#120465000000
1!
1%
#120470000000
0!
0%
#120475000000
1!
1%
#120480000000
0!
0%
#120485000000
1!
1%
#120490000000
0!
0%
#120495000000
1!
1%
#120500000000
0!
0%
#120505000000
1!
1%
#120510000000
0!
0%
#120515000000
1!
1%
#120520000000
0!
0%
#120525000000
1!
1%
#120530000000
0!
0%
#120535000000
1!
1%
#120540000000
0!
0%
#120545000000
1!
1%
#120550000000
0!
0%
#120555000000
1!
1%
#120560000000
0!
0%
#120565000000
1!
1%
#120570000000
0!
0%
#120575000000
1!
1%
#120580000000
0!
0%
#120585000000
1!
1%
#120590000000
0!
0%
#120595000000
1!
1%
#120600000000
0!
0%
#120605000000
1!
1%
#120610000000
0!
0%
#120615000000
1!
1%
#120620000000
0!
0%
#120625000000
1!
1%
#120630000000
0!
0%
#120635000000
1!
1%
#120640000000
0!
0%
#120645000000
1!
1%
#120650000000
0!
0%
#120655000000
1!
1%
#120660000000
0!
0%
#120665000000
1!
1%
#120670000000
0!
0%
#120675000000
1!
1%
#120680000000
0!
0%
#120685000000
1!
1%
#120690000000
0!
0%
#120695000000
1!
1%
#120700000000
0!
0%
#120705000000
1!
1%
#120710000000
0!
0%
#120715000000
1!
1%
#120720000000
0!
0%
#120725000000
1!
1%
#120730000000
0!
0%
#120735000000
1!
1%
#120740000000
0!
0%
#120745000000
1!
1%
#120750000000
0!
0%
#120755000000
1!
1%
#120760000000
0!
0%
#120765000000
1!
1%
#120770000000
0!
0%
#120775000000
1!
1%
#120780000000
0!
0%
#120785000000
1!
1%
#120790000000
0!
0%
#120795000000
1!
1%
#120800000000
0!
0%
#120805000000
1!
1%
#120810000000
0!
0%
#120815000000
1!
1%
#120820000000
0!
0%
#120825000000
1!
1%
#120830000000
0!
0%
#120835000000
1!
1%
#120840000000
0!
0%
#120845000000
1!
1%
#120850000000
0!
0%
#120855000000
1!
1%
#120860000000
0!
0%
#120865000000
1!
1%
#120870000000
0!
0%
#120875000000
1!
1%
#120880000000
0!
0%
#120885000000
1!
1%
#120890000000
0!
0%
#120895000000
1!
1%
#120900000000
0!
0%
#120905000000
1!
1%
#120910000000
0!
0%
#120915000000
1!
1%
#120920000000
0!
0%
#120925000000
1!
1%
#120930000000
0!
0%
#120935000000
1!
1%
#120940000000
0!
0%
#120945000000
1!
1%
#120950000000
0!
0%
#120955000000
1!
1%
#120960000000
0!
0%
#120965000000
1!
1%
#120970000000
0!
0%
#120975000000
1!
1%
#120980000000
0!
0%
#120985000000
1!
1%
#120990000000
0!
0%
#120995000000
1!
1%
#121000000000
0!
0%
#121005000000
1!
1%
#121010000000
0!
0%
#121015000000
1!
1%
#121020000000
0!
0%
#121025000000
1!
1%
#121030000000
0!
0%
#121035000000
1!
1%
#121040000000
0!
0%
#121045000000
1!
1%
#121050000000
0!
0%
#121055000000
1!
1%
#121060000000
0!
0%
#121065000000
1!
1%
#121070000000
0!
0%
#121075000000
1!
1%
#121080000000
0!
0%
#121085000000
1!
1%
#121090000000
0!
0%
#121095000000
1!
1%
#121100000000
0!
0%
#121105000000
1!
1%
#121110000000
0!
0%
#121115000000
1!
1%
#121120000000
0!
0%
#121125000000
1!
1%
#121130000000
0!
0%
#121135000000
1!
1%
#121140000000
0!
0%
#121145000000
1!
1%
#121150000000
0!
0%
#121155000000
1!
1%
#121160000000
0!
0%
#121165000000
1!
1%
#121170000000
0!
0%
#121175000000
1!
1%
#121180000000
0!
0%
#121185000000
1!
1%
#121190000000
0!
0%
#121195000000
1!
1%
#121200000000
0!
0%
#121205000000
1!
1%
#121210000000
0!
0%
#121215000000
1!
1%
#121220000000
0!
0%
#121225000000
1!
1%
#121230000000
0!
0%
#121235000000
1!
1%
#121240000000
0!
0%
#121245000000
1!
1%
#121250000000
0!
0%
#121255000000
1!
1%
#121260000000
0!
0%
#121265000000
1!
1%
#121270000000
0!
0%
#121275000000
1!
1%
#121280000000
0!
0%
#121285000000
1!
1%
#121290000000
0!
0%
#121295000000
1!
1%
#121300000000
0!
0%
#121305000000
1!
1%
#121310000000
0!
0%
#121315000000
1!
1%
#121320000000
0!
0%
#121325000000
1!
1%
#121330000000
0!
0%
#121335000000
1!
1%
#121340000000
0!
0%
#121345000000
1!
1%
#121350000000
0!
0%
#121355000000
1!
1%
#121360000000
0!
0%
#121365000000
1!
1%
#121370000000
0!
0%
#121375000000
1!
1%
#121380000000
0!
0%
#121385000000
1!
1%
#121390000000
0!
0%
#121395000000
1!
1%
#121400000000
0!
0%
#121405000000
1!
1%
#121410000000
0!
0%
#121415000000
1!
1%
#121420000000
0!
0%
#121425000000
1!
1%
#121430000000
0!
0%
#121435000000
1!
1%
#121440000000
0!
0%
#121445000000
1!
1%
#121450000000
0!
0%
#121455000000
1!
1%
#121460000000
0!
0%
#121465000000
1!
1%
#121470000000
0!
0%
#121475000000
1!
1%
#121480000000
0!
0%
#121485000000
1!
1%
#121490000000
0!
0%
#121495000000
1!
1%
#121500000000
0!
0%
#121505000000
1!
1%
#121510000000
0!
0%
#121515000000
1!
1%
#121520000000
0!
0%
#121525000000
1!
1%
#121530000000
0!
0%
#121535000000
1!
1%
#121540000000
0!
0%
#121545000000
1!
1%
#121550000000
0!
0%
#121555000000
1!
1%
#121560000000
0!
0%
#121565000000
1!
1%
#121570000000
0!
0%
#121575000000
1!
1%
#121580000000
0!
0%
#121585000000
1!
1%
#121590000000
0!
0%
#121595000000
1!
1%
#121600000000
0!
0%
#121605000000
1!
1%
#121610000000
0!
0%
#121615000000
1!
1%
#121620000000
0!
0%
#121625000000
1!
1%
#121630000000
0!
0%
#121635000000
1!
1%
#121640000000
0!
0%
#121645000000
1!
1%
#121650000000
0!
0%
#121655000000
1!
1%
#121660000000
0!
0%
#121665000000
1!
1%
#121670000000
0!
0%
#121675000000
1!
1%
#121680000000
0!
0%
#121685000000
1!
1%
#121690000000
0!
0%
#121695000000
1!
1%
#121700000000
0!
0%
#121705000000
1!
1%
#121710000000
0!
0%
#121715000000
1!
1%
#121720000000
0!
0%
#121725000000
1!
1%
#121730000000
0!
0%
#121735000000
1!
1%
#121740000000
0!
0%
#121745000000
1!
1%
#121750000000
0!
0%
#121755000000
1!
1%
#121760000000
0!
0%
#121765000000
1!
1%
#121770000000
0!
0%
#121775000000
1!
1%
#121780000000
0!
0%
#121785000000
1!
1%
#121790000000
0!
0%
#121795000000
1!
1%
#121800000000
0!
0%
#121805000000
1!
1%
#121810000000
0!
0%
#121815000000
1!
1%
#121820000000
0!
0%
#121825000000
1!
1%
#121830000000
0!
0%
#121835000000
1!
1%
#121840000000
0!
0%
#121845000000
1!
1%
#121850000000
0!
0%
#121855000000
1!
1%
#121860000000
0!
0%
#121865000000
1!
1%
#121870000000
0!
0%
#121875000000
1!
1%
#121880000000
0!
0%
#121885000000
1!
1%
#121890000000
0!
0%
#121895000000
1!
1%
#121900000000
0!
0%
#121905000000
1!
1%
#121910000000
0!
0%
#121915000000
1!
1%
#121920000000
0!
0%
#121925000000
1!
1%
#121930000000
0!
0%
#121935000000
1!
1%
#121940000000
0!
0%
#121945000000
1!
1%
#121950000000
0!
0%
#121955000000
1!
1%
#121960000000
0!
0%
#121965000000
1!
1%
#121970000000
0!
0%
#121975000000
1!
1%
#121980000000
0!
0%
#121985000000
1!
1%
#121990000000
0!
0%
#121995000000
1!
1%
#122000000000
0!
0%
#122005000000
1!
1%
#122010000000
0!
0%
#122015000000
1!
1%
#122020000000
0!
0%
#122025000000
1!
1%
#122030000000
0!
0%
#122035000000
1!
1%
#122040000000
0!
0%
#122045000000
1!
1%
#122050000000
0!
0%
#122055000000
1!
1%
#122060000000
0!
0%
#122065000000
1!
1%
#122070000000
0!
0%
#122075000000
1!
1%
#122080000000
0!
0%
#122085000000
1!
1%
#122090000000
0!
0%
#122095000000
1!
1%
#122100000000
0!
0%
#122105000000
1!
1%
#122110000000
0!
0%
#122115000000
1!
1%
#122120000000
0!
0%
#122125000000
1!
1%
#122130000000
0!
0%
#122135000000
1!
1%
#122140000000
0!
0%
#122145000000
1!
1%
#122150000000
0!
0%
#122155000000
1!
1%
#122160000000
0!
0%
#122165000000
1!
1%
#122170000000
0!
0%
#122175000000
1!
1%
#122180000000
0!
0%
#122185000000
1!
1%
#122190000000
0!
0%
#122195000000
1!
1%
#122200000000
0!
0%
#122205000000
1!
1%
#122210000000
0!
0%
#122215000000
1!
1%
#122220000000
0!
0%
#122225000000
1!
1%
#122230000000
0!
0%
#122235000000
1!
1%
#122240000000
0!
0%
#122245000000
1!
1%
#122250000000
0!
0%
#122255000000
1!
1%
#122260000000
0!
0%
#122265000000
1!
1%
#122270000000
0!
0%
#122275000000
1!
1%
#122280000000
0!
0%
#122285000000
1!
1%
#122290000000
0!
0%
#122295000000
1!
1%
#122300000000
0!
0%
#122305000000
1!
1%
#122310000000
0!
0%
#122315000000
1!
1%
#122320000000
0!
0%
#122325000000
1!
1%
#122330000000
0!
0%
#122335000000
1!
1%
#122340000000
0!
0%
#122345000000
1!
1%
#122350000000
0!
0%
#122355000000
1!
1%
#122360000000
0!
0%
#122365000000
1!
1%
#122370000000
0!
0%
#122375000000
1!
1%
#122380000000
0!
0%
#122385000000
1!
1%
#122390000000
0!
0%
#122395000000
1!
1%
#122400000000
0!
0%
#122405000000
1!
1%
#122410000000
0!
0%
#122415000000
1!
1%
#122420000000
0!
0%
#122425000000
1!
1%
#122430000000
0!
0%
#122435000000
1!
1%
#122440000000
0!
0%
#122445000000
1!
1%
#122450000000
0!
0%
#122455000000
1!
1%
#122460000000
0!
0%
#122465000000
1!
1%
#122470000000
0!
0%
#122475000000
1!
1%
#122480000000
0!
0%
#122485000000
1!
1%
#122490000000
0!
0%
#122495000000
1!
1%
#122500000000
0!
0%
#122505000000
1!
1%
#122510000000
0!
0%
#122515000000
1!
1%
#122520000000
0!
0%
#122525000000
1!
1%
#122530000000
0!
0%
#122535000000
1!
1%
#122540000000
0!
0%
#122545000000
1!
1%
#122550000000
0!
0%
#122555000000
1!
1%
#122560000000
0!
0%
#122565000000
1!
1%
#122570000000
0!
0%
#122575000000
1!
1%
#122580000000
0!
0%
#122585000000
1!
1%
#122590000000
0!
0%
#122595000000
1!
1%
#122600000000
0!
0%
#122605000000
1!
1%
#122610000000
0!
0%
#122615000000
1!
1%
#122620000000
0!
0%
#122625000000
1!
1%
#122630000000
0!
0%
#122635000000
1!
1%
#122640000000
0!
0%
#122645000000
1!
1%
#122650000000
0!
0%
#122655000000
1!
1%
#122660000000
0!
0%
#122665000000
1!
1%
#122670000000
0!
0%
#122675000000
1!
1%
#122680000000
0!
0%
#122685000000
1!
1%
#122690000000
0!
0%
#122695000000
1!
1%
#122700000000
0!
0%
#122705000000
1!
1%
#122710000000
0!
0%
#122715000000
1!
1%
#122720000000
0!
0%
#122725000000
1!
1%
#122730000000
0!
0%
#122735000000
1!
1%
#122740000000
0!
0%
#122745000000
1!
1%
#122750000000
0!
0%
#122755000000
1!
1%
#122760000000
0!
0%
#122765000000
1!
1%
#122770000000
0!
0%
#122775000000
1!
1%
#122780000000
0!
0%
#122785000000
1!
1%
#122790000000
0!
0%
#122795000000
1!
1%
#122800000000
0!
0%
#122805000000
1!
1%
#122810000000
0!
0%
#122815000000
1!
1%
#122820000000
0!
0%
#122825000000
1!
1%
#122830000000
0!
0%
#122835000000
1!
1%
#122840000000
0!
0%
#122845000000
1!
1%
#122850000000
0!
0%
#122855000000
1!
1%
#122860000000
0!
0%
#122865000000
1!
1%
#122870000000
0!
0%
#122875000000
1!
1%
#122880000000
0!
0%
#122885000000
1!
1%
#122890000000
0!
0%
#122895000000
1!
1%
#122900000000
0!
0%
#122905000000
1!
1%
#122910000000
0!
0%
#122915000000
1!
1%
#122920000000
0!
0%
#122925000000
1!
1%
#122930000000
0!
0%
#122935000000
1!
1%
#122940000000
0!
0%
#122945000000
1!
1%
#122950000000
0!
0%
#122955000000
1!
1%
#122960000000
0!
0%
#122965000000
1!
1%
#122970000000
0!
0%
#122975000000
1!
1%
#122980000000
0!
0%
#122985000000
1!
1%
#122990000000
0!
0%
#122995000000
1!
1%
#123000000000
0!
0%
#123005000000
1!
1%
#123010000000
0!
0%
#123015000000
1!
1%
#123020000000
0!
0%
#123025000000
1!
1%
#123030000000
0!
0%
#123035000000
1!
1%
#123040000000
0!
0%
#123045000000
1!
1%
#123050000000
0!
0%
#123055000000
1!
1%
#123060000000
0!
0%
#123065000000
1!
1%
#123070000000
0!
0%
#123075000000
1!
1%
#123080000000
0!
0%
#123085000000
1!
1%
#123090000000
0!
0%
#123095000000
1!
1%
#123100000000
0!
0%
#123105000000
1!
1%
#123110000000
0!
0%
#123115000000
1!
1%
#123120000000
0!
0%
#123125000000
1!
1%
#123130000000
0!
0%
#123135000000
1!
1%
#123140000000
0!
0%
#123145000000
1!
1%
#123150000000
0!
0%
#123155000000
1!
1%
#123160000000
0!
0%
#123165000000
1!
1%
#123170000000
0!
0%
#123175000000
1!
1%
#123180000000
0!
0%
#123185000000
1!
1%
#123190000000
0!
0%
#123195000000
1!
1%
#123200000000
0!
0%
#123205000000
1!
1%
#123210000000
0!
0%
#123215000000
1!
1%
#123220000000
0!
0%
#123225000000
1!
1%
#123230000000
0!
0%
#123235000000
1!
1%
#123240000000
0!
0%
#123245000000
1!
1%
#123250000000
0!
0%
#123255000000
1!
1%
#123260000000
0!
0%
#123265000000
1!
1%
#123270000000
0!
0%
#123275000000
1!
1%
#123280000000
0!
0%
#123285000000
1!
1%
#123290000000
0!
0%
#123295000000
1!
1%
#123300000000
0!
0%
#123305000000
1!
1%
#123310000000
0!
0%
#123315000000
1!
1%
#123320000000
0!
0%
#123325000000
1!
1%
#123330000000
0!
0%
#123335000000
1!
1%
#123340000000
0!
0%
#123345000000
1!
1%
#123350000000
0!
0%
#123355000000
1!
1%
#123360000000
0!
0%
#123365000000
1!
1%
#123370000000
0!
0%
#123375000000
1!
1%
#123380000000
0!
0%
#123385000000
1!
1%
#123390000000
0!
0%
#123395000000
1!
1%
#123400000000
0!
0%
#123405000000
1!
1%
#123410000000
0!
0%
#123415000000
1!
1%
#123420000000
0!
0%
#123425000000
1!
1%
#123430000000
0!
0%
#123435000000
1!
1%
#123440000000
0!
0%
#123445000000
1!
1%
#123450000000
0!
0%
#123455000000
1!
1%
#123460000000
0!
0%
#123465000000
1!
1%
#123470000000
0!
0%
#123475000000
1!
1%
#123480000000
0!
0%
#123485000000
1!
1%
#123490000000
0!
0%
#123495000000
1!
1%
#123500000000
0!
0%
#123505000000
1!
1%
#123510000000
0!
0%
#123515000000
1!
1%
#123520000000
0!
0%
#123525000000
1!
1%
#123530000000
0!
0%
#123535000000
1!
1%
#123540000000
0!
0%
#123545000000
1!
1%
#123550000000
0!
0%
#123555000000
1!
1%
#123560000000
0!
0%
#123565000000
1!
1%
#123570000000
0!
0%
#123575000000
1!
1%
#123580000000
0!
0%
#123585000000
1!
1%
#123590000000
0!
0%
#123595000000
1!
1%
#123600000000
0!
0%
#123605000000
1!
1%
#123610000000
0!
0%
#123615000000
1!
1%
#123620000000
0!
0%
#123625000000
1!
1%
#123630000000
0!
0%
#123635000000
1!
1%
#123640000000
0!
0%
#123645000000
1!
1%
#123650000000
0!
0%
#123655000000
1!
1%
#123660000000
0!
0%
#123665000000
1!
1%
#123670000000
0!
0%
#123675000000
1!
1%
#123680000000
0!
0%
#123685000000
1!
1%
#123690000000
0!
0%
#123695000000
1!
1%
#123700000000
0!
0%
#123705000000
1!
1%
#123710000000
0!
0%
#123715000000
1!
1%
#123720000000
0!
0%
#123725000000
1!
1%
#123730000000
0!
0%
#123735000000
1!
1%
#123740000000
0!
0%
#123745000000
1!
1%
#123750000000
0!
0%
#123755000000
1!
1%
#123760000000
0!
0%
#123765000000
1!
1%
#123770000000
0!
0%
#123775000000
1!
1%
#123780000000
0!
0%
#123785000000
1!
1%
#123790000000
0!
0%
#123795000000
1!
1%
#123800000000
0!
0%
#123805000000
1!
1%
#123810000000
0!
0%
#123815000000
1!
1%
#123820000000
0!
0%
#123825000000
1!
1%
#123830000000
0!
0%
#123835000000
1!
1%
#123840000000
0!
0%
#123845000000
1!
1%
#123850000000
0!
0%
#123855000000
1!
1%
#123860000000
0!
0%
#123865000000
1!
1%
#123870000000
0!
0%
#123875000000
1!
1%
#123880000000
0!
0%
#123885000000
1!
1%
#123890000000
0!
0%
#123895000000
1!
1%
#123900000000
0!
0%
#123905000000
1!
1%
#123910000000
0!
0%
#123915000000
1!
1%
#123920000000
0!
0%
#123925000000
1!
1%
#123930000000
0!
0%
#123935000000
1!
1%
#123940000000
0!
0%
#123945000000
1!
1%
#123950000000
0!
0%
#123955000000
1!
1%
#123960000000
0!
0%
#123965000000
1!
1%
#123970000000
0!
0%
#123975000000
1!
1%
#123980000000
0!
0%
#123985000000
1!
1%
#123990000000
0!
0%
#123995000000
1!
1%
#124000000000
0!
0%
#124005000000
1!
1%
#124010000000
0!
0%
#124015000000
1!
1%
#124020000000
0!
0%
#124025000000
1!
1%
#124030000000
0!
0%
#124035000000
1!
1%
#124040000000
0!
0%
#124045000000
1!
1%
#124050000000
0!
0%
#124055000000
1!
1%
#124060000000
0!
0%
#124065000000
1!
1%
#124070000000
0!
0%
#124075000000
1!
1%
#124080000000
0!
0%
#124085000000
1!
1%
#124090000000
0!
0%
#124095000000
1!
1%
#124100000000
0!
0%
#124105000000
1!
1%
#124110000000
0!
0%
#124115000000
1!
1%
#124120000000
0!
0%
#124125000000
1!
1%
#124130000000
0!
0%
#124135000000
1!
1%
#124140000000
0!
0%
#124145000000
1!
1%
#124150000000
0!
0%
#124155000000
1!
1%
#124160000000
0!
0%
#124165000000
1!
1%
#124170000000
0!
0%
#124175000000
1!
1%
#124180000000
0!
0%
#124185000000
1!
1%
#124190000000
0!
0%
#124195000000
1!
1%
#124200000000
0!
0%
#124205000000
1!
1%
#124210000000
0!
0%
#124215000000
1!
1%
#124220000000
0!
0%
#124225000000
1!
1%
#124230000000
0!
0%
#124235000000
1!
1%
#124240000000
0!
0%
#124245000000
1!
1%
#124250000000
0!
0%
#124255000000
1!
1%
#124260000000
0!
0%
#124265000000
1!
1%
#124270000000
0!
0%
#124275000000
1!
1%
#124280000000
0!
0%
#124285000000
1!
1%
#124290000000
0!
0%
#124295000000
1!
1%
#124300000000
0!
0%
#124305000000
1!
1%
#124310000000
0!
0%
#124315000000
1!
1%
#124320000000
0!
0%
#124325000000
1!
1%
#124330000000
0!
0%
#124335000000
1!
1%
#124340000000
0!
0%
#124345000000
1!
1%
#124350000000
0!
0%
#124355000000
1!
1%
#124360000000
0!
0%
#124365000000
1!
1%
#124370000000
0!
0%
#124375000000
1!
1%
#124380000000
0!
0%
#124385000000
1!
1%
#124390000000
0!
0%
#124395000000
1!
1%
#124400000000
0!
0%
#124405000000
1!
1%
#124410000000
0!
0%
#124415000000
1!
1%
#124420000000
0!
0%
#124425000000
1!
1%
#124430000000
0!
0%
#124435000000
1!
1%
#124440000000
0!
0%
#124445000000
1!
1%
#124450000000
0!
0%
#124455000000
1!
1%
#124460000000
0!
0%
#124465000000
1!
1%
#124470000000
0!
0%
#124475000000
1!
1%
#124480000000
0!
0%
#124485000000
1!
1%
#124490000000
0!
0%
#124495000000
1!
1%
#124500000000
0!
0%
#124505000000
1!
1%
#124510000000
0!
0%
#124515000000
1!
1%
#124520000000
0!
0%
#124525000000
1!
1%
#124530000000
0!
0%
#124535000000
1!
1%
#124540000000
0!
0%
#124545000000
1!
1%
#124550000000
0!
0%
#124555000000
1!
1%
#124560000000
0!
0%
#124565000000
1!
1%
#124570000000
0!
0%
#124575000000
1!
1%
#124580000000
0!
0%
#124585000000
1!
1%
#124590000000
0!
0%
#124595000000
1!
1%
#124600000000
0!
0%
#124605000000
1!
1%
#124610000000
0!
0%
#124615000000
1!
1%
#124620000000
0!
0%
#124625000000
1!
1%
#124630000000
0!
0%
#124635000000
1!
1%
#124640000000
0!
0%
#124645000000
1!
1%
#124650000000
0!
0%
#124655000000
1!
1%
#124660000000
0!
0%
#124665000000
1!
1%
#124670000000
0!
0%
#124675000000
1!
1%
#124680000000
0!
0%
#124685000000
1!
1%
#124690000000
0!
0%
#124695000000
1!
1%
#124700000000
0!
0%
#124705000000
1!
1%
#124710000000
0!
0%
#124715000000
1!
1%
#124720000000
0!
0%
#124725000000
1!
1%
#124730000000
0!
0%
#124735000000
1!
1%
#124740000000
0!
0%
#124745000000
1!
1%
#124750000000
0!
0%
#124755000000
1!
1%
#124760000000
0!
0%
#124765000000
1!
1%
#124770000000
0!
0%
#124775000000
1!
1%
#124780000000
0!
0%
#124785000000
1!
1%
#124790000000
0!
0%
#124795000000
1!
1%
#124800000000
0!
0%
#124805000000
1!
1%
#124810000000
0!
0%
#124815000000
1!
1%
#124820000000
0!
0%
#124825000000
1!
1%
#124830000000
0!
0%
#124835000000
1!
1%
#124840000000
0!
0%
#124845000000
1!
1%
#124850000000
0!
0%
#124855000000
1!
1%
#124860000000
0!
0%
#124865000000
1!
1%
#124870000000
0!
0%
#124875000000
1!
1%
#124880000000
0!
0%
#124885000000
1!
1%
#124890000000
0!
0%
#124895000000
1!
1%
#124900000000
0!
0%
#124905000000
1!
1%
#124910000000
0!
0%
#124915000000
1!
1%
#124920000000
0!
0%
#124925000000
1!
1%
#124930000000
0!
0%
#124935000000
1!
1%
#124940000000
0!
0%
#124945000000
1!
1%
#124950000000
0!
0%
#124955000000
1!
1%
#124960000000
0!
0%
#124965000000
1!
1%
#124970000000
0!
0%
#124975000000
1!
1%
#124980000000
0!
0%
#124985000000
1!
1%
#124990000000
0!
0%
#124995000000
1!
1%
#125000000000
0!
0%
#125005000000
1!
1%
#125010000000
0!
0%
#125015000000
1!
1%
#125020000000
0!
0%
#125025000000
1!
1%
#125030000000
0!
0%
#125035000000
1!
1%
#125040000000
0!
0%
#125045000000
1!
1%
#125050000000
0!
0%
#125055000000
1!
1%
#125060000000
0!
0%
#125065000000
1!
1%
#125070000000
0!
0%
#125075000000
1!
1%
#125080000000
0!
0%
#125085000000
1!
1%
#125090000000
0!
0%
#125095000000
1!
1%
#125100000000
0!
0%
#125105000000
1!
1%
#125110000000
0!
0%
#125115000000
1!
1%
#125120000000
0!
0%
#125125000000
1!
1%
#125130000000
0!
0%
#125135000000
1!
1%
#125140000000
0!
0%
#125145000000
1!
1%
#125150000000
0!
0%
#125155000000
1!
1%
#125160000000
0!
0%
#125165000000
1!
1%
#125170000000
0!
0%
#125175000000
1!
1%
#125180000000
0!
0%
#125185000000
1!
1%
#125190000000
0!
0%
#125195000000
1!
1%
#125200000000
0!
0%
#125205000000
1!
1%
#125210000000
0!
0%
#125215000000
1!
1%
#125220000000
0!
0%
#125225000000
1!
1%
#125230000000
0!
0%
#125235000000
1!
1%
#125240000000
0!
0%
#125245000000
1!
1%
#125250000000
0!
0%
#125255000000
1!
1%
#125260000000
0!
0%
#125265000000
1!
1%
#125270000000
0!
0%
#125275000000
1!
1%
#125280000000
0!
0%
#125285000000
1!
1%
#125290000000
0!
0%
#125295000000
1!
1%
#125300000000
0!
0%
#125305000000
1!
1%
#125310000000
0!
0%
#125315000000
1!
1%
#125320000000
0!
0%
#125325000000
1!
1%
#125330000000
0!
0%
#125335000000
1!
1%
#125340000000
0!
0%
#125345000000
1!
1%
#125350000000
0!
0%
#125355000000
1!
1%
#125360000000
0!
0%
#125365000000
1!
1%
#125370000000
0!
0%
#125375000000
1!
1%
#125380000000
0!
0%
#125385000000
1!
1%
#125390000000
0!
0%
#125395000000
1!
1%
#125400000000
0!
0%
#125405000000
1!
1%
#125410000000
0!
0%
#125415000000
1!
1%
#125420000000
0!
0%
#125425000000
1!
1%
#125430000000
0!
0%
#125435000000
1!
1%
#125440000000
0!
0%
#125445000000
1!
1%
#125450000000
0!
0%
#125455000000
1!
1%
#125460000000
0!
0%
#125465000000
1!
1%
#125470000000
0!
0%
#125475000000
1!
1%
#125480000000
0!
0%
#125485000000
1!
1%
#125490000000
0!
0%
#125495000000
1!
1%
#125500000000
0!
0%
#125505000000
1!
1%
#125510000000
0!
0%
#125515000000
1!
1%
#125520000000
0!
0%
#125525000000
1!
1%
#125530000000
0!
0%
#125535000000
1!
1%
#125540000000
0!
0%
#125545000000
1!
1%
#125550000000
0!
0%
#125555000000
1!
1%
#125560000000
0!
0%
#125565000000
1!
1%
#125570000000
0!
0%
#125575000000
1!
1%
#125580000000
0!
0%
#125585000000
1!
1%
#125590000000
0!
0%
#125595000000
1!
1%
#125600000000
0!
0%
#125605000000
1!
1%
#125610000000
0!
0%
#125615000000
1!
1%
#125620000000
0!
0%
#125625000000
1!
1%
#125630000000
0!
0%
#125635000000
1!
1%
#125640000000
0!
0%
#125645000000
1!
1%
#125650000000
0!
0%
#125655000000
1!
1%
#125660000000
0!
0%
#125665000000
1!
1%
#125670000000
0!
0%
#125675000000
1!
1%
#125680000000
0!
0%
#125685000000
1!
1%
#125690000000
0!
0%
#125695000000
1!
1%
#125700000000
0!
0%
#125705000000
1!
1%
#125710000000
0!
0%
#125715000000
1!
1%
#125720000000
0!
0%
#125725000000
1!
1%
#125730000000
0!
0%
#125735000000
1!
1%
#125740000000
0!
0%
#125745000000
1!
1%
#125750000000
0!
0%
#125755000000
1!
1%
#125760000000
0!
0%
#125765000000
1!
1%
#125770000000
0!
0%
#125775000000
1!
1%
#125780000000
0!
0%
#125785000000
1!
1%
#125790000000
0!
0%
#125795000000
1!
1%
#125800000000
0!
0%
#125805000000
1!
1%
#125810000000
0!
0%
#125815000000
1!
1%
#125820000000
0!
0%
#125825000000
1!
1%
#125830000000
0!
0%
#125835000000
1!
1%
#125840000000
0!
0%
#125845000000
1!
1%
#125850000000
0!
0%
#125855000000
1!
1%
#125860000000
0!
0%
#125865000000
1!
1%
#125870000000
0!
0%
#125875000000
1!
1%
#125880000000
0!
0%
#125885000000
1!
1%
#125890000000
0!
0%
#125895000000
1!
1%
#125900000000
0!
0%
#125905000000
1!
1%
#125910000000
0!
0%
#125915000000
1!
1%
#125920000000
0!
0%
#125925000000
1!
1%
#125930000000
0!
0%
#125935000000
1!
1%
#125940000000
0!
0%
#125945000000
1!
1%
#125950000000
0!
0%
#125955000000
1!
1%
#125960000000
0!
0%
#125965000000
1!
1%
#125970000000
0!
0%
#125975000000
1!
1%
#125980000000
0!
0%
#125985000000
1!
1%
#125990000000
0!
0%
#125995000000
1!
1%
#126000000000
0!
0%
#126005000000
1!
1%
#126010000000
0!
0%
#126015000000
1!
1%
#126020000000
0!
0%
#126025000000
1!
1%
#126030000000
0!
0%
#126035000000
1!
1%
#126040000000
0!
0%
#126045000000
1!
1%
#126050000000
0!
0%
#126055000000
1!
1%
#126060000000
0!
0%
#126065000000
1!
1%
#126070000000
0!
0%
#126075000000
1!
1%
#126080000000
0!
0%
#126085000000
1!
1%
#126090000000
0!
0%
#126095000000
1!
1%
#126100000000
0!
0%
#126105000000
1!
1%
#126110000000
0!
0%
#126115000000
1!
1%
#126120000000
0!
0%
#126125000000
1!
1%
#126130000000
0!
0%
#126135000000
1!
1%
#126140000000
0!
0%
#126145000000
1!
1%
#126150000000
0!
0%
#126155000000
1!
1%
#126160000000
0!
0%
#126165000000
1!
1%
#126170000000
0!
0%
#126175000000
1!
1%
#126180000000
0!
0%
#126185000000
1!
1%
#126190000000
0!
0%
#126195000000
1!
1%
#126200000000
0!
0%
#126205000000
1!
1%
#126210000000
0!
0%
#126215000000
1!
1%
#126220000000
0!
0%
#126225000000
1!
1%
#126230000000
0!
0%
#126235000000
1!
1%
#126240000000
0!
0%
#126245000000
1!
1%
#126250000000
0!
0%
#126255000000
1!
1%
#126260000000
0!
0%
#126265000000
1!
1%
#126270000000
0!
0%
#126275000000
1!
1%
#126280000000
0!
0%
#126285000000
1!
1%
#126290000000
0!
0%
#126295000000
1!
1%
#126300000000
0!
0%
#126305000000
1!
1%
#126310000000
0!
0%
#126315000000
1!
1%
#126320000000
0!
0%
#126325000000
1!
1%
#126330000000
0!
0%
#126335000000
1!
1%
#126340000000
0!
0%
#126345000000
1!
1%
#126350000000
0!
0%
#126355000000
1!
1%
#126360000000
0!
0%
#126365000000
1!
1%
#126370000000
0!
0%
#126375000000
1!
1%
#126380000000
0!
0%
#126385000000
1!
1%
#126390000000
0!
0%
#126395000000
1!
1%
#126400000000
0!
0%
#126405000000
1!
1%
#126410000000
0!
0%
#126415000000
1!
1%
#126420000000
0!
0%
#126425000000
1!
1%
#126430000000
0!
0%
#126435000000
1!
1%
#126440000000
0!
0%
#126445000000
1!
1%
#126450000000
0!
0%
#126455000000
1!
1%
#126460000000
0!
0%
#126465000000
1!
1%
#126470000000
0!
0%
#126475000000
1!
1%
#126480000000
0!
0%
#126485000000
1!
1%
#126490000000
0!
0%
#126495000000
1!
1%
#126500000000
0!
0%
#126505000000
1!
1%
#126510000000
0!
0%
#126515000000
1!
1%
#126520000000
0!
0%
#126525000000
1!
1%
#126530000000
0!
0%
#126535000000
1!
1%
#126540000000
0!
0%
#126545000000
1!
1%
#126550000000
0!
0%
#126555000000
1!
1%
#126560000000
0!
0%
#126565000000
1!
1%
#126570000000
0!
0%
#126575000000
1!
1%
#126580000000
0!
0%
#126585000000
1!
1%
#126590000000
0!
0%
#126595000000
1!
1%
#126600000000
0!
0%
#126605000000
1!
1%
#126610000000
0!
0%
#126615000000
1!
1%
#126620000000
0!
0%
#126625000000
1!
1%
#126630000000
0!
0%
#126635000000
1!
1%
#126640000000
0!
0%
#126645000000
1!
1%
#126650000000
0!
0%
#126655000000
1!
1%
#126660000000
0!
0%
#126665000000
1!
1%
#126670000000
0!
0%
#126675000000
1!
1%
#126680000000
0!
0%
#126685000000
1!
1%
#126690000000
0!
0%
#126695000000
1!
1%
#126700000000
0!
0%
#126705000000
1!
1%
#126710000000
0!
0%
#126715000000
1!
1%
#126720000000
0!
0%
#126725000000
1!
1%
#126730000000
0!
0%
#126735000000
1!
1%
#126740000000
0!
0%
#126745000000
1!
1%
#126750000000
0!
0%
#126755000000
1!
1%
#126760000000
0!
0%
#126765000000
1!
1%
#126770000000
0!
0%
#126775000000
1!
1%
#126780000000
0!
0%
#126785000000
1!
1%
#126790000000
0!
0%
#126795000000
1!
1%
#126800000000
0!
0%
#126805000000
1!
1%
#126810000000
0!
0%
#126815000000
1!
1%
#126820000000
0!
0%
#126825000000
1!
1%
#126830000000
0!
0%
#126835000000
1!
1%
#126840000000
0!
0%
#126845000000
1!
1%
#126850000000
0!
0%
#126855000000
1!
1%
#126860000000
0!
0%
#126865000000
1!
1%
#126870000000
0!
0%
#126875000000
1!
1%
#126880000000
0!
0%
#126885000000
1!
1%
#126890000000
0!
0%
#126895000000
1!
1%
#126900000000
0!
0%
#126905000000
1!
1%
#126910000000
0!
0%
#126915000000
1!
1%
#126920000000
0!
0%
#126925000000
1!
1%
#126930000000
0!
0%
#126935000000
1!
1%
#126940000000
0!
0%
#126945000000
1!
1%
#126950000000
0!
0%
#126955000000
1!
1%
#126960000000
0!
0%
#126965000000
1!
1%
#126970000000
0!
0%
#126975000000
1!
1%
#126980000000
0!
0%
#126985000000
1!
1%
#126990000000
0!
0%
#126995000000
1!
1%
#127000000000
0!
0%
#127005000000
1!
1%
#127010000000
0!
0%
#127015000000
1!
1%
#127020000000
0!
0%
#127025000000
1!
1%
#127030000000
0!
0%
#127035000000
1!
1%
#127040000000
0!
0%
#127045000000
1!
1%
#127050000000
0!
0%
#127055000000
1!
1%
#127060000000
0!
0%
#127065000000
1!
1%
#127070000000
0!
0%
#127075000000
1!
1%
#127080000000
0!
0%
#127085000000
1!
1%
#127090000000
0!
0%
#127095000000
1!
1%
#127100000000
0!
0%
#127105000000
1!
1%
#127110000000
0!
0%
#127115000000
1!
1%
#127120000000
0!
0%
#127125000000
1!
1%
#127130000000
0!
0%
#127135000000
1!
1%
#127140000000
0!
0%
#127145000000
1!
1%
#127150000000
0!
0%
#127155000000
1!
1%
#127160000000
0!
0%
#127165000000
1!
1%
#127170000000
0!
0%
#127175000000
1!
1%
#127180000000
0!
0%
#127185000000
1!
1%
#127190000000
0!
0%
#127195000000
1!
1%
#127200000000
0!
0%
#127205000000
1!
1%
#127210000000
0!
0%
#127215000000
1!
1%
#127220000000
0!
0%
#127225000000
1!
1%
#127230000000
0!
0%
#127235000000
1!
1%
#127240000000
0!
0%
#127245000000
1!
1%
#127250000000
0!
0%
#127255000000
1!
1%
#127260000000
0!
0%
#127265000000
1!
1%
#127270000000
0!
0%
#127275000000
1!
1%
#127280000000
0!
0%
#127285000000
1!
1%
#127290000000
0!
0%
#127295000000
1!
1%
#127300000000
0!
0%
#127305000000
1!
1%
#127310000000
0!
0%
#127315000000
1!
1%
#127320000000
0!
0%
#127325000000
1!
1%
#127330000000
0!
0%
#127335000000
1!
1%
#127340000000
0!
0%
#127345000000
1!
1%
#127350000000
0!
0%
#127355000000
1!
1%
#127360000000
0!
0%
#127365000000
1!
1%
#127370000000
0!
0%
#127375000000
1!
1%
#127380000000
0!
0%
#127385000000
1!
1%
#127390000000
0!
0%
#127395000000
1!
1%
#127400000000
0!
0%
#127405000000
1!
1%
#127410000000
0!
0%
#127415000000
1!
1%
#127420000000
0!
0%
#127425000000
1!
1%
#127430000000
0!
0%
#127435000000
1!
1%
#127440000000
0!
0%
#127445000000
1!
1%
#127450000000
0!
0%
#127455000000
1!
1%
#127460000000
0!
0%
#127465000000
1!
1%
#127470000000
0!
0%
#127475000000
1!
1%
#127480000000
0!
0%
#127485000000
1!
1%
#127490000000
0!
0%
#127495000000
1!
1%
#127500000000
0!
0%
#127505000000
1!
1%
#127510000000
0!
0%
#127515000000
1!
1%
#127520000000
0!
0%
#127525000000
1!
1%
#127530000000
0!
0%
#127535000000
1!
1%
#127540000000
0!
0%
#127545000000
1!
1%
#127550000000
0!
0%
#127555000000
1!
1%
#127560000000
0!
0%
#127565000000
1!
1%
#127570000000
0!
0%
#127575000000
1!
1%
#127580000000
0!
0%
#127585000000
1!
1%
#127590000000
0!
0%
#127595000000
1!
1%
#127600000000
0!
0%
#127605000000
1!
1%
#127610000000
0!
0%
#127615000000
1!
1%
#127620000000
0!
0%
#127625000000
1!
1%
#127630000000
0!
0%
#127635000000
1!
1%
#127640000000
0!
0%
#127645000000
1!
1%
#127650000000
0!
0%
#127655000000
1!
1%
#127660000000
0!
0%
#127665000000
1!
1%
#127670000000
0!
0%
#127675000000
1!
1%
#127680000000
0!
0%
#127685000000
1!
1%
#127690000000
0!
0%
#127695000000
1!
1%
#127700000000
0!
0%
#127705000000
1!
1%
#127710000000
0!
0%
#127715000000
1!
1%
#127720000000
0!
0%
#127725000000
1!
1%
#127730000000
0!
0%
#127735000000
1!
1%
#127740000000
0!
0%
#127745000000
1!
1%
#127750000000
0!
0%
#127755000000
1!
1%
#127760000000
0!
0%
#127765000000
1!
1%
#127770000000
0!
0%
#127775000000
1!
1%
#127780000000
0!
0%
#127785000000
1!
1%
#127790000000
0!
0%
#127795000000
1!
1%
#127800000000
0!
0%
#127805000000
1!
1%
#127810000000
0!
0%
#127815000000
1!
1%
#127820000000
0!
0%
#127825000000
1!
1%
#127830000000
0!
0%
#127835000000
1!
1%
#127840000000
0!
0%
#127845000000
1!
1%
#127850000000
0!
0%
#127855000000
1!
1%
#127860000000
0!
0%
#127865000000
1!
1%
#127870000000
0!
0%
#127875000000
1!
1%
#127880000000
0!
0%
#127885000000
1!
1%
#127890000000
0!
0%
#127895000000
1!
1%
#127900000000
0!
0%
#127905000000
1!
1%
#127910000000
0!
0%
#127915000000
1!
1%
#127920000000
0!
0%
#127925000000
1!
1%
#127930000000
0!
0%
#127935000000
1!
1%
#127940000000
0!
0%
#127945000000
1!
1%
#127950000000
0!
0%
#127955000000
1!
1%
#127960000000
0!
0%
#127965000000
1!
1%
#127970000000
0!
0%
#127975000000
1!
1%
#127980000000
0!
0%
#127985000000
1!
1%
#127990000000
0!
0%
#127995000000
1!
1%
#128000000000
0!
0%
#128005000000
1!
1%
#128010000000
0!
0%
#128015000000
1!
1%
#128020000000
0!
0%
#128025000000
1!
1%
#128030000000
0!
0%
#128035000000
1!
1%
#128040000000
0!
0%
#128045000000
1!
1%
#128050000000
0!
0%
#128055000000
1!
1%
#128060000000
0!
0%
#128065000000
1!
1%
#128070000000
0!
0%
#128075000000
1!
1%
#128080000000
0!
0%
#128085000000
1!
1%
#128090000000
0!
0%
#128095000000
1!
1%
#128100000000
0!
0%
#128105000000
1!
1%
#128110000000
0!
0%
#128115000000
1!
1%
#128120000000
0!
0%
#128125000000
1!
1%
#128130000000
0!
0%
#128135000000
1!
1%
#128140000000
0!
0%
#128145000000
1!
1%
#128150000000
0!
0%
#128155000000
1!
1%
#128160000000
0!
0%
#128165000000
1!
1%
#128170000000
0!
0%
#128175000000
1!
1%
#128180000000
0!
0%
#128185000000
1!
1%
#128190000000
0!
0%
#128195000000
1!
1%
#128200000000
0!
0%
#128205000000
1!
1%
#128210000000
0!
0%
#128215000000
1!
1%
#128220000000
0!
0%
#128225000000
1!
1%
#128230000000
0!
0%
#128235000000
1!
1%
#128240000000
0!
0%
#128245000000
1!
1%
#128250000000
0!
0%
#128255000000
1!
1%
#128260000000
0!
0%
#128265000000
1!
1%
#128270000000
0!
0%
#128275000000
1!
1%
#128280000000
0!
0%
#128285000000
1!
1%
#128290000000
0!
0%
#128295000000
1!
1%
#128300000000
0!
0%
#128305000000
1!
1%
#128310000000
0!
0%
#128315000000
1!
1%
#128320000000
0!
0%
#128325000000
1!
1%
#128330000000
0!
0%
#128335000000
1!
1%
#128340000000
0!
0%
#128345000000
1!
1%
#128350000000
0!
0%
#128355000000
1!
1%
#128360000000
0!
0%
#128365000000
1!
1%
#128370000000
0!
0%
#128375000000
1!
1%
#128380000000
0!
0%
#128385000000
1!
1%
#128390000000
0!
0%
#128395000000
1!
1%
#128400000000
0!
0%
#128405000000
1!
1%
#128410000000
0!
0%
#128415000000
1!
1%
#128420000000
0!
0%
#128425000000
1!
1%
#128430000000
0!
0%
#128435000000
1!
1%
#128440000000
0!
0%
#128445000000
1!
1%
#128450000000
0!
0%
#128455000000
1!
1%
#128460000000
0!
0%
#128465000000
1!
1%
#128470000000
0!
0%
#128475000000
1!
1%
#128480000000
0!
0%
#128485000000
1!
1%
#128490000000
0!
0%
#128495000000
1!
1%
#128500000000
0!
0%
#128505000000
1!
1%
#128510000000
0!
0%
#128515000000
1!
1%
#128520000000
0!
0%
#128525000000
1!
1%
#128530000000
0!
0%
#128535000000
1!
1%
#128540000000
0!
0%
#128545000000
1!
1%
#128550000000
0!
0%
#128555000000
1!
1%
#128560000000
0!
0%
#128565000000
1!
1%
#128570000000
0!
0%
#128575000000
1!
1%
#128580000000
0!
0%
#128585000000
1!
1%
#128590000000
0!
0%
#128595000000
1!
1%
#128600000000
0!
0%
#128605000000
1!
1%
#128610000000
0!
0%
#128615000000
1!
1%
#128620000000
0!
0%
#128625000000
1!
1%
#128630000000
0!
0%
#128635000000
1!
1%
#128640000000
0!
0%
#128645000000
1!
1%
#128650000000
0!
0%
#128655000000
1!
1%
#128660000000
0!
0%
#128665000000
1!
1%
#128670000000
0!
0%
#128675000000
1!
1%
#128680000000
0!
0%
#128685000000
1!
1%
#128690000000
0!
0%
#128695000000
1!
1%
#128700000000
0!
0%
#128705000000
1!
1%
#128710000000
0!
0%
#128715000000
1!
1%
#128720000000
0!
0%
#128725000000
1!
1%
#128730000000
0!
0%
#128735000000
1!
1%
#128740000000
0!
0%
#128745000000
1!
1%
#128750000000
0!
0%
#128755000000
1!
1%
#128760000000
0!
0%
#128765000000
1!
1%
#128770000000
0!
0%
#128775000000
1!
1%
#128780000000
0!
0%
#128785000000
1!
1%
#128790000000
0!
0%
#128795000000
1!
1%
#128800000000
0!
0%
#128805000000
1!
1%
#128810000000
0!
0%
#128815000000
1!
1%
#128820000000
0!
0%
#128825000000
1!
1%
#128830000000
0!
0%
#128835000000
1!
1%
#128840000000
0!
0%
#128845000000
1!
1%
#128850000000
0!
0%
#128855000000
1!
1%
#128860000000
0!
0%
#128865000000
1!
1%
#128870000000
0!
0%
#128875000000
1!
1%
#128880000000
0!
0%
#128885000000
1!
1%
#128890000000
0!
0%
#128895000000
1!
1%
#128900000000
0!
0%
#128905000000
1!
1%
#128910000000
0!
0%
#128915000000
1!
1%
#128920000000
0!
0%
#128925000000
1!
1%
#128930000000
0!
0%
#128935000000
1!
1%
#128940000000
0!
0%
#128945000000
1!
1%
#128950000000
0!
0%
#128955000000
1!
1%
#128960000000
0!
0%
#128965000000
1!
1%
#128970000000
0!
0%
#128975000000
1!
1%
#128980000000
0!
0%
#128985000000
1!
1%
#128990000000
0!
0%
#128995000000
1!
1%
#129000000000
0!
0%
#129005000000
1!
1%
#129010000000
0!
0%
#129015000000
1!
1%
#129020000000
0!
0%
#129025000000
1!
1%
#129030000000
0!
0%
#129035000000
1!
1%
#129040000000
0!
0%
#129045000000
1!
1%
#129050000000
0!
0%
#129055000000
1!
1%
#129060000000
0!
0%
#129065000000
1!
1%
#129070000000
0!
0%
#129075000000
1!
1%
#129080000000
0!
0%
#129085000000
1!
1%
#129090000000
0!
0%
#129095000000
1!
1%
#129100000000
0!
0%
#129105000000
1!
1%
#129110000000
0!
0%
#129115000000
1!
1%
#129120000000
0!
0%
#129125000000
1!
1%
#129130000000
0!
0%
#129135000000
1!
1%
#129140000000
0!
0%
#129145000000
1!
1%
#129150000000
0!
0%
#129155000000
1!
1%
#129160000000
0!
0%
#129165000000
1!
1%
#129170000000
0!
0%
#129175000000
1!
1%
#129180000000
0!
0%
#129185000000
1!
1%
#129190000000
0!
0%
#129195000000
1!
1%
#129200000000
0!
0%
#129205000000
1!
1%
#129210000000
0!
0%
#129215000000
1!
1%
#129220000000
0!
0%
#129225000000
1!
1%
#129230000000
0!
0%
#129235000000
1!
1%
#129240000000
0!
0%
#129245000000
1!
1%
#129250000000
0!
0%
#129255000000
1!
1%
#129260000000
0!
0%
#129265000000
1!
1%
#129270000000
0!
0%
#129275000000
1!
1%
#129280000000
0!
0%
#129285000000
1!
1%
#129290000000
0!
0%
#129295000000
1!
1%
#129300000000
0!
0%
#129305000000
1!
1%
#129310000000
0!
0%
#129315000000
1!
1%
#129320000000
0!
0%
#129325000000
1!
1%
#129330000000
0!
0%
#129335000000
1!
1%
#129340000000
0!
0%
#129345000000
1!
1%
#129350000000
0!
0%
#129355000000
1!
1%
#129360000000
0!
0%
#129365000000
1!
1%
#129370000000
0!
0%
#129375000000
1!
1%
#129380000000
0!
0%
#129385000000
1!
1%
#129390000000
0!
0%
#129395000000
1!
1%
#129400000000
0!
0%
#129405000000
1!
1%
#129410000000
0!
0%
#129415000000
1!
1%
#129420000000
0!
0%
#129425000000
1!
1%
#129430000000
0!
0%
#129435000000
1!
1%
#129440000000
0!
0%
#129445000000
1!
1%
#129450000000
0!
0%
#129455000000
1!
1%
#129460000000
0!
0%
#129465000000
1!
1%
#129470000000
0!
0%
#129475000000
1!
1%
#129480000000
0!
0%
#129485000000
1!
1%
#129490000000
0!
0%
#129495000000
1!
1%
#129500000000
0!
0%
#129505000000
1!
1%
#129510000000
0!
0%
#129515000000
1!
1%
#129520000000
0!
0%
#129525000000
1!
1%
#129530000000
0!
0%
#129535000000
1!
1%
#129540000000
0!
0%
#129545000000
1!
1%
#129550000000
0!
0%
#129555000000
1!
1%
#129560000000
0!
0%
#129565000000
1!
1%
#129570000000
0!
0%
#129575000000
1!
1%
#129580000000
0!
0%
#129585000000
1!
1%
#129590000000
0!
0%
#129595000000
1!
1%
#129600000000
0!
0%
#129605000000
1!
1%
#129610000000
0!
0%
#129615000000
1!
1%
#129620000000
0!
0%
#129625000000
1!
1%
#129630000000
0!
0%
#129635000000
1!
1%
#129640000000
0!
0%
#129645000000
1!
1%
#129650000000
0!
0%
#129655000000
1!
1%
#129660000000
0!
0%
#129665000000
1!
1%
#129670000000
0!
0%
#129675000000
1!
1%
#129680000000
0!
0%
#129685000000
1!
1%
#129690000000
0!
0%
#129695000000
1!
1%
#129700000000
0!
0%
#129705000000
1!
1%
#129710000000
0!
0%
#129715000000
1!
1%
#129720000000
0!
0%
#129725000000
1!
1%
#129730000000
0!
0%
#129735000000
1!
1%
#129740000000
0!
0%
#129745000000
1!
1%
#129750000000
0!
0%
#129755000000
1!
1%
#129760000000
0!
0%
#129765000000
1!
1%
#129770000000
0!
0%
#129775000000
1!
1%
#129780000000
0!
0%
#129785000000
1!
1%
#129790000000
0!
0%
#129795000000
1!
1%
#129800000000
0!
0%
#129805000000
1!
1%
#129810000000
0!
0%
#129815000000
1!
1%
#129820000000
0!
0%
#129825000000
1!
1%
#129830000000
0!
0%
#129835000000
1!
1%
#129840000000
0!
0%
#129845000000
1!
1%
#129850000000
0!
0%
#129855000000
1!
1%
#129860000000
0!
0%
#129865000000
1!
1%
#129870000000
0!
0%
#129875000000
1!
1%
#129880000000
0!
0%
#129885000000
1!
1%
#129890000000
0!
0%
#129895000000
1!
1%
#129900000000
0!
0%
#129905000000
1!
1%
#129910000000
0!
0%
#129915000000
1!
1%
#129920000000
0!
0%
#129925000000
1!
1%
#129930000000
0!
0%
#129935000000
1!
1%
#129940000000
0!
0%
#129945000000
1!
1%
#129950000000
0!
0%
#129955000000
1!
1%
#129960000000
0!
0%
#129965000000
1!
1%
#129970000000
0!
0%
#129975000000
1!
1%
#129980000000
0!
0%
#129985000000
1!
1%
#129990000000
0!
0%
#129995000000
1!
1%
#130000000000
0!
0%
#130005000000
1!
1%
#130010000000
0!
0%
#130015000000
1!
1%
#130020000000
0!
0%
#130025000000
1!
1%
#130030000000
0!
0%
#130035000000
1!
1%
#130040000000
0!
0%
#130045000000
1!
1%
#130050000000
0!
0%
#130055000000
1!
1%
#130060000000
0!
0%
#130065000000
1!
1%
#130070000000
0!
0%
#130075000000
1!
1%
#130080000000
0!
0%
#130085000000
1!
1%
#130090000000
0!
0%
#130095000000
1!
1%
#130100000000
0!
0%
#130105000000
1!
1%
#130110000000
0!
0%
#130115000000
1!
1%
#130120000000
0!
0%
#130125000000
1!
1%
#130130000000
0!
0%
#130135000000
1!
1%
#130140000000
0!
0%
#130145000000
1!
1%
#130150000000
0!
0%
#130155000000
1!
1%
#130160000000
0!
0%
#130165000000
1!
1%
#130170000000
0!
0%
#130175000000
1!
1%
#130180000000
0!
0%
#130185000000
1!
1%
#130190000000
0!
0%
#130195000000
1!
1%
#130200000000
0!
0%
#130205000000
1!
1%
#130210000000
0!
0%
#130215000000
1!
1%
#130220000000
0!
0%
#130225000000
1!
1%
#130230000000
0!
0%
#130235000000
1!
1%
#130240000000
0!
0%
#130245000000
1!
1%
#130250000000
0!
0%
#130255000000
1!
1%
#130260000000
0!
0%
#130265000000
1!
1%
#130270000000
0!
0%
#130275000000
1!
1%
#130280000000
0!
0%
#130285000000
1!
1%
#130290000000
0!
0%
#130295000000
1!
1%
#130300000000
0!
0%
#130305000000
1!
1%
#130310000000
0!
0%
#130315000000
1!
1%
#130320000000
0!
0%
#130325000000
1!
1%
#130330000000
0!
0%
#130335000000
1!
1%
#130340000000
0!
0%
#130345000000
1!
1%
#130350000000
0!
0%
#130355000000
1!
1%
#130360000000
0!
0%
#130365000000
1!
1%
#130370000000
0!
0%
#130375000000
1!
1%
#130380000000
0!
0%
#130385000000
1!
1%
#130390000000
0!
0%
#130395000000
1!
1%
#130400000000
0!
0%
#130405000000
1!
1%
#130410000000
0!
0%
#130415000000
1!
1%
#130420000000
0!
0%
#130425000000
1!
1%
#130430000000
0!
0%
#130435000000
1!
1%
#130440000000
0!
0%
#130445000000
1!
1%
#130450000000
0!
0%
#130455000000
1!
1%
#130460000000
0!
0%
#130465000000
1!
1%
#130470000000
0!
0%
#130475000000
1!
1%
#130480000000
0!
0%
#130485000000
1!
1%
#130490000000
0!
0%
#130495000000
1!
1%
#130500000000
0!
0%
#130505000000
1!
1%
#130510000000
0!
0%
#130515000000
1!
1%
#130520000000
0!
0%
#130525000000
1!
1%
#130530000000
0!
0%
#130535000000
1!
1%
#130540000000
0!
0%
#130545000000
1!
1%
#130550000000
0!
0%
#130555000000
1!
1%
#130560000000
0!
0%
#130565000000
1!
1%
#130570000000
0!
0%
#130575000000
1!
1%
#130580000000
0!
0%
#130585000000
1!
1%
#130590000000
0!
0%
#130595000000
1!
1%
#130600000000
0!
0%
#130605000000
1!
1%
#130610000000
0!
0%
#130615000000
1!
1%
#130620000000
0!
0%
#130625000000
1!
1%
#130630000000
0!
0%
#130635000000
1!
1%
#130640000000
0!
0%
#130645000000
1!
1%
#130650000000
0!
0%
#130655000000
1!
1%
#130660000000
0!
0%
#130665000000
1!
1%
#130670000000
0!
0%
#130675000000
1!
1%
#130680000000
0!
0%
#130685000000
1!
1%
#130690000000
0!
0%
#130695000000
1!
1%
#130700000000
0!
0%
#130705000000
1!
1%
#130710000000
0!
0%
#130715000000
1!
1%
#130720000000
0!
0%
#130725000000
1!
1%
#130730000000
0!
0%
#130735000000
1!
1%
#130740000000
0!
0%
#130745000000
1!
1%
#130750000000
0!
0%
#130755000000
1!
1%
#130760000000
0!
0%
#130765000000
1!
1%
#130770000000
0!
0%
#130775000000
1!
1%
#130780000000
0!
0%
#130785000000
1!
1%
#130790000000
0!
0%
#130795000000
1!
1%
#130800000000
0!
0%
#130805000000
1!
1%
#130810000000
0!
0%
#130815000000
1!
1%
#130820000000
0!
0%
#130825000000
1!
1%
#130830000000
0!
0%
#130835000000
1!
1%
#130840000000
0!
0%
#130845000000
1!
1%
#130850000000
0!
0%
#130855000000
1!
1%
#130860000000
0!
0%
#130865000000
1!
1%
#130870000000
0!
0%
#130875000000
1!
1%
#130880000000
0!
0%
#130885000000
1!
1%
#130890000000
0!
0%
#130895000000
1!
1%
#130900000000
0!
0%
#130905000000
1!
1%
#130910000000
0!
0%
#130915000000
1!
1%
#130920000000
0!
0%
#130925000000
1!
1%
#130930000000
0!
0%
#130935000000
1!
1%
#130940000000
0!
0%
#130945000000
1!
1%
#130950000000
0!
0%
#130955000000
1!
1%
#130960000000
0!
0%
#130965000000
1!
1%
#130970000000
0!
0%
#130975000000
1!
1%
#130980000000
0!
0%
#130985000000
1!
1%
#130990000000
0!
0%
#130995000000
1!
1%
#131000000000
0!
0%
#131005000000
1!
1%
#131010000000
0!
0%
#131015000000
1!
1%
#131020000000
0!
0%
#131025000000
1!
1%
#131030000000
0!
0%
#131035000000
1!
1%
#131040000000
0!
0%
#131045000000
1!
1%
#131050000000
0!
0%
#131055000000
1!
1%
#131060000000
0!
0%
#131065000000
1!
1%
#131070000000
0!
0%
#131075000000
1!
1%
#131080000000
0!
0%
#131085000000
1!
1%
#131090000000
0!
0%
#131095000000
1!
1%
#131100000000
0!
0%
#131105000000
1!
1%
#131110000000
0!
0%
#131115000000
1!
1%
#131120000000
0!
0%
#131125000000
1!
1%
#131130000000
0!
0%
#131135000000
1!
1%
#131140000000
0!
0%
#131145000000
1!
1%
#131150000000
0!
0%
#131155000000
1!
1%
#131160000000
0!
0%
#131165000000
1!
1%
#131170000000
0!
0%
#131175000000
1!
1%
#131180000000
0!
0%
#131185000000
1!
1%
#131190000000
0!
0%
#131195000000
1!
1%
#131200000000
0!
0%
#131205000000
1!
1%
#131210000000
0!
0%
#131215000000
1!
1%
#131220000000
0!
0%
#131225000000
1!
1%
#131230000000
0!
0%
#131235000000
1!
1%
#131240000000
0!
0%
#131245000000
1!
1%
#131250000000
0!
0%
#131255000000
1!
1%
#131260000000
0!
0%
#131265000000
1!
1%
#131270000000
0!
0%
#131275000000
1!
1%
#131280000000
0!
0%
#131285000000
1!
1%
#131290000000
0!
0%
#131295000000
1!
1%
#131300000000
0!
0%
#131305000000
1!
1%
#131310000000
0!
0%
#131315000000
1!
1%
#131320000000
0!
0%
#131325000000
1!
1%
#131330000000
0!
0%
#131335000000
1!
1%
#131340000000
0!
0%
#131345000000
1!
1%
#131350000000
0!
0%
#131355000000
1!
1%
#131360000000
0!
0%
#131365000000
1!
1%
#131370000000
0!
0%
#131375000000
1!
1%
#131380000000
0!
0%
#131385000000
1!
1%
#131390000000
0!
0%
#131395000000
1!
1%
#131400000000
0!
0%
#131405000000
1!
1%
#131410000000
0!
0%
#131415000000
1!
1%
#131420000000
0!
0%
#131425000000
1!
1%
#131430000000
0!
0%
#131435000000
1!
1%
#131440000000
0!
0%
#131445000000
1!
1%
#131450000000
0!
0%
#131455000000
1!
1%
#131460000000
0!
0%
#131465000000
1!
1%
#131470000000
0!
0%
#131475000000
1!
1%
#131480000000
0!
0%
#131485000000
1!
1%
#131490000000
0!
0%
#131495000000
1!
1%
#131500000000
0!
0%
#131505000000
1!
1%
#131510000000
0!
0%
#131515000000
1!
1%
#131520000000
0!
0%
#131525000000
1!
1%
#131530000000
0!
0%
#131535000000
1!
1%
#131540000000
0!
0%
#131545000000
1!
1%
#131550000000
0!
0%
#131555000000
1!
1%
#131560000000
0!
0%
#131565000000
1!
1%
#131570000000
0!
0%
#131575000000
1!
1%
#131580000000
0!
0%
#131585000000
1!
1%
#131590000000
0!
0%
#131595000000
1!
1%
#131600000000
0!
0%
#131605000000
1!
1%
#131610000000
0!
0%
#131615000000
1!
1%
#131620000000
0!
0%
#131625000000
1!
1%
#131630000000
0!
0%
#131635000000
1!
1%
#131640000000
0!
0%
#131645000000
1!
1%
#131650000000
0!
0%
#131655000000
1!
1%
#131660000000
0!
0%
#131665000000
1!
1%
#131670000000
0!
0%
#131675000000
1!
1%
#131680000000
0!
0%
#131685000000
1!
1%
#131690000000
0!
0%
#131695000000
1!
1%
#131700000000
0!
0%
#131705000000
1!
1%
#131710000000
0!
0%
#131715000000
1!
1%
#131720000000
0!
0%
#131725000000
1!
1%
#131730000000
0!
0%
#131735000000
1!
1%
#131740000000
0!
0%
#131745000000
1!
1%
#131750000000
0!
0%
#131755000000
1!
1%
#131760000000
0!
0%
#131765000000
1!
1%
#131770000000
0!
0%
#131775000000
1!
1%
#131780000000
0!
0%
#131785000000
1!
1%
#131790000000
0!
0%
#131795000000
1!
1%
#131800000000
0!
0%
#131805000000
1!
1%
#131810000000
0!
0%
#131815000000
1!
1%
#131820000000
0!
0%
#131825000000
1!
1%
#131830000000
0!
0%
#131835000000
1!
1%
#131840000000
0!
0%
#131845000000
1!
1%
#131850000000
0!
0%
#131855000000
1!
1%
#131860000000
0!
0%
#131865000000
1!
1%
#131870000000
0!
0%
#131875000000
1!
1%
#131880000000
0!
0%
#131885000000
1!
1%
#131890000000
0!
0%
#131895000000
1!
1%
#131900000000
0!
0%
#131905000000
1!
1%
#131910000000
0!
0%
#131915000000
1!
1%
#131920000000
0!
0%
#131925000000
1!
1%
#131930000000
0!
0%
#131935000000
1!
1%
#131940000000
0!
0%
#131945000000
1!
1%
#131950000000
0!
0%
#131955000000
1!
1%
#131960000000
0!
0%
#131965000000
1!
1%
#131970000000
0!
0%
#131975000000
1!
1%
#131980000000
0!
0%
#131985000000
1!
1%
#131990000000
0!
0%
#131995000000
1!
1%
#132000000000
0!
0%
#132005000000
1!
1%
#132010000000
0!
0%
#132015000000
1!
1%
#132020000000
0!
0%
#132025000000
1!
1%
#132030000000
0!
0%
#132035000000
1!
1%
#132040000000
0!
0%
#132045000000
1!
1%
#132050000000
0!
0%
#132055000000
1!
1%
#132060000000
0!
0%
#132065000000
1!
1%
#132070000000
0!
0%
#132075000000
1!
1%
#132080000000
0!
0%
#132085000000
1!
1%
#132090000000
0!
0%
#132095000000
1!
1%
#132100000000
0!
0%
#132105000000
1!
1%
#132110000000
0!
0%
#132115000000
1!
1%
#132120000000
0!
0%
#132125000000
1!
1%
#132130000000
0!
0%
#132135000000
1!
1%
#132140000000
0!
0%
#132145000000
1!
1%
#132150000000
0!
0%
#132155000000
1!
1%
#132160000000
0!
0%
#132165000000
1!
1%
#132170000000
0!
0%
#132175000000
1!
1%
#132180000000
0!
0%
#132185000000
1!
1%
#132190000000
0!
0%
#132195000000
1!
1%
#132200000000
0!
0%
#132205000000
1!
1%
#132210000000
0!
0%
#132215000000
1!
1%
#132220000000
0!
0%
#132225000000
1!
1%
#132230000000
0!
0%
#132235000000
1!
1%
#132240000000
0!
0%
#132245000000
1!
1%
#132250000000
0!
0%
#132255000000
1!
1%
#132260000000
0!
0%
#132265000000
1!
1%
#132270000000
0!
0%
#132275000000
1!
1%
#132280000000
0!
0%
#132285000000
1!
1%
#132290000000
0!
0%
#132295000000
1!
1%
#132300000000
0!
0%
#132305000000
1!
1%
#132310000000
0!
0%
#132315000000
1!
1%
#132320000000
0!
0%
#132325000000
1!
1%
#132330000000
0!
0%
#132335000000
1!
1%
#132340000000
0!
0%
#132345000000
1!
1%
#132350000000
0!
0%
#132355000000
1!
1%
#132360000000
0!
0%
#132365000000
1!
1%
#132370000000
0!
0%
#132375000000
1!
1%
#132380000000
0!
0%
#132385000000
1!
1%
#132390000000
0!
0%
#132395000000
1!
1%
#132400000000
0!
0%
#132405000000
1!
1%
#132410000000
0!
0%
#132415000000
1!
1%
#132420000000
0!
0%
#132425000000
1!
1%
#132430000000
0!
0%
#132435000000
1!
1%
#132440000000
0!
0%
#132445000000
1!
1%
#132450000000
0!
0%
#132455000000
1!
1%
#132460000000
0!
0%
#132465000000
1!
1%
#132470000000
0!
0%
#132475000000
1!
1%
#132480000000
0!
0%
#132485000000
1!
1%
#132490000000
0!
0%
#132495000000
1!
1%
#132500000000
0!
0%
#132505000000
1!
1%
#132510000000
0!
0%
#132515000000
1!
1%
#132520000000
0!
0%
#132525000000
1!
1%
#132530000000
0!
0%
#132535000000
1!
1%
#132540000000
0!
0%
#132545000000
1!
1%
#132550000000
0!
0%
#132555000000
1!
1%
#132560000000
0!
0%
#132565000000
1!
1%
#132570000000
0!
0%
#132575000000
1!
1%
#132580000000
0!
0%
#132585000000
1!
1%
#132590000000
0!
0%
#132595000000
1!
1%
#132600000000
0!
0%
#132605000000
1!
1%
#132610000000
0!
0%
#132615000000
1!
1%
#132620000000
0!
0%
#132625000000
1!
1%
#132630000000
0!
0%
#132635000000
1!
1%
#132640000000
0!
0%
#132645000000
1!
1%
#132650000000
0!
0%
#132655000000
1!
1%
#132660000000
0!
0%
#132665000000
1!
1%
#132670000000
0!
0%
#132675000000
1!
1%
#132680000000
0!
0%
#132685000000
1!
1%
#132690000000
0!
0%
#132695000000
1!
1%
#132700000000
0!
0%
#132705000000
1!
1%
#132710000000
0!
0%
#132715000000
1!
1%
#132720000000
0!
0%
#132725000000
1!
1%
#132730000000
0!
0%
#132735000000
1!
1%
#132740000000
0!
0%
#132745000000
1!
1%
#132750000000
0!
0%
#132755000000
1!
1%
#132760000000
0!
0%
#132765000000
1!
1%
#132770000000
0!
0%
#132775000000
1!
1%
#132780000000
0!
0%
#132785000000
1!
1%
#132790000000
0!
0%
#132795000000
1!
1%
#132800000000
0!
0%
#132805000000
1!
1%
#132810000000
0!
0%
#132815000000
1!
1%
#132820000000
0!
0%
#132825000000
1!
1%
#132830000000
0!
0%
#132835000000
1!
1%
#132840000000
0!
0%
#132845000000
1!
1%
#132850000000
0!
0%
#132855000000
1!
1%
#132860000000
0!
0%
#132865000000
1!
1%
#132870000000
0!
0%
#132875000000
1!
1%
#132880000000
0!
0%
#132885000000
1!
1%
#132890000000
0!
0%
#132895000000
1!
1%
#132900000000
0!
0%
#132905000000
1!
1%
#132910000000
0!
0%
#132915000000
1!
1%
#132920000000
0!
0%
#132925000000
1!
1%
#132930000000
0!
0%
#132935000000
1!
1%
#132940000000
0!
0%
#132945000000
1!
1%
#132950000000
0!
0%
#132955000000
1!
1%
#132960000000
0!
0%
#132965000000
1!
1%
#132970000000
0!
0%
#132975000000
1!
1%
#132980000000
0!
0%
#132985000000
1!
1%
#132990000000
0!
0%
#132995000000
1!
1%
#133000000000
0!
0%
#133005000000
1!
1%
#133010000000
0!
0%
#133015000000
1!
1%
#133020000000
0!
0%
#133025000000
1!
1%
#133030000000
0!
0%
#133035000000
1!
1%
#133040000000
0!
0%
#133045000000
1!
1%
#133050000000
0!
0%
#133055000000
1!
1%
#133060000000
0!
0%
#133065000000
1!
1%
#133070000000
0!
0%
#133075000000
1!
1%
#133080000000
0!
0%
#133085000000
1!
1%
#133090000000
0!
0%
#133095000000
1!
1%
#133100000000
0!
0%
#133105000000
1!
1%
#133110000000
0!
0%
#133115000000
1!
1%
#133120000000
0!
0%
#133125000000
1!
1%
#133130000000
0!
0%
#133135000000
1!
1%
#133140000000
0!
0%
#133145000000
1!
1%
#133150000000
0!
0%
#133155000000
1!
1%
#133160000000
0!
0%
#133165000000
1!
1%
#133170000000
0!
0%
#133175000000
1!
1%
#133180000000
0!
0%
#133185000000
1!
1%
#133190000000
0!
0%
#133195000000
1!
1%
#133200000000
0!
0%
#133205000000
1!
1%
#133210000000
0!
0%
#133215000000
1!
1%
#133220000000
0!
0%
#133225000000
1!
1%
#133230000000
0!
0%
#133235000000
1!
1%
#133240000000
0!
0%
#133245000000
1!
1%
#133250000000
0!
0%
#133255000000
1!
1%
#133260000000
0!
0%
#133265000000
1!
1%
#133270000000
0!
0%
#133275000000
1!
1%
#133280000000
0!
0%
#133285000000
1!
1%
#133290000000
0!
0%
#133295000000
1!
1%
#133300000000
0!
0%
#133305000000
1!
1%
#133310000000
0!
0%
#133315000000
1!
1%
#133320000000
0!
0%
#133325000000
1!
1%
#133330000000
0!
0%
#133335000000
1!
1%
#133340000000
0!
0%
#133345000000
1!
1%
#133350000000
0!
0%
#133355000000
1!
1%
#133360000000
0!
0%
#133365000000
1!
1%
#133370000000
0!
0%
#133375000000
1!
1%
#133380000000
0!
0%
#133385000000
1!
1%
#133390000000
0!
0%
#133395000000
1!
1%
#133400000000
0!
0%
#133405000000
1!
1%
#133410000000
0!
0%
#133415000000
1!
1%
#133420000000
0!
0%
#133425000000
1!
1%
#133430000000
0!
0%
#133435000000
1!
1%
#133440000000
0!
0%
#133445000000
1!
1%
#133450000000
0!
0%
#133455000000
1!
1%
#133460000000
0!
0%
#133465000000
1!
1%
#133470000000
0!
0%
#133475000000
1!
1%
#133480000000
0!
0%
#133485000000
1!
1%
#133490000000
0!
0%
#133495000000
1!
1%
#133500000000
0!
0%
#133505000000
1!
1%
#133510000000
0!
0%
#133515000000
1!
1%
#133520000000
0!
0%
#133525000000
1!
1%
#133530000000
0!
0%
#133535000000
1!
1%
#133540000000
0!
0%
#133545000000
1!
1%
#133550000000
0!
0%
#133555000000
1!
1%
#133560000000
0!
0%
#133565000000
1!
1%
#133570000000
0!
0%
#133575000000
1!
1%
#133580000000
0!
0%
#133585000000
1!
1%
#133590000000
0!
0%
#133595000000
1!
1%
#133600000000
0!
0%
#133605000000
1!
1%
#133610000000
0!
0%
#133615000000
1!
1%
#133620000000
0!
0%
#133625000000
1!
1%
#133630000000
0!
0%
#133635000000
1!
1%
#133640000000
0!
0%
#133645000000
1!
1%
#133650000000
0!
0%
#133655000000
1!
1%
#133660000000
0!
0%
#133665000000
1!
1%
#133670000000
0!
0%
#133675000000
1!
1%
#133680000000
0!
0%
#133685000000
1!
1%
#133690000000
0!
0%
#133695000000
1!
1%
#133700000000
0!
0%
#133705000000
1!
1%
#133710000000
0!
0%
#133715000000
1!
1%
#133720000000
0!
0%
#133725000000
1!
1%
#133730000000
0!
0%
#133735000000
1!
1%
#133740000000
0!
0%
#133745000000
1!
1%
#133750000000
0!
0%
#133755000000
1!
1%
#133760000000
0!
0%
#133765000000
1!
1%
#133770000000
0!
0%
#133775000000
1!
1%
#133780000000
0!
0%
#133785000000
1!
1%
#133790000000
0!
0%
#133795000000
1!
1%
#133800000000
0!
0%
#133805000000
1!
1%
#133810000000
0!
0%
#133815000000
1!
1%
#133820000000
0!
0%
#133825000000
1!
1%
#133830000000
0!
0%
#133835000000
1!
1%
#133840000000
0!
0%
#133845000000
1!
1%
#133850000000
0!
0%
#133855000000
1!
1%
#133860000000
0!
0%
#133865000000
1!
1%
#133870000000
0!
0%
#133875000000
1!
1%
#133880000000
0!
0%
#133885000000
1!
1%
#133890000000
0!
0%
#133895000000
1!
1%
#133900000000
0!
0%
#133905000000
1!
1%
#133910000000
0!
0%
#133915000000
1!
1%
#133920000000
0!
0%
#133925000000
1!
1%
#133930000000
0!
0%
#133935000000
1!
1%
#133940000000
0!
0%
#133945000000
1!
1%
#133950000000
0!
0%
#133955000000
1!
1%
#133960000000
0!
0%
#133965000000
1!
1%
#133970000000
0!
0%
#133975000000
1!
1%
#133980000000
0!
0%
#133985000000
1!
1%
#133990000000
0!
0%
#133995000000
1!
1%
#134000000000
0!
0%
#134005000000
1!
1%
#134010000000
0!
0%
#134015000000
1!
1%
#134020000000
0!
0%
#134025000000
1!
1%
#134030000000
0!
0%
#134035000000
1!
1%
#134040000000
0!
0%
#134045000000
1!
1%
#134050000000
0!
0%
#134055000000
1!
1%
#134060000000
0!
0%
#134065000000
1!
1%
#134070000000
0!
0%
#134075000000
1!
1%
#134080000000
0!
0%
#134085000000
1!
1%
#134090000000
0!
0%
#134095000000
1!
1%
#134100000000
0!
0%
#134105000000
1!
1%
#134110000000
0!
0%
#134115000000
1!
1%
#134120000000
0!
0%
#134125000000
1!
1%
#134130000000
0!
0%
#134135000000
1!
1%
#134140000000
0!
0%
#134145000000
1!
1%
#134150000000
0!
0%
#134155000000
1!
1%
#134160000000
0!
0%
#134165000000
1!
1%
#134170000000
0!
0%
#134175000000
1!
1%
#134180000000
0!
0%
#134185000000
1!
1%
#134190000000
0!
0%
#134195000000
1!
1%
#134200000000
0!
0%
#134205000000
1!
1%
#134210000000
0!
0%
#134215000000
1!
1%
#134220000000
0!
0%
#134225000000
1!
1%
#134230000000
0!
0%
#134235000000
1!
1%
#134240000000
0!
0%
#134245000000
1!
1%
#134250000000
0!
0%
#134255000000
1!
1%
#134260000000
0!
0%
#134265000000
1!
1%
#134270000000
0!
0%
#134275000000
1!
1%
#134280000000
0!
0%
#134285000000
1!
1%
#134290000000
0!
0%
#134295000000
1!
1%
#134300000000
0!
0%
#134305000000
1!
1%
#134310000000
0!
0%
#134315000000
1!
1%
#134320000000
0!
0%
#134325000000
1!
1%
#134330000000
0!
0%
#134335000000
1!
1%
#134340000000
0!
0%
#134345000000
1!
1%
#134350000000
0!
0%
#134355000000
1!
1%
#134360000000
0!
0%
#134365000000
1!
1%
#134370000000
0!
0%
#134375000000
1!
1%
#134380000000
0!
0%
#134385000000
1!
1%
#134390000000
0!
0%
#134395000000
1!
1%
#134400000000
0!
0%
#134405000000
1!
1%
#134410000000
0!
0%
#134415000000
1!
1%
#134420000000
0!
0%
#134425000000
1!
1%
#134430000000
0!
0%
#134435000000
1!
1%
#134440000000
0!
0%
#134445000000
1!
1%
#134450000000
0!
0%
#134455000000
1!
1%
#134460000000
0!
0%
#134465000000
1!
1%
#134470000000
0!
0%
#134475000000
1!
1%
#134480000000
0!
0%
#134485000000
1!
1%
#134490000000
0!
0%
#134495000000
1!
1%
#134500000000
0!
0%
#134505000000
1!
1%
#134510000000
0!
0%
#134515000000
1!
1%
#134520000000
0!
0%
#134525000000
1!
1%
#134530000000
0!
0%
#134535000000
1!
1%
#134540000000
0!
0%
#134545000000
1!
1%
#134550000000
0!
0%
#134555000000
1!
1%
#134560000000
0!
0%
#134565000000
1!
1%
#134570000000
0!
0%
#134575000000
1!
1%
#134580000000
0!
0%
#134585000000
1!
1%
#134590000000
0!
0%
#134595000000
1!
1%
#134600000000
0!
0%
#134605000000
1!
1%
#134610000000
0!
0%
#134615000000
1!
1%
#134620000000
0!
0%
#134625000000
1!
1%
#134630000000
0!
0%
#134635000000
1!
1%
#134640000000
0!
0%
#134645000000
1!
1%
#134650000000
0!
0%
#134655000000
1!
1%
#134660000000
0!
0%
#134665000000
1!
1%
#134670000000
0!
0%
#134675000000
1!
1%
#134680000000
0!
0%
#134685000000
1!
1%
#134690000000
0!
0%
#134695000000
1!
1%
#134700000000
0!
0%
#134705000000
1!
1%
#134710000000
0!
0%
#134715000000
1!
1%
#134720000000
0!
0%
#134725000000
1!
1%
#134730000000
0!
0%
#134735000000
1!
1%
#134740000000
0!
0%
#134745000000
1!
1%
#134750000000
0!
0%
#134755000000
1!
1%
#134760000000
0!
0%
#134765000000
1!
1%
#134770000000
0!
0%
#134775000000
1!
1%
#134780000000
0!
0%
#134785000000
1!
1%
#134790000000
0!
0%
#134795000000
1!
1%
#134800000000
0!
0%
#134805000000
1!
1%
#134810000000
0!
0%
#134815000000
1!
1%
#134820000000
0!
0%
#134825000000
1!
1%
#134830000000
0!
0%
#134835000000
1!
1%
#134840000000
0!
0%
#134845000000
1!
1%
#134850000000
0!
0%
#134855000000
1!
1%
#134860000000
0!
0%
#134865000000
1!
1%
#134870000000
0!
0%
#134875000000
1!
1%
#134880000000
0!
0%
#134885000000
1!
1%
#134890000000
0!
0%
#134895000000
1!
1%
#134900000000
0!
0%
#134905000000
1!
1%
#134910000000
0!
0%
#134915000000
1!
1%
#134920000000
0!
0%
#134925000000
1!
1%
#134930000000
0!
0%
#134935000000
1!
1%
#134940000000
0!
0%
#134945000000
1!
1%
#134950000000
0!
0%
#134955000000
1!
1%
#134960000000
0!
0%
#134965000000
1!
1%
#134970000000
0!
0%
#134975000000
1!
1%
#134980000000
0!
0%
#134985000000
1!
1%
#134990000000
0!
0%
#134995000000
1!
1%
#135000000000
0!
0%
#135005000000
1!
1%
#135010000000
0!
0%
#135015000000
1!
1%
#135020000000
0!
0%
#135025000000
1!
1%
#135030000000
0!
0%
#135035000000
1!
1%
#135040000000
0!
0%
#135045000000
1!
1%
#135050000000
0!
0%
#135055000000
1!
1%
#135060000000
0!
0%
#135065000000
1!
1%
#135070000000
0!
0%
#135075000000
1!
1%
#135080000000
0!
0%
#135085000000
1!
1%
#135090000000
0!
0%
#135095000000
1!
1%
#135100000000
0!
0%
#135105000000
1!
1%
#135110000000
0!
0%
#135115000000
1!
1%
#135120000000
0!
0%
#135125000000
1!
1%
#135130000000
0!
0%
#135135000000
1!
1%
#135140000000
0!
0%
#135145000000
1!
1%
#135150000000
0!
0%
#135155000000
1!
1%
#135160000000
0!
0%
#135165000000
1!
1%
#135170000000
0!
0%
#135175000000
1!
1%
#135180000000
0!
0%
#135185000000
1!
1%
#135190000000
0!
0%
#135195000000
1!
1%
#135200000000
0!
0%
#135205000000
1!
1%
#135210000000
0!
0%
#135215000000
1!
1%
#135220000000
0!
0%
#135225000000
1!
1%
#135230000000
0!
0%
#135235000000
1!
1%
#135240000000
0!
0%
#135245000000
1!
1%
#135250000000
0!
0%
#135255000000
1!
1%
#135260000000
0!
0%
#135265000000
1!
1%
#135270000000
0!
0%
#135275000000
1!
1%
#135280000000
0!
0%
#135285000000
1!
1%
#135290000000
0!
0%
#135295000000
1!
1%
#135300000000
0!
0%
#135305000000
1!
1%
#135310000000
0!
0%
#135315000000
1!
1%
#135320000000
0!
0%
#135325000000
1!
1%
#135330000000
0!
0%
#135335000000
1!
1%
#135340000000
0!
0%
#135345000000
1!
1%
#135350000000
0!
0%
#135355000000
1!
1%
#135360000000
0!
0%
#135365000000
1!
1%
#135370000000
0!
0%
#135375000000
1!
1%
#135380000000
0!
0%
#135385000000
1!
1%
#135390000000
0!
0%
#135395000000
1!
1%
#135400000000
0!
0%
#135405000000
1!
1%
#135410000000
0!
0%
#135415000000
1!
1%
#135420000000
0!
0%
#135425000000
1!
1%
#135430000000
0!
0%
#135435000000
1!
1%
#135440000000
0!
0%
#135445000000
1!
1%
#135450000000
0!
0%
#135455000000
1!
1%
#135460000000
0!
0%
#135465000000
1!
1%
#135470000000
0!
0%
#135475000000
1!
1%
#135480000000
0!
0%
#135485000000
1!
1%
#135490000000
0!
0%
#135495000000
1!
1%
#135500000000
0!
0%
#135505000000
1!
1%
#135510000000
0!
0%
#135515000000
1!
1%
#135520000000
0!
0%
#135525000000
1!
1%
#135530000000
0!
0%
#135535000000
1!
1%
#135540000000
0!
0%
#135545000000
1!
1%
#135550000000
0!
0%
#135555000000
1!
1%
#135560000000
0!
0%
#135565000000
1!
1%
#135570000000
0!
0%
#135575000000
1!
1%
#135580000000
0!
0%
#135585000000
1!
1%
#135590000000
0!
0%
#135595000000
1!
1%
#135600000000
0!
0%
#135605000000
1!
1%
#135610000000
0!
0%
#135615000000
1!
1%
#135620000000
0!
0%
#135625000000
1!
1%
#135630000000
0!
0%
#135635000000
1!
1%
#135640000000
0!
0%
#135645000000
1!
1%
#135650000000
0!
0%
#135655000000
1!
1%
#135660000000
0!
0%
#135665000000
1!
1%
#135670000000
0!
0%
#135675000000
1!
1%
#135680000000
0!
0%
#135685000000
1!
1%
#135690000000
0!
0%
#135695000000
1!
1%
#135700000000
0!
0%
#135705000000
1!
1%
#135710000000
0!
0%
#135715000000
1!
1%
#135720000000
0!
0%
#135725000000
1!
1%
#135730000000
0!
0%
#135735000000
1!
1%
#135740000000
0!
0%
#135745000000
1!
1%
#135750000000
0!
0%
#135755000000
1!
1%
#135760000000
0!
0%
#135765000000
1!
1%
#135770000000
0!
0%
#135775000000
1!
1%
#135780000000
0!
0%
#135785000000
1!
1%
#135790000000
0!
0%
#135795000000
1!
1%
#135800000000
0!
0%
#135805000000
1!
1%
#135810000000
0!
0%
#135815000000
1!
1%
#135820000000
0!
0%
#135825000000
1!
1%
#135830000000
0!
0%
#135835000000
1!
1%
#135840000000
0!
0%
#135845000000
1!
1%
#135850000000
0!
0%
#135855000000
1!
1%
#135860000000
0!
0%
#135865000000
1!
1%
#135870000000
0!
0%
#135875000000
1!
1%
#135880000000
0!
0%
#135885000000
1!
1%
#135890000000
0!
0%
#135895000000
1!
1%
#135900000000
0!
0%
#135905000000
1!
1%
#135910000000
0!
0%
#135915000000
1!
1%
#135920000000
0!
0%
#135925000000
1!
1%
#135930000000
0!
0%
#135935000000
1!
1%
#135940000000
0!
0%
#135945000000
1!
1%
#135950000000
0!
0%
#135955000000
1!
1%
#135960000000
0!
0%
#135965000000
1!
1%
#135970000000
0!
0%
#135975000000
1!
1%
#135980000000
0!
0%
#135985000000
1!
1%
#135990000000
0!
0%
#135995000000
1!
1%
#136000000000
0!
0%
#136005000000
1!
1%
#136010000000
0!
0%
#136015000000
1!
1%
#136020000000
0!
0%
#136025000000
1!
1%
#136030000000
0!
0%
#136035000000
1!
1%
#136040000000
0!
0%
#136045000000
1!
1%
#136050000000
0!
0%
#136055000000
1!
1%
#136060000000
0!
0%
#136065000000
1!
1%
#136070000000
0!
0%
#136075000000
1!
1%
#136080000000
0!
0%
#136085000000
1!
1%
#136090000000
0!
0%
#136095000000
1!
1%
#136100000000
0!
0%
#136105000000
1!
1%
#136110000000
0!
0%
#136115000000
1!
1%
#136120000000
0!
0%
#136125000000
1!
1%
#136130000000
0!
0%
#136135000000
1!
1%
#136140000000
0!
0%
#136145000000
1!
1%
#136150000000
0!
0%
#136155000000
1!
1%
#136160000000
0!
0%
#136165000000
1!
1%
#136170000000
0!
0%
#136175000000
1!
1%
#136180000000
0!
0%
#136185000000
1!
1%
#136190000000
0!
0%
#136195000000
1!
1%
#136200000000
0!
0%
#136205000000
1!
1%
#136210000000
0!
0%
#136215000000
1!
1%
#136220000000
0!
0%
#136225000000
1!
1%
#136230000000
0!
0%
#136235000000
1!
1%
#136240000000
0!
0%
#136245000000
1!
1%
#136250000000
0!
0%
#136255000000
1!
1%
#136260000000
0!
0%
#136265000000
1!
1%
#136270000000
0!
0%
#136275000000
1!
1%
#136280000000
0!
0%
#136285000000
1!
1%
#136290000000
0!
0%
#136295000000
1!
1%
#136300000000
0!
0%
#136305000000
1!
1%
#136310000000
0!
0%
#136315000000
1!
1%
#136320000000
0!
0%
#136325000000
1!
1%
#136330000000
0!
0%
#136335000000
1!
1%
#136340000000
0!
0%
#136345000000
1!
1%
#136350000000
0!
0%
#136355000000
1!
1%
#136360000000
0!
0%
#136365000000
1!
1%
#136370000000
0!
0%
#136375000000
1!
1%
#136380000000
0!
0%
#136385000000
1!
1%
#136390000000
0!
0%
#136395000000
1!
1%
#136400000000
0!
0%
#136405000000
1!
1%
#136410000000
0!
0%
#136415000000
1!
1%
#136420000000
0!
0%
#136425000000
1!
1%
#136430000000
0!
0%
#136435000000
1!
1%
#136440000000
0!
0%
#136445000000
1!
1%
#136450000000
0!
0%
#136455000000
1!
1%
#136460000000
0!
0%
#136465000000
1!
1%
#136470000000
0!
0%
#136475000000
1!
1%
#136480000000
0!
0%
#136485000000
1!
1%
#136490000000
0!
0%
#136495000000
1!
1%
#136500000000
0!
0%
#136505000000
1!
1%
#136510000000
0!
0%
#136515000000
1!
1%
#136520000000
0!
0%
#136525000000
1!
1%
#136530000000
0!
0%
#136535000000
1!
1%
#136540000000
0!
0%
#136545000000
1!
1%
#136550000000
0!
0%
#136555000000
1!
1%
#136560000000
0!
0%
#136565000000
1!
1%
#136570000000
0!
0%
#136575000000
1!
1%
#136580000000
0!
0%
#136585000000
1!
1%
#136590000000
0!
0%
#136595000000
1!
1%
#136600000000
0!
0%
#136605000000
1!
1%
#136610000000
0!
0%
#136615000000
1!
1%
#136620000000
0!
0%
#136625000000
1!
1%
#136630000000
0!
0%
#136635000000
1!
1%
#136640000000
0!
0%
#136645000000
1!
1%
#136650000000
0!
0%
#136655000000
1!
1%
#136660000000
0!
0%
#136665000000
1!
1%
#136670000000
0!
0%
#136675000000
1!
1%
#136680000000
0!
0%
#136685000000
1!
1%
#136690000000
0!
0%
#136695000000
1!
1%
#136700000000
0!
0%
#136705000000
1!
1%
#136710000000
0!
0%
#136715000000
1!
1%
#136720000000
0!
0%
#136725000000
1!
1%
#136730000000
0!
0%
#136735000000
1!
1%
#136740000000
0!
0%
#136745000000
1!
1%
#136750000000
0!
0%
#136755000000
1!
1%
#136760000000
0!
0%
#136765000000
1!
1%
#136770000000
0!
0%
#136775000000
1!
1%
#136780000000
0!
0%
#136785000000
1!
1%
#136790000000
0!
0%
#136795000000
1!
1%
#136800000000
0!
0%
#136805000000
1!
1%
#136810000000
0!
0%
#136815000000
1!
1%
#136820000000
0!
0%
#136825000000
1!
1%
#136830000000
0!
0%
#136835000000
1!
1%
#136840000000
0!
0%
#136845000000
1!
1%
#136850000000
0!
0%
#136855000000
1!
1%
#136860000000
0!
0%
#136865000000
1!
1%
#136870000000
0!
0%
#136875000000
1!
1%
#136880000000
0!
0%
#136885000000
1!
1%
#136890000000
0!
0%
#136895000000
1!
1%
#136900000000
0!
0%
#136905000000
1!
1%
#136910000000
0!
0%
#136915000000
1!
1%
#136920000000
0!
0%
#136925000000
1!
1%
#136930000000
0!
0%
#136935000000
1!
1%
#136940000000
0!
0%
#136945000000
1!
1%
#136950000000
0!
0%
#136955000000
1!
1%
#136960000000
0!
0%
#136965000000
1!
1%
#136970000000
0!
0%
#136975000000
1!
1%
#136980000000
0!
0%
#136985000000
1!
1%
#136990000000
0!
0%
#136995000000
1!
1%
#137000000000
0!
0%
#137005000000
1!
1%
#137010000000
0!
0%
#137015000000
1!
1%
#137020000000
0!
0%
#137025000000
1!
1%
#137030000000
0!
0%
#137035000000
1!
1%
#137040000000
0!
0%
#137045000000
1!
1%
#137050000000
0!
0%
#137055000000
1!
1%
#137060000000
0!
0%
#137065000000
1!
1%
#137070000000
0!
0%
#137075000000
1!
1%
#137080000000
0!
0%
#137085000000
1!
1%
#137090000000
0!
0%
#137095000000
1!
1%
#137100000000
0!
0%
#137105000000
1!
1%
#137110000000
0!
0%
#137115000000
1!
1%
#137120000000
0!
0%
#137125000000
1!
1%
#137130000000
0!
0%
#137135000000
1!
1%
#137140000000
0!
0%
#137145000000
1!
1%
#137150000000
0!
0%
#137155000000
1!
1%
#137160000000
0!
0%
#137165000000
1!
1%
#137170000000
0!
0%
#137175000000
1!
1%
#137180000000
0!
0%
#137185000000
1!
1%
#137190000000
0!
0%
#137195000000
1!
1%
#137200000000
0!
0%
#137205000000
1!
1%
#137210000000
0!
0%
#137215000000
1!
1%
#137220000000
0!
0%
#137225000000
1!
1%
#137230000000
0!
0%
#137235000000
1!
1%
#137240000000
0!
0%
#137245000000
1!
1%
#137250000000
0!
0%
#137255000000
1!
1%
#137260000000
0!
0%
#137265000000
1!
1%
#137270000000
0!
0%
#137275000000
1!
1%
#137280000000
0!
0%
#137285000000
1!
1%
#137290000000
0!
0%
#137295000000
1!
1%
#137300000000
0!
0%
#137305000000
1!
1%
#137310000000
0!
0%
#137315000000
1!
1%
#137320000000
0!
0%
#137325000000
1!
1%
#137330000000
0!
0%
#137335000000
1!
1%
#137340000000
0!
0%
#137345000000
1!
1%
#137350000000
0!
0%
#137355000000
1!
1%
#137360000000
0!
0%
#137365000000
1!
1%
#137370000000
0!
0%
#137375000000
1!
1%
#137380000000
0!
0%
#137385000000
1!
1%
#137390000000
0!
0%
#137395000000
1!
1%
#137400000000
0!
0%
#137405000000
1!
1%
#137410000000
0!
0%
#137415000000
1!
1%
#137420000000
0!
0%
#137425000000
1!
1%
#137430000000
0!
0%
#137435000000
1!
1%
#137440000000
0!
0%
#137445000000
1!
1%
#137450000000
0!
0%
#137455000000
1!
1%
#137460000000
0!
0%
#137465000000
1!
1%
#137470000000
0!
0%
#137475000000
1!
1%
#137480000000
0!
0%
#137485000000
1!
1%
#137490000000
0!
0%
#137495000000
1!
1%
#137500000000
0!
0%
#137505000000
1!
1%
#137510000000
0!
0%
#137515000000
1!
1%
#137520000000
0!
0%
#137525000000
1!
1%
#137530000000
0!
0%
#137535000000
1!
1%
#137540000000
0!
0%
#137545000000
1!
1%
#137550000000
0!
0%
#137555000000
1!
1%
#137560000000
0!
0%
#137565000000
1!
1%
#137570000000
0!
0%
#137575000000
1!
1%
#137580000000
0!
0%
#137585000000
1!
1%
#137590000000
0!
0%
#137595000000
1!
1%
#137600000000
0!
0%
#137605000000
1!
1%
#137610000000
0!
0%
#137615000000
1!
1%
#137620000000
0!
0%
#137625000000
1!
1%
#137630000000
0!
0%
#137635000000
1!
1%
#137640000000
0!
0%
#137645000000
1!
1%
#137650000000
0!
0%
#137655000000
1!
1%
#137660000000
0!
0%
#137665000000
1!
1%
#137670000000
0!
0%
#137675000000
1!
1%
#137680000000
0!
0%
#137685000000
1!
1%
#137690000000
0!
0%
#137695000000
1!
1%
#137700000000
0!
0%
#137705000000
1!
1%
#137710000000
0!
0%
#137715000000
1!
1%
#137720000000
0!
0%
#137725000000
1!
1%
#137730000000
0!
0%
#137735000000
1!
1%
#137740000000
0!
0%
#137745000000
1!
1%
#137750000000
0!
0%
#137755000000
1!
1%
#137760000000
0!
0%
#137765000000
1!
1%
#137770000000
0!
0%
#137775000000
1!
1%
#137780000000
0!
0%
#137785000000
1!
1%
#137790000000
0!
0%
#137795000000
1!
1%
#137800000000
0!
0%
#137805000000
1!
1%
#137810000000
0!
0%
#137815000000
1!
1%
#137820000000
0!
0%
#137825000000
1!
1%
#137830000000
0!
0%
#137835000000
1!
1%
#137840000000
0!
0%
#137845000000
1!
1%
#137850000000
0!
0%
#137855000000
1!
1%
#137860000000
0!
0%
#137865000000
1!
1%
#137870000000
0!
0%
#137875000000
1!
1%
#137880000000
0!
0%
#137885000000
1!
1%
#137890000000
0!
0%
#137895000000
1!
1%
#137900000000
0!
0%
#137905000000
1!
1%
#137910000000
0!
0%
#137915000000
1!
1%
#137920000000
0!
0%
#137925000000
1!
1%
#137930000000
0!
0%
#137935000000
1!
1%
#137940000000
0!
0%
#137945000000
1!
1%
#137950000000
0!
0%
#137955000000
1!
1%
#137960000000
0!
0%
#137965000000
1!
1%
#137970000000
0!
0%
#137975000000
1!
1%
#137980000000
0!
0%
#137985000000
1!
1%
#137990000000
0!
0%
#137995000000
1!
1%
#138000000000
0!
0%
#138005000000
1!
1%
#138010000000
0!
0%
#138015000000
1!
1%
#138020000000
0!
0%
#138025000000
1!
1%
#138030000000
0!
0%
#138035000000
1!
1%
#138040000000
0!
0%
#138045000000
1!
1%
#138050000000
0!
0%
#138055000000
1!
1%
#138060000000
0!
0%
#138065000000
1!
1%
#138070000000
0!
0%
#138075000000
1!
1%
#138080000000
0!
0%
#138085000000
1!
1%
#138090000000
0!
0%
#138095000000
1!
1%
#138100000000
0!
0%
#138105000000
1!
1%
#138110000000
0!
0%
#138115000000
1!
1%
#138120000000
0!
0%
#138125000000
1!
1%
#138130000000
0!
0%
#138135000000
1!
1%
#138140000000
0!
0%
#138145000000
1!
1%
#138150000000
0!
0%
#138155000000
1!
1%
#138160000000
0!
0%
#138165000000
1!
1%
#138170000000
0!
0%
#138175000000
1!
1%
#138180000000
0!
0%
#138185000000
1!
1%
#138190000000
0!
0%
#138195000000
1!
1%
#138200000000
0!
0%
#138205000000
1!
1%
#138210000000
0!
0%
#138215000000
1!
1%
#138220000000
0!
0%
#138225000000
1!
1%
#138230000000
0!
0%
#138235000000
1!
1%
#138240000000
0!
0%
#138245000000
1!
1%
#138250000000
0!
0%
#138255000000
1!
1%
#138260000000
0!
0%
#138265000000
1!
1%
#138270000000
0!
0%
#138275000000
1!
1%
#138280000000
0!
0%
#138285000000
1!
1%
#138290000000
0!
0%
#138295000000
1!
1%
#138300000000
0!
0%
#138305000000
1!
1%
#138310000000
0!
0%
#138315000000
1!
1%
#138320000000
0!
0%
#138325000000
1!
1%
#138330000000
0!
0%
#138335000000
1!
1%
#138340000000
0!
0%
#138345000000
1!
1%
#138350000000
0!
0%
#138355000000
1!
1%
#138360000000
0!
0%
#138365000000
1!
1%
#138370000000
0!
0%
#138375000000
1!
1%
#138380000000
0!
0%
#138385000000
1!
1%
#138390000000
0!
0%
#138395000000
1!
1%
#138400000000
0!
0%
#138405000000
1!
1%
#138410000000
0!
0%
#138415000000
1!
1%
#138420000000
0!
0%
#138425000000
1!
1%
#138430000000
0!
0%
#138435000000
1!
1%
#138440000000
0!
0%
#138445000000
1!
1%
#138450000000
0!
0%
#138455000000
1!
1%
#138460000000
0!
0%
#138465000000
1!
1%
#138470000000
0!
0%
#138475000000
1!
1%
#138480000000
0!
0%
#138485000000
1!
1%
#138490000000
0!
0%
#138495000000
1!
1%
#138500000000
0!
0%
#138505000000
1!
1%
#138510000000
0!
0%
#138515000000
1!
1%
#138520000000
0!
0%
#138525000000
1!
1%
#138530000000
0!
0%
#138535000000
1!
1%
#138540000000
0!
0%
#138545000000
1!
1%
#138550000000
0!
0%
#138555000000
1!
1%
#138560000000
0!
0%
#138565000000
1!
1%
#138570000000
0!
0%
#138575000000
1!
1%
#138580000000
0!
0%
#138585000000
1!
1%
#138590000000
0!
0%
#138595000000
1!
1%
#138600000000
0!
0%
#138605000000
1!
1%
#138610000000
0!
0%
#138615000000
1!
1%
#138620000000
0!
0%
#138625000000
1!
1%
#138630000000
0!
0%
#138635000000
1!
1%
#138640000000
0!
0%
#138645000000
1!
1%
#138650000000
0!
0%
#138655000000
1!
1%
#138660000000
0!
0%
#138665000000
1!
1%
#138670000000
0!
0%
#138675000000
1!
1%
#138680000000
0!
0%
#138685000000
1!
1%
#138690000000
0!
0%
#138695000000
1!
1%
#138700000000
0!
0%
#138705000000
1!
1%
#138710000000
0!
0%
#138715000000
1!
1%
#138720000000
0!
0%
#138725000000
1!
1%
#138730000000
0!
0%
#138735000000
1!
1%
#138740000000
0!
0%
#138745000000
1!
1%
#138750000000
0!
0%
#138755000000
1!
1%
#138760000000
0!
0%
#138765000000
1!
1%
#138770000000
0!
0%
#138775000000
1!
1%
#138780000000
0!
0%
#138785000000
1!
1%
#138790000000
0!
0%
#138795000000
1!
1%
#138800000000
0!
0%
#138805000000
1!
1%
#138810000000
0!
0%
#138815000000
1!
1%
#138820000000
0!
0%
#138825000000
1!
1%
#138830000000
0!
0%
#138835000000
1!
1%
#138840000000
0!
0%
#138845000000
1!
1%
#138850000000
0!
0%
#138855000000
1!
1%
#138860000000
0!
0%
#138865000000
1!
1%
#138870000000
0!
0%
#138875000000
1!
1%
#138880000000
0!
0%
#138885000000
1!
1%
#138890000000
0!
0%
#138895000000
1!
1%
#138900000000
0!
0%
#138905000000
1!
1%
#138910000000
0!
0%
#138915000000
1!
1%
#138920000000
0!
0%
#138925000000
1!
1%
#138930000000
0!
0%
#138935000000
1!
1%
#138940000000
0!
0%
#138945000000
1!
1%
#138950000000
0!
0%
#138955000000
1!
1%
#138960000000
0!
0%
#138965000000
1!
1%
#138970000000
0!
0%
#138975000000
1!
1%
#138980000000
0!
0%
#138985000000
1!
1%
#138990000000
0!
0%
#138995000000
1!
1%
#139000000000
0!
0%
#139005000000
1!
1%
#139010000000
0!
0%
#139015000000
1!
1%
#139020000000
0!
0%
#139025000000
1!
1%
#139030000000
0!
0%
#139035000000
1!
1%
#139040000000
0!
0%
#139045000000
1!
1%
#139050000000
0!
0%
#139055000000
1!
1%
#139060000000
0!
0%
#139065000000
1!
1%
#139070000000
0!
0%
#139075000000
1!
1%
#139080000000
0!
0%
#139085000000
1!
1%
#139090000000
0!
0%
#139095000000
1!
1%
#139100000000
0!
0%
#139105000000
1!
1%
#139110000000
0!
0%
#139115000000
1!
1%
#139120000000
0!
0%
#139125000000
1!
1%
#139130000000
0!
0%
#139135000000
1!
1%
#139140000000
0!
0%
#139145000000
1!
1%
#139150000000
0!
0%
#139155000000
1!
1%
#139160000000
0!
0%
#139165000000
1!
1%
#139170000000
0!
0%
#139175000000
1!
1%
#139180000000
0!
0%
#139185000000
1!
1%
#139190000000
0!
0%
#139195000000
1!
1%
#139200000000
0!
0%
#139205000000
1!
1%
#139210000000
0!
0%
#139215000000
1!
1%
#139220000000
0!
0%
#139225000000
1!
1%
#139230000000
0!
0%
#139235000000
1!
1%
#139240000000
0!
0%
#139245000000
1!
1%
#139250000000
0!
0%
#139255000000
1!
1%
#139260000000
0!
0%
#139265000000
1!
1%
#139270000000
0!
0%
#139275000000
1!
1%
#139280000000
0!
0%
#139285000000
1!
1%
#139290000000
0!
0%
#139295000000
1!
1%
#139300000000
0!
0%
#139305000000
1!
1%
#139310000000
0!
0%
#139315000000
1!
1%
#139320000000
0!
0%
#139325000000
1!
1%
#139330000000
0!
0%
#139335000000
1!
1%
#139340000000
0!
0%
#139345000000
1!
1%
#139350000000
0!
0%
#139355000000
1!
1%
#139360000000
0!
0%
#139365000000
1!
1%
#139370000000
0!
0%
#139375000000
1!
1%
#139380000000
0!
0%
#139385000000
1!
1%
#139390000000
0!
0%
#139395000000
1!
1%
#139400000000
0!
0%
#139405000000
1!
1%
#139410000000
0!
0%
#139415000000
1!
1%
#139420000000
0!
0%
#139425000000
1!
1%
#139430000000
0!
0%
#139435000000
1!
1%
#139440000000
0!
0%
#139445000000
1!
1%
#139450000000
0!
0%
#139455000000
1!
1%
#139460000000
0!
0%
#139465000000
1!
1%
#139470000000
0!
0%
#139475000000
1!
1%
#139480000000
0!
0%
#139485000000
1!
1%
#139490000000
0!
0%
#139495000000
1!
1%
#139500000000
0!
0%
#139505000000
1!
1%
#139510000000
0!
0%
#139515000000
1!
1%
#139520000000
0!
0%
#139525000000
1!
1%
#139530000000
0!
0%
#139535000000
1!
1%
#139540000000
0!
0%
#139545000000
1!
1%
#139550000000
0!
0%
#139555000000
1!
1%
#139560000000
0!
0%
#139565000000
1!
1%
#139570000000
0!
0%
#139575000000
1!
1%
#139580000000
0!
0%
#139585000000
1!
1%
#139590000000
0!
0%
#139595000000
1!
1%
#139600000000
0!
0%
#139605000000
1!
1%
#139610000000
0!
0%
#139615000000
1!
1%
#139620000000
0!
0%
#139625000000
1!
1%
#139630000000
0!
0%
#139635000000
1!
1%
#139640000000
0!
0%
#139645000000
1!
1%
#139650000000
0!
0%
#139655000000
1!
1%
#139660000000
0!
0%
#139665000000
1!
1%
#139670000000
0!
0%
#139675000000
1!
1%
#139680000000
0!
0%
#139685000000
1!
1%
#139690000000
0!
0%
#139695000000
1!
1%
#139700000000
0!
0%
#139705000000
1!
1%
#139710000000
0!
0%
#139715000000
1!
1%
#139720000000
0!
0%
#139725000000
1!
1%
#139730000000
0!
0%
#139735000000
1!
1%
#139740000000
0!
0%
#139745000000
1!
1%
#139750000000
0!
0%
#139755000000
1!
1%
#139760000000
0!
0%
#139765000000
1!
1%
#139770000000
0!
0%
#139775000000
1!
1%
#139780000000
0!
0%
#139785000000
1!
1%
#139790000000
0!
0%
#139795000000
1!
1%
#139800000000
0!
0%
#139805000000
1!
1%
#139810000000
0!
0%
#139815000000
1!
1%
#139820000000
0!
0%
#139825000000
1!
1%
#139830000000
0!
0%
#139835000000
1!
1%
#139840000000
0!
0%
#139845000000
1!
1%
#139850000000
0!
0%
#139855000000
1!
1%
#139860000000
0!
0%
#139865000000
1!
1%
#139870000000
0!
0%
#139875000000
1!
1%
#139880000000
0!
0%
#139885000000
1!
1%
#139890000000
0!
0%
#139895000000
1!
1%
#139900000000
0!
0%
#139905000000
1!
1%
#139910000000
0!
0%
#139915000000
1!
1%
#139920000000
0!
0%
#139925000000
1!
1%
#139930000000
0!
0%
#139935000000
1!
1%
#139940000000
0!
0%
#139945000000
1!
1%
#139950000000
0!
0%
#139955000000
1!
1%
#139960000000
0!
0%
#139965000000
1!
1%
#139970000000
0!
0%
#139975000000
1!
1%
#139980000000
0!
0%
#139985000000
1!
1%
#139990000000
0!
0%
#139995000000
1!
1%
#140000000000
0!
0%
#140005000000
1!
1%
#140010000000
0!
0%
#140015000000
1!
1%
#140020000000
0!
0%
#140025000000
1!
1%
#140030000000
0!
0%
#140035000000
1!
1%
#140040000000
0!
0%
#140045000000
1!
1%
#140050000000
0!
0%
#140055000000
1!
1%
#140060000000
0!
0%
#140065000000
1!
1%
#140070000000
0!
0%
#140075000000
1!
1%
#140080000000
0!
0%
#140085000000
1!
1%
#140090000000
0!
0%
#140095000000
1!
1%
#140100000000
0!
0%
#140105000000
1!
1%
#140110000000
0!
0%
#140115000000
1!
1%
#140120000000
0!
0%
#140125000000
1!
1%
#140130000000
0!
0%
#140135000000
1!
1%
#140140000000
0!
0%
#140145000000
1!
1%
#140150000000
0!
0%
#140155000000
1!
1%
#140160000000
0!
0%
#140165000000
1!
1%
#140170000000
0!
0%
#140175000000
1!
1%
#140180000000
0!
0%
#140185000000
1!
1%
#140190000000
0!
0%
#140195000000
1!
1%
#140200000000
0!
0%
#140205000000
1!
1%
#140210000000
0!
0%
#140215000000
1!
1%
#140220000000
0!
0%
#140225000000
1!
1%
#140230000000
0!
0%
#140235000000
1!
1%
#140240000000
0!
0%
#140245000000
1!
1%
#140250000000
0!
0%
#140255000000
1!
1%
#140260000000
0!
0%
#140265000000
1!
1%
#140270000000
0!
0%
#140275000000
1!
1%
#140280000000
0!
0%
#140285000000
1!
1%
#140290000000
0!
0%
#140295000000
1!
1%
#140300000000
0!
0%
#140305000000
1!
1%
#140310000000
0!
0%
#140315000000
1!
1%
#140320000000
0!
0%
#140325000000
1!
1%
#140330000000
0!
0%
#140335000000
1!
1%
#140340000000
0!
0%
#140345000000
1!
1%
#140350000000
0!
0%
#140355000000
1!
1%
#140360000000
0!
0%
#140365000000
1!
1%
#140370000000
0!
0%
#140375000000
1!
1%
#140380000000
0!
0%
#140385000000
1!
1%
#140390000000
0!
0%
#140395000000
1!
1%
#140400000000
0!
0%
#140405000000
1!
1%
#140410000000
0!
0%
#140415000000
1!
1%
#140420000000
0!
0%
#140425000000
1!
1%
#140430000000
0!
0%
#140435000000
1!
1%
#140440000000
0!
0%
#140445000000
1!
1%
#140450000000
0!
0%
#140455000000
1!
1%
#140460000000
0!
0%
#140465000000
1!
1%
#140470000000
0!
0%
#140475000000
1!
1%
#140480000000
0!
0%
#140485000000
1!
1%
#140490000000
0!
0%
#140495000000
1!
1%
#140500000000
0!
0%
#140505000000
1!
1%
#140510000000
0!
0%
#140515000000
1!
1%
#140520000000
0!
0%
#140525000000
1!
1%
#140530000000
0!
0%
#140535000000
1!
1%
#140540000000
0!
0%
#140545000000
1!
1%
#140550000000
0!
0%
#140555000000
1!
1%
#140560000000
0!
0%
#140565000000
1!
1%
#140570000000
0!
0%
#140575000000
1!
1%
#140580000000
0!
0%
#140585000000
1!
1%
#140590000000
0!
0%
#140595000000
1!
1%
#140600000000
0!
0%
#140605000000
1!
1%
#140610000000
0!
0%
#140615000000
1!
1%
#140620000000
0!
0%
#140625000000
1!
1%
#140630000000
0!
0%
#140635000000
1!
1%
#140640000000
0!
0%
#140645000000
1!
1%
#140650000000
0!
0%
#140655000000
1!
1%
#140660000000
0!
0%
#140665000000
1!
1%
#140670000000
0!
0%
#140675000000
1!
1%
#140680000000
0!
0%
#140685000000
1!
1%
#140690000000
0!
0%
#140695000000
1!
1%
#140700000000
0!
0%
#140705000000
1!
1%
#140710000000
0!
0%
#140715000000
1!
1%
#140720000000
0!
0%
#140725000000
1!
1%
#140730000000
0!
0%
#140735000000
1!
1%
#140740000000
0!
0%
#140745000000
1!
1%
#140750000000
0!
0%
#140755000000
1!
1%
#140760000000
0!
0%
#140765000000
1!
1%
#140770000000
0!
0%
#140775000000
1!
1%
#140780000000
0!
0%
#140785000000
1!
1%
#140790000000
0!
0%
#140795000000
1!
1%
#140800000000
0!
0%
#140805000000
1!
1%
#140810000000
0!
0%
#140815000000
1!
1%
#140820000000
0!
0%
#140825000000
1!
1%
#140830000000
0!
0%
#140835000000
1!
1%
#140840000000
0!
0%
#140845000000
1!
1%
#140850000000
0!
0%
#140855000000
1!
1%
#140860000000
0!
0%
#140865000000
1!
1%
#140870000000
0!
0%
#140875000000
1!
1%
#140880000000
0!
0%
#140885000000
1!
1%
#140890000000
0!
0%
#140895000000
1!
1%
#140900000000
0!
0%
#140905000000
1!
1%
#140910000000
0!
0%
#140915000000
1!
1%
#140920000000
0!
0%
#140925000000
1!
1%
#140930000000
0!
0%
#140935000000
1!
1%
#140940000000
0!
0%
#140945000000
1!
1%
#140950000000
0!
0%
#140955000000
1!
1%
#140960000000
0!
0%
#140965000000
1!
1%
#140970000000
0!
0%
#140975000000
1!
1%
#140980000000
0!
0%
#140985000000
1!
1%
#140990000000
0!
0%
#140995000000
1!
1%
#141000000000
0!
0%
#141005000000
1!
1%
#141010000000
0!
0%
#141015000000
1!
1%
#141020000000
0!
0%
#141025000000
1!
1%
#141030000000
0!
0%
#141035000000
1!
1%
#141040000000
0!
0%
#141045000000
1!
1%
#141050000000
0!
0%
#141055000000
1!
1%
#141060000000
0!
0%
#141065000000
1!
1%
#141070000000
0!
0%
#141075000000
1!
1%
#141080000000
0!
0%
#141085000000
1!
1%
#141090000000
0!
0%
#141095000000
1!
1%
#141100000000
0!
0%
#141105000000
1!
1%
#141110000000
0!
0%
#141115000000
1!
1%
#141120000000
0!
0%
#141125000000
1!
1%
#141130000000
0!
0%
#141135000000
1!
1%
#141140000000
0!
0%
#141145000000
1!
1%
#141150000000
0!
0%
#141155000000
1!
1%
#141160000000
0!
0%
#141165000000
1!
1%
#141170000000
0!
0%
#141175000000
1!
1%
#141180000000
0!
0%
#141185000000
1!
1%
#141190000000
0!
0%
#141195000000
1!
1%
#141200000000
0!
0%
#141205000000
1!
1%
#141210000000
0!
0%
#141215000000
1!
1%
#141220000000
0!
0%
#141225000000
1!
1%
#141230000000
0!
0%
#141235000000
1!
1%
#141240000000
0!
0%
#141245000000
1!
1%
#141250000000
0!
0%
#141255000000
1!
1%
#141260000000
0!
0%
#141265000000
1!
1%
#141270000000
0!
0%
#141275000000
1!
1%
#141280000000
0!
0%
#141285000000
1!
1%
#141290000000
0!
0%
#141295000000
1!
1%
#141300000000
0!
0%
#141305000000
1!
1%
#141310000000
0!
0%
#141315000000
1!
1%
#141320000000
0!
0%
#141325000000
1!
1%
#141330000000
0!
0%
#141335000000
1!
1%
#141340000000
0!
0%
#141345000000
1!
1%
#141350000000
0!
0%
#141355000000
1!
1%
#141360000000
0!
0%
#141365000000
1!
1%
#141370000000
0!
0%
#141375000000
1!
1%
#141380000000
0!
0%
#141385000000
1!
1%
#141390000000
0!
0%
#141395000000
1!
1%
#141400000000
0!
0%
#141405000000
1!
1%
#141410000000
0!
0%
#141415000000
1!
1%
#141420000000
0!
0%
#141425000000
1!
1%
#141430000000
0!
0%
#141435000000
1!
1%
#141440000000
0!
0%
#141445000000
1!
1%
#141450000000
0!
0%
#141455000000
1!
1%
#141460000000
0!
0%
#141465000000
1!
1%
#141470000000
0!
0%
#141475000000
1!
1%
#141480000000
0!
0%
#141485000000
1!
1%
#141490000000
0!
0%
#141495000000
1!
1%
#141500000000
0!
0%
#141505000000
1!
1%
#141510000000
0!
0%
#141515000000
1!
1%
#141520000000
0!
0%
#141525000000
1!
1%
#141530000000
0!
0%
#141535000000
1!
1%
#141540000000
0!
0%
#141545000000
1!
1%
#141550000000
0!
0%
#141555000000
1!
1%
#141560000000
0!
0%
#141565000000
1!
1%
#141570000000
0!
0%
#141575000000
1!
1%
#141580000000
0!
0%
#141585000000
1!
1%
#141590000000
0!
0%
#141595000000
1!
1%
#141600000000
0!
0%
#141605000000
1!
1%
#141610000000
0!
0%
#141615000000
1!
1%
#141620000000
0!
0%
#141625000000
1!
1%
#141630000000
0!
0%
#141635000000
1!
1%
#141640000000
0!
0%
#141645000000
1!
1%
#141650000000
0!
0%
#141655000000
1!
1%
#141660000000
0!
0%
#141665000000
1!
1%
#141670000000
0!
0%
#141675000000
1!
1%
#141680000000
0!
0%
#141685000000
1!
1%
#141690000000
0!
0%
#141695000000
1!
1%
#141700000000
0!
0%
#141705000000
1!
1%
#141710000000
0!
0%
#141715000000
1!
1%
#141720000000
0!
0%
#141725000000
1!
1%
#141730000000
0!
0%
#141735000000
1!
1%
#141740000000
0!
0%
#141745000000
1!
1%
#141750000000
0!
0%
#141755000000
1!
1%
#141760000000
0!
0%
#141765000000
1!
1%
#141770000000
0!
0%
#141775000000
1!
1%
#141780000000
0!
0%
#141785000000
1!
1%
#141790000000
0!
0%
#141795000000
1!
1%
#141800000000
0!
0%
#141805000000
1!
1%
#141810000000
0!
0%
#141815000000
1!
1%
#141820000000
0!
0%
#141825000000
1!
1%
#141830000000
0!
0%
#141835000000
1!
1%
#141840000000
0!
0%
#141845000000
1!
1%
#141850000000
0!
0%
#141855000000
1!
1%
#141860000000
0!
0%
#141865000000
1!
1%
#141870000000
0!
0%
#141875000000
1!
1%
#141880000000
0!
0%
#141885000000
1!
1%
#141890000000
0!
0%
#141895000000
1!
1%
#141900000000
0!
0%
#141905000000
1!
1%
#141910000000
0!
0%
#141915000000
1!
1%
#141920000000
0!
0%
#141925000000
1!
1%
#141930000000
0!
0%
#141935000000
1!
1%
#141940000000
0!
0%
#141945000000
1!
1%
#141950000000
0!
0%
#141955000000
1!
1%
#141960000000
0!
0%
#141965000000
1!
1%
#141970000000
0!
0%
#141975000000
1!
1%
#141980000000
0!
0%
#141985000000
1!
1%
#141990000000
0!
0%
#141995000000
1!
1%
#142000000000
0!
0%
#142005000000
1!
1%
#142010000000
0!
0%
#142015000000
1!
1%
#142020000000
0!
0%
#142025000000
1!
1%
#142030000000
0!
0%
#142035000000
1!
1%
#142040000000
0!
0%
#142045000000
1!
1%
#142050000000
0!
0%
#142055000000
1!
1%
#142060000000
0!
0%
#142065000000
1!
1%
#142070000000
0!
0%
#142075000000
1!
1%
#142080000000
0!
0%
#142085000000
1!
1%
#142090000000
0!
0%
#142095000000
1!
1%
#142100000000
0!
0%
#142105000000
1!
1%
#142110000000
0!
0%
#142115000000
1!
1%
#142120000000
0!
0%
#142125000000
1!
1%
#142130000000
0!
0%
#142135000000
1!
1%
#142140000000
0!
0%
#142145000000
1!
1%
#142150000000
0!
0%
#142155000000
1!
1%
#142160000000
0!
0%
#142165000000
1!
1%
#142170000000
0!
0%
#142175000000
1!
1%
#142180000000
0!
0%
#142185000000
1!
1%
#142190000000
0!
0%
#142195000000
1!
1%
#142200000000
0!
0%
#142205000000
1!
1%
#142210000000
0!
0%
#142215000000
1!
1%
#142220000000
0!
0%
#142225000000
1!
1%
#142230000000
0!
0%
#142235000000
1!
1%
#142240000000
0!
0%
#142245000000
1!
1%
#142250000000
0!
0%
#142255000000
1!
1%
#142260000000
0!
0%
#142265000000
1!
1%
#142270000000
0!
0%
#142275000000
1!
1%
#142280000000
0!
0%
#142285000000
1!
1%
#142290000000
0!
0%
#142295000000
1!
1%
#142300000000
0!
0%
#142305000000
1!
1%
#142310000000
0!
0%
#142315000000
1!
1%
#142320000000
0!
0%
#142325000000
1!
1%
#142330000000
0!
0%
#142335000000
1!
1%
#142340000000
0!
0%
#142345000000
1!
1%
#142350000000
0!
0%
#142355000000
1!
1%
#142360000000
0!
0%
#142365000000
1!
1%
#142370000000
0!
0%
#142375000000
1!
1%
#142380000000
0!
0%
#142385000000
1!
1%
#142390000000
0!
0%
#142395000000
1!
1%
#142400000000
0!
0%
#142405000000
1!
1%
#142410000000
0!
0%
#142415000000
1!
1%
#142420000000
0!
0%
#142425000000
1!
1%
#142430000000
0!
0%
#142435000000
1!
1%
#142440000000
0!
0%
#142445000000
1!
1%
#142450000000
0!
0%
#142455000000
1!
1%
#142460000000
0!
0%
#142465000000
1!
1%
#142470000000
0!
0%
#142475000000
1!
1%
#142480000000
0!
0%
#142485000000
1!
1%
#142490000000
0!
0%
#142495000000
1!
1%
#142500000000
0!
0%
#142505000000
1!
1%
#142510000000
0!
0%
#142515000000
1!
1%
#142520000000
0!
0%
#142525000000
1!
1%
#142530000000
0!
0%
#142535000000
1!
1%
#142540000000
0!
0%
#142545000000
1!
1%
#142550000000
0!
0%
#142555000000
1!
1%
#142560000000
0!
0%
#142565000000
1!
1%
#142570000000
0!
0%
#142575000000
1!
1%
#142580000000
0!
0%
#142585000000
1!
1%
#142590000000
0!
0%
#142595000000
1!
1%
#142600000000
0!
0%
#142605000000
1!
1%
#142610000000
0!
0%
#142615000000
1!
1%
#142620000000
0!
0%
#142625000000
1!
1%
#142630000000
0!
0%
#142635000000
1!
1%
#142640000000
0!
0%
#142645000000
1!
1%
#142650000000
0!
0%
#142655000000
1!
1%
#142660000000
0!
0%
#142665000000
1!
1%
#142670000000
0!
0%
#142675000000
1!
1%
#142680000000
0!
0%
#142685000000
1!
1%
#142690000000
0!
0%
#142695000000
1!
1%
#142700000000
0!
0%
#142705000000
1!
1%
#142710000000
0!
0%
#142715000000
1!
1%
#142720000000
0!
0%
#142725000000
1!
1%
#142730000000
0!
0%
#142735000000
1!
1%
#142740000000
0!
0%
#142745000000
1!
1%
#142750000000
0!
0%
#142755000000
1!
1%
#142760000000
0!
0%
#142765000000
1!
1%
#142770000000
0!
0%
#142775000000
1!
1%
#142780000000
0!
0%
#142785000000
1!
1%
#142790000000
0!
0%
#142795000000
1!
1%
#142800000000
0!
0%
#142805000000
1!
1%
#142810000000
0!
0%
#142815000000
1!
1%
#142820000000
0!
0%
#142825000000
1!
1%
#142830000000
0!
0%
#142835000000
1!
1%
#142840000000
0!
0%
#142845000000
1!
1%
#142850000000
0!
0%
#142855000000
1!
1%
#142860000000
0!
0%
#142865000000
1!
1%
#142870000000
0!
0%
#142875000000
1!
1%
#142880000000
0!
0%
#142885000000
1!
1%
#142890000000
0!
0%
#142895000000
1!
1%
#142900000000
0!
0%
#142905000000
1!
1%
#142910000000
0!
0%
#142915000000
1!
1%
#142920000000
0!
0%
#142925000000
1!
1%
#142930000000
0!
0%
#142935000000
1!
1%
#142940000000
0!
0%
#142945000000
1!
1%
#142950000000
0!
0%
#142955000000
1!
1%
#142960000000
0!
0%
#142965000000
1!
1%
#142970000000
0!
0%
#142975000000
1!
1%
#142980000000
0!
0%
#142985000000
1!
1%
#142990000000
0!
0%
#142995000000
1!
1%
#143000000000
0!
0%
#143005000000
1!
1%
#143010000000
0!
0%
#143015000000
1!
1%
#143020000000
0!
0%
#143025000000
1!
1%
#143030000000
0!
0%
#143035000000
1!
1%
#143040000000
0!
0%
#143045000000
1!
1%
#143050000000
0!
0%
#143055000000
1!
1%
#143060000000
0!
0%
#143065000000
1!
1%
#143070000000
0!
0%
#143075000000
1!
1%
#143080000000
0!
0%
#143085000000
1!
1%
#143090000000
0!
0%
#143095000000
1!
1%
#143100000000
0!
0%
#143105000000
1!
1%
#143110000000
0!
0%
#143115000000
1!
1%
#143120000000
0!
0%
#143125000000
1!
1%
#143130000000
0!
0%
#143135000000
1!
1%
#143140000000
0!
0%
#143145000000
1!
1%
#143150000000
0!
0%
#143155000000
1!
1%
#143160000000
0!
0%
#143165000000
1!
1%
#143170000000
0!
0%
#143175000000
1!
1%
#143180000000
0!
0%
#143185000000
1!
1%
#143190000000
0!
0%
#143195000000
1!
1%
#143200000000
0!
0%
#143205000000
1!
1%
#143210000000
0!
0%
#143215000000
1!
1%
#143220000000
0!
0%
#143225000000
1!
1%
#143230000000
0!
0%
#143235000000
1!
1%
#143240000000
0!
0%
#143245000000
1!
1%
#143250000000
0!
0%
#143255000000
1!
1%
#143260000000
0!
0%
#143265000000
1!
1%
#143270000000
0!
0%
#143275000000
1!
1%
#143280000000
0!
0%
#143285000000
1!
1%
#143290000000
0!
0%
#143295000000
1!
1%
#143300000000
0!
0%
#143305000000
1!
1%
#143310000000
0!
0%
#143315000000
1!
1%
#143320000000
0!
0%
#143325000000
1!
1%
#143330000000
0!
0%
#143335000000
1!
1%
#143340000000
0!
0%
#143345000000
1!
1%
#143350000000
0!
0%
#143355000000
1!
1%
#143360000000
0!
0%
#143365000000
1!
1%
#143370000000
0!
0%
#143375000000
1!
1%
#143380000000
0!
0%
#143385000000
1!
1%
#143390000000
0!
0%
#143395000000
1!
1%
#143400000000
0!
0%
#143405000000
1!
1%
#143410000000
0!
0%
#143415000000
1!
1%
#143420000000
0!
0%
#143425000000
1!
1%
#143430000000
0!
0%
#143435000000
1!
1%
#143440000000
0!
0%
#143445000000
1!
1%
#143450000000
0!
0%
#143455000000
1!
1%
#143460000000
0!
0%
#143465000000
1!
1%
#143470000000
0!
0%
#143475000000
1!
1%
#143480000000
0!
0%
#143485000000
1!
1%
#143490000000
0!
0%
#143495000000
1!
1%
#143500000000
0!
0%
#143505000000
1!
1%
#143510000000
0!
0%
#143515000000
1!
1%
#143520000000
0!
0%
#143525000000
1!
1%
#143530000000
0!
0%
#143535000000
1!
1%
#143540000000
0!
0%
#143545000000
1!
1%
#143550000000
0!
0%
#143555000000
1!
1%
#143560000000
0!
0%
#143565000000
1!
1%
#143570000000
0!
0%
#143575000000
1!
1%
#143580000000
0!
0%
#143585000000
1!
1%
#143590000000
0!
0%
#143595000000
1!
1%
#143600000000
0!
0%
#143605000000
1!
1%
#143610000000
0!
0%
#143615000000
1!
1%
#143620000000
0!
0%
#143625000000
1!
1%
#143630000000
0!
0%
#143635000000
1!
1%
#143640000000
0!
0%
#143645000000
1!
1%
#143650000000
0!
0%
#143655000000
1!
1%
#143660000000
0!
0%
#143665000000
1!
1%
#143670000000
0!
0%
#143675000000
1!
1%
#143680000000
0!
0%
#143685000000
1!
1%
#143690000000
0!
0%
#143695000000
1!
1%
#143700000000
0!
0%
#143705000000
1!
1%
#143710000000
0!
0%
#143715000000
1!
1%
#143720000000
0!
0%
#143725000000
1!
1%
#143730000000
0!
0%
#143735000000
1!
1%
#143740000000
0!
0%
#143745000000
1!
1%
#143750000000
0!
0%
#143755000000
1!
1%
#143760000000
0!
0%
#143765000000
1!
1%
#143770000000
0!
0%
#143775000000
1!
1%
#143780000000
0!
0%
#143785000000
1!
1%
#143790000000
0!
0%
#143795000000
1!
1%
#143800000000
0!
0%
#143805000000
1!
1%
#143810000000
0!
0%
#143815000000
1!
1%
#143820000000
0!
0%
#143825000000
1!
1%
#143830000000
0!
0%
#143835000000
1!
1%
#143840000000
0!
0%
#143845000000
1!
1%
#143850000000
0!
0%
#143855000000
1!
1%
#143860000000
0!
0%
#143865000000
1!
1%
#143870000000
0!
0%
#143875000000
1!
1%
#143880000000
0!
0%
#143885000000
1!
1%
#143890000000
0!
0%
#143895000000
1!
1%
#143900000000
0!
0%
#143905000000
1!
1%
#143910000000
0!
0%
#143915000000
1!
1%
#143920000000
0!
0%
#143925000000
1!
1%
#143930000000
0!
0%
#143935000000
1!
1%
#143940000000
0!
0%
#143945000000
1!
1%
#143950000000
0!
0%
#143955000000
1!
1%
#143960000000
0!
0%
#143965000000
1!
1%
#143970000000
0!
0%
#143975000000
1!
1%
#143980000000
0!
0%
#143985000000
1!
1%
#143990000000
0!
0%
#143995000000
1!
1%
#144000000000
0!
0%
#144005000000
1!
1%
#144010000000
0!
0%
#144015000000
1!
1%
#144020000000
0!
0%
#144025000000
1!
1%
#144030000000
0!
0%
#144035000000
1!
1%
#144040000000
0!
0%
#144045000000
1!
1%
#144050000000
0!
0%
#144055000000
1!
1%
#144060000000
0!
0%
#144065000000
1!
1%
#144070000000
0!
0%
#144075000000
1!
1%
#144080000000
0!
0%
#144085000000
1!
1%
#144090000000
0!
0%
#144095000000
1!
1%
#144100000000
0!
0%
#144105000000
1!
1%
#144110000000
0!
0%
#144115000000
1!
1%
#144120000000
0!
0%
#144125000000
1!
1%
#144130000000
0!
0%
#144135000000
1!
1%
#144140000000
0!
0%
#144145000000
1!
1%
#144150000000
0!
0%
#144155000000
1!
1%
#144160000000
0!
0%
#144165000000
1!
1%
#144170000000
0!
0%
#144175000000
1!
1%
#144180000000
0!
0%
#144185000000
1!
1%
#144190000000
0!
0%
#144195000000
1!
1%
#144200000000
0!
0%
#144205000000
1!
1%
#144210000000
0!
0%
#144215000000
1!
1%
#144220000000
0!
0%
#144225000000
1!
1%
#144230000000
0!
0%
#144235000000
1!
1%
#144240000000
0!
0%
#144245000000
1!
1%
#144250000000
0!
0%
#144255000000
1!
1%
#144260000000
0!
0%
#144265000000
1!
1%
#144270000000
0!
0%
#144275000000
1!
1%
#144280000000
0!
0%
#144285000000
1!
1%
#144290000000
0!
0%
#144295000000
1!
1%
#144300000000
0!
0%
#144305000000
1!
1%
#144310000000
0!
0%
#144315000000
1!
1%
#144320000000
0!
0%
#144325000000
1!
1%
#144330000000
0!
0%
#144335000000
1!
1%
#144340000000
0!
0%
#144345000000
1!
1%
#144350000000
0!
0%
#144355000000
1!
1%
#144360000000
0!
0%
#144365000000
1!
1%
#144370000000
0!
0%
#144375000000
1!
1%
#144380000000
0!
0%
#144385000000
1!
1%
#144390000000
0!
0%
#144395000000
1!
1%
#144400000000
0!
0%
#144405000000
1!
1%
#144410000000
0!
0%
#144415000000
1!
1%
#144420000000
0!
0%
#144425000000
1!
1%
#144430000000
0!
0%
#144435000000
1!
1%
#144440000000
0!
0%
#144445000000
1!
1%
#144450000000
0!
0%
#144455000000
1!
1%
#144460000000
0!
0%
#144465000000
1!
1%
#144470000000
0!
0%
#144475000000
1!
1%
#144480000000
0!
0%
#144485000000
1!
1%
#144490000000
0!
0%
#144495000000
1!
1%
#144500000000
0!
0%
#144505000000
1!
1%
#144510000000
0!
0%
#144515000000
1!
1%
#144520000000
0!
0%
#144525000000
1!
1%
#144530000000
0!
0%
#144535000000
1!
1%
#144540000000
0!
0%
#144545000000
1!
1%
#144550000000
0!
0%
#144555000000
1!
1%
#144560000000
0!
0%
#144565000000
1!
1%
#144570000000
0!
0%
#144575000000
1!
1%
#144580000000
0!
0%
#144585000000
1!
1%
#144590000000
0!
0%
#144595000000
1!
1%
#144600000000
0!
0%
#144605000000
1!
1%
#144610000000
0!
0%
#144615000000
1!
1%
#144620000000
0!
0%
#144625000000
1!
1%
#144630000000
0!
0%
#144635000000
1!
1%
#144640000000
0!
0%
#144645000000
1!
1%
#144650000000
0!
0%
#144655000000
1!
1%
#144660000000
0!
0%
#144665000000
1!
1%
#144670000000
0!
0%
#144675000000
1!
1%
#144680000000
0!
0%
#144685000000
1!
1%
#144690000000
0!
0%
#144695000000
1!
1%
#144700000000
0!
0%
#144705000000
1!
1%
#144710000000
0!
0%
#144715000000
1!
1%
#144720000000
0!
0%
#144725000000
1!
1%
#144730000000
0!
0%
#144735000000
1!
1%
#144740000000
0!
0%
#144745000000
1!
1%
#144750000000
0!
0%
#144755000000
1!
1%
#144760000000
0!
0%
#144765000000
1!
1%
#144770000000
0!
0%
#144775000000
1!
1%
#144780000000
0!
0%
#144785000000
1!
1%
#144790000000
0!
0%
#144795000000
1!
1%
#144800000000
0!
0%
#144805000000
1!
1%
#144810000000
0!
0%
#144815000000
1!
1%
#144820000000
0!
0%
#144825000000
1!
1%
#144830000000
0!
0%
#144835000000
1!
1%
#144840000000
0!
0%
#144845000000
1!
1%
#144850000000
0!
0%
#144855000000
1!
1%
#144860000000
0!
0%
#144865000000
1!
1%
#144870000000
0!
0%
#144875000000
1!
1%
#144880000000
0!
0%
#144885000000
1!
1%
#144890000000
0!
0%
#144895000000
1!
1%
#144900000000
0!
0%
#144905000000
1!
1%
#144910000000
0!
0%
#144915000000
1!
1%
#144920000000
0!
0%
#144925000000
1!
1%
#144930000000
0!
0%
#144935000000
1!
1%
#144940000000
0!
0%
#144945000000
1!
1%
#144950000000
0!
0%
#144955000000
1!
1%
#144960000000
0!
0%
#144965000000
1!
1%
#144970000000
0!
0%
#144975000000
1!
1%
#144980000000
0!
0%
#144985000000
1!
1%
#144990000000
0!
0%
#144995000000
1!
1%
#145000000000
0!
0%
#145005000000
1!
1%
#145010000000
0!
0%
#145015000000
1!
1%
#145020000000
0!
0%
#145025000000
1!
1%
#145030000000
0!
0%
#145035000000
1!
1%
#145040000000
0!
0%
#145045000000
1!
1%
#145050000000
0!
0%
#145055000000
1!
1%
#145060000000
0!
0%
#145065000000
1!
1%
#145070000000
0!
0%
#145075000000
1!
1%
#145080000000
0!
0%
#145085000000
1!
1%
#145090000000
0!
0%
#145095000000
1!
1%
#145100000000
0!
0%
#145105000000
1!
1%
#145110000000
0!
0%
#145115000000
1!
1%
#145120000000
0!
0%
#145125000000
1!
1%
#145130000000
0!
0%
#145135000000
1!
1%
#145140000000
0!
0%
#145145000000
1!
1%
#145150000000
0!
0%
#145155000000
1!
1%
#145160000000
0!
0%
#145165000000
1!
1%
#145170000000
0!
0%
#145175000000
1!
1%
#145180000000
0!
0%
#145185000000
1!
1%
#145190000000
0!
0%
#145195000000
1!
1%
#145200000000
0!
0%
#145205000000
1!
1%
#145210000000
0!
0%
#145215000000
1!
1%
#145220000000
0!
0%
#145225000000
1!
1%
#145230000000
0!
0%
#145235000000
1!
1%
#145240000000
0!
0%
#145245000000
1!
1%
#145250000000
0!
0%
#145255000000
1!
1%
#145260000000
0!
0%
#145265000000
1!
1%
#145270000000
0!
0%
#145275000000
1!
1%
#145280000000
0!
0%
#145285000000
1!
1%
#145290000000
0!
0%
#145295000000
1!
1%
#145300000000
0!
0%
#145305000000
1!
1%
#145310000000
0!
0%
#145315000000
1!
1%
#145320000000
0!
0%
#145325000000
1!
1%
#145330000000
0!
0%
#145335000000
1!
1%
#145340000000
0!
0%
#145345000000
1!
1%
#145350000000
0!
0%
#145355000000
1!
1%
#145360000000
0!
0%
#145365000000
1!
1%
#145370000000
0!
0%
#145375000000
1!
1%
#145380000000
0!
0%
#145385000000
1!
1%
#145390000000
0!
0%
#145395000000
1!
1%
#145400000000
0!
0%
#145405000000
1!
1%
#145410000000
0!
0%
#145415000000
1!
1%
#145420000000
0!
0%
#145425000000
1!
1%
#145430000000
0!
0%
#145435000000
1!
1%
#145440000000
0!
0%
#145445000000
1!
1%
#145450000000
0!
0%
#145455000000
1!
1%
#145460000000
0!
0%
#145465000000
1!
1%
#145470000000
0!
0%
#145475000000
1!
1%
#145480000000
0!
0%
#145485000000
1!
1%
#145490000000
0!
0%
#145495000000
1!
1%
#145500000000
0!
0%
#145505000000
1!
1%
#145510000000
0!
0%
#145515000000
1!
1%
#145520000000
0!
0%
#145525000000
1!
1%
#145530000000
0!
0%
#145535000000
1!
1%
#145540000000
0!
0%
#145545000000
1!
1%
#145550000000
0!
0%
#145555000000
1!
1%
#145560000000
0!
0%
#145565000000
1!
1%
#145570000000
0!
0%
#145575000000
1!
1%
#145580000000
0!
0%
#145585000000
1!
1%
#145590000000
0!
0%
#145595000000
1!
1%
#145600000000
0!
0%
#145605000000
1!
1%
#145610000000
0!
0%
#145615000000
1!
1%
#145620000000
0!
0%
#145625000000
1!
1%
#145630000000
0!
0%
#145635000000
1!
1%
#145640000000
0!
0%
#145645000000
1!
1%
#145650000000
0!
0%
#145655000000
1!
1%
#145660000000
0!
0%
#145665000000
1!
1%
#145670000000
0!
0%
#145675000000
1!
1%
#145680000000
0!
0%
#145685000000
1!
1%
#145690000000
0!
0%
#145695000000
1!
1%
#145700000000
0!
0%
#145705000000
1!
1%
#145710000000
0!
0%
#145715000000
1!
1%
#145720000000
0!
0%
#145725000000
1!
1%
#145730000000
0!
0%
#145735000000
1!
1%
#145740000000
0!
0%
#145745000000
1!
1%
#145750000000
0!
0%
#145755000000
1!
1%
#145760000000
0!
0%
#145765000000
1!
1%
#145770000000
0!
0%
#145775000000
1!
1%
#145780000000
0!
0%
#145785000000
1!
1%
#145790000000
0!
0%
#145795000000
1!
1%
#145800000000
0!
0%
#145805000000
1!
1%
#145810000000
0!
0%
#145815000000
1!
1%
#145820000000
0!
0%
#145825000000
1!
1%
#145830000000
0!
0%
#145835000000
1!
1%
#145840000000
0!
0%
#145845000000
1!
1%
#145850000000
0!
0%
#145855000000
1!
1%
#145860000000
0!
0%
#145865000000
1!
1%
#145870000000
0!
0%
#145875000000
1!
1%
#145880000000
0!
0%
#145885000000
1!
1%
#145890000000
0!
0%
#145895000000
1!
1%
#145900000000
0!
0%
#145905000000
1!
1%
#145910000000
0!
0%
#145915000000
1!
1%
#145920000000
0!
0%
#145925000000
1!
1%
#145930000000
0!
0%
#145935000000
1!
1%
#145940000000
0!
0%
#145945000000
1!
1%
#145950000000
0!
0%
#145955000000
1!
1%
#145960000000
0!
0%
#145965000000
1!
1%
#145970000000
0!
0%
#145975000000
1!
1%
#145980000000
0!
0%
#145985000000
1!
1%
#145990000000
0!
0%
#145995000000
1!
1%
#146000000000
0!
0%
#146005000000
1!
1%
#146010000000
0!
0%
#146015000000
1!
1%
#146020000000
0!
0%
#146025000000
1!
1%
#146030000000
0!
0%
#146035000000
1!
1%
#146040000000
0!
0%
#146045000000
1!
1%
#146050000000
0!
0%
#146055000000
1!
1%
#146060000000
0!
0%
#146065000000
1!
1%
#146070000000
0!
0%
#146075000000
1!
1%
#146080000000
0!
0%
#146085000000
1!
1%
#146090000000
0!
0%
#146095000000
1!
1%
#146100000000
0!
0%
#146105000000
1!
1%
#146110000000
0!
0%
#146115000000
1!
1%
#146120000000
0!
0%
#146125000000
1!
1%
#146130000000
0!
0%
#146135000000
1!
1%
#146140000000
0!
0%
#146145000000
1!
1%
#146150000000
0!
0%
#146155000000
1!
1%
#146160000000
0!
0%
#146165000000
1!
1%
#146170000000
0!
0%
#146175000000
1!
1%
#146180000000
0!
0%
#146185000000
1!
1%
#146190000000
0!
0%
#146195000000
1!
1%
#146200000000
0!
0%
#146205000000
1!
1%
#146210000000
0!
0%
#146215000000
1!
1%
#146220000000
0!
0%
#146225000000
1!
1%
#146230000000
0!
0%
#146235000000
1!
1%
#146240000000
0!
0%
#146245000000
1!
1%
#146250000000
0!
0%
#146255000000
1!
1%
#146260000000
0!
0%
#146265000000
1!
1%
#146270000000
0!
0%
#146275000000
1!
1%
#146280000000
0!
0%
#146285000000
1!
1%
#146290000000
0!
0%
#146295000000
1!
1%
#146300000000
0!
0%
#146305000000
1!
1%
#146310000000
0!
0%
#146315000000
1!
1%
#146320000000
0!
0%
#146325000000
1!
1%
#146330000000
0!
0%
#146335000000
1!
1%
#146340000000
0!
0%
#146345000000
1!
1%
#146350000000
0!
0%
#146355000000
1!
1%
#146360000000
0!
0%
#146365000000
1!
1%
#146370000000
0!
0%
#146375000000
1!
1%
#146380000000
0!
0%
#146385000000
1!
1%
#146390000000
0!
0%
#146395000000
1!
1%
#146400000000
0!
0%
#146405000000
1!
1%
#146410000000
0!
0%
#146415000000
1!
1%
#146420000000
0!
0%
#146425000000
1!
1%
#146430000000
0!
0%
#146435000000
1!
1%
#146440000000
0!
0%
#146445000000
1!
1%
#146450000000
0!
0%
#146455000000
1!
1%
#146460000000
0!
0%
#146465000000
1!
1%
#146470000000
0!
0%
#146475000000
1!
1%
#146480000000
0!
0%
#146485000000
1!
1%
#146490000000
0!
0%
#146495000000
1!
1%
#146500000000
0!
0%
#146505000000
1!
1%
#146510000000
0!
0%
#146515000000
1!
1%
#146520000000
0!
0%
#146525000000
1!
1%
#146530000000
0!
0%
#146535000000
1!
1%
#146540000000
0!
0%
#146545000000
1!
1%
#146550000000
0!
0%
#146555000000
1!
1%
#146560000000
0!
0%
#146565000000
1!
1%
#146570000000
0!
0%
#146575000000
1!
1%
#146580000000
0!
0%
#146585000000
1!
1%
#146590000000
0!
0%
#146595000000
1!
1%
#146600000000
0!
0%
#146605000000
1!
1%
#146610000000
0!
0%
#146615000000
1!
1%
#146620000000
0!
0%
#146625000000
1!
1%
#146630000000
0!
0%
#146635000000
1!
1%
#146640000000
0!
0%
#146645000000
1!
1%
#146650000000
0!
0%
#146655000000
1!
1%
#146660000000
0!
0%
#146665000000
1!
1%
#146670000000
0!
0%
#146675000000
1!
1%
#146680000000
0!
0%
#146685000000
1!
1%
#146690000000
0!
0%
#146695000000
1!
1%
#146700000000
0!
0%
#146705000000
1!
1%
#146710000000
0!
0%
#146715000000
1!
1%
#146720000000
0!
0%
#146725000000
1!
1%
#146730000000
0!
0%
#146735000000
1!
1%
#146740000000
0!
0%
#146745000000
1!
1%
#146750000000
0!
0%
#146755000000
1!
1%
#146760000000
0!
0%
#146765000000
1!
1%
#146770000000
0!
0%
#146775000000
1!
1%
#146780000000
0!
0%
#146785000000
1!
1%
#146790000000
0!
0%
#146795000000
1!
1%
#146800000000
0!
0%
#146805000000
1!
1%
#146810000000
0!
0%
#146815000000
1!
1%
#146820000000
0!
0%
#146825000000
1!
1%
#146830000000
0!
0%
#146835000000
1!
1%
#146840000000
0!
0%
#146845000000
1!
1%
#146850000000
0!
0%
#146855000000
1!
1%
#146860000000
0!
0%
#146865000000
1!
1%
#146870000000
0!
0%
#146875000000
1!
1%
#146880000000
0!
0%
#146885000000
1!
1%
#146890000000
0!
0%
#146895000000
1!
1%
#146900000000
0!
0%
#146905000000
1!
1%
#146910000000
0!
0%
#146915000000
1!
1%
#146920000000
0!
0%
#146925000000
1!
1%
#146930000000
0!
0%
#146935000000
1!
1%
#146940000000
0!
0%
#146945000000
1!
1%
#146950000000
0!
0%
#146955000000
1!
1%
#146960000000
0!
0%
#146965000000
1!
1%
#146970000000
0!
0%
#146975000000
1!
1%
#146980000000
0!
0%
#146985000000
1!
1%
#146990000000
0!
0%
#146995000000
1!
1%
#147000000000
0!
0%
#147005000000
1!
1%
#147010000000
0!
0%
#147015000000
1!
1%
#147020000000
0!
0%
#147025000000
1!
1%
#147030000000
0!
0%
#147035000000
1!
1%
#147040000000
0!
0%
#147045000000
1!
1%
#147050000000
0!
0%
#147055000000
1!
1%
#147060000000
0!
0%
#147065000000
1!
1%
#147070000000
0!
0%
#147075000000
1!
1%
#147080000000
0!
0%
#147085000000
1!
1%
#147090000000
0!
0%
#147095000000
1!
1%
#147100000000
0!
0%
#147105000000
1!
1%
#147110000000
0!
0%
#147115000000
1!
1%
#147120000000
0!
0%
#147125000000
1!
1%
#147130000000
0!
0%
#147135000000
1!
1%
#147140000000
0!
0%
#147145000000
1!
1%
#147150000000
0!
0%
#147155000000
1!
1%
#147160000000
0!
0%
#147165000000
1!
1%
#147170000000
0!
0%
#147175000000
1!
1%
#147180000000
0!
0%
#147185000000
1!
1%
#147190000000
0!
0%
#147195000000
1!
1%
#147200000000
0!
0%
#147205000000
1!
1%
#147210000000
0!
0%
#147215000000
1!
1%
#147220000000
0!
0%
#147225000000
1!
1%
#147230000000
0!
0%
#147235000000
1!
1%
#147240000000
0!
0%
#147245000000
1!
1%
#147250000000
0!
0%
#147255000000
1!
1%
#147260000000
0!
0%
#147265000000
1!
1%
#147270000000
0!
0%
#147275000000
1!
1%
#147280000000
0!
0%
#147285000000
1!
1%
#147290000000
0!
0%
#147295000000
1!
1%
#147300000000
0!
0%
#147305000000
1!
1%
#147310000000
0!
0%
#147315000000
1!
1%
#147320000000
0!
0%
#147325000000
1!
1%
#147330000000
0!
0%
#147335000000
1!
1%
#147340000000
0!
0%
#147345000000
1!
1%
#147350000000
0!
0%
#147355000000
1!
1%
#147360000000
0!
0%
#147365000000
1!
1%
#147370000000
0!
0%
#147375000000
1!
1%
#147380000000
0!
0%
#147385000000
1!
1%
#147390000000
0!
0%
#147395000000
1!
1%
#147400000000
0!
0%
#147405000000
1!
1%
#147410000000
0!
0%
#147415000000
1!
1%
#147420000000
0!
0%
#147425000000
1!
1%
#147430000000
0!
0%
#147435000000
1!
1%
#147440000000
0!
0%
#147445000000
1!
1%
#147450000000
0!
0%
#147455000000
1!
1%
#147460000000
0!
0%
#147465000000
1!
1%
#147470000000
0!
0%
#147475000000
1!
1%
#147480000000
0!
0%
#147485000000
1!
1%
#147490000000
0!
0%
#147495000000
1!
1%
#147500000000
0!
0%
#147505000000
1!
1%
#147510000000
0!
0%
#147515000000
1!
1%
#147520000000
0!
0%
#147525000000
1!
1%
#147530000000
0!
0%
#147535000000
1!
1%
#147540000000
0!
0%
#147545000000
1!
1%
#147550000000
0!
0%
#147555000000
1!
1%
#147560000000
0!
0%
#147565000000
1!
1%
#147570000000
0!
0%
#147575000000
1!
1%
#147580000000
0!
0%
#147585000000
1!
1%
#147590000000
0!
0%
#147595000000
1!
1%
#147600000000
0!
0%
#147605000000
1!
1%
#147610000000
0!
0%
#147615000000
1!
1%
#147620000000
0!
0%
#147625000000
1!
1%
#147630000000
0!
0%
#147635000000
1!
1%
#147640000000
0!
0%
#147645000000
1!
1%
#147650000000
0!
0%
#147655000000
1!
1%
#147660000000
0!
0%
#147665000000
1!
1%
#147670000000
0!
0%
#147675000000
1!
1%
#147680000000
0!
0%
#147685000000
1!
1%
#147690000000
0!
0%
#147695000000
1!
1%
#147700000000
0!
0%
#147705000000
1!
1%
#147710000000
0!
0%
#147715000000
1!
1%
#147720000000
0!
0%
#147725000000
1!
1%
#147730000000
0!
0%
#147735000000
1!
1%
#147740000000
0!
0%
#147745000000
1!
1%
#147750000000
0!
0%
#147755000000
1!
1%
#147760000000
0!
0%
#147765000000
1!
1%
#147770000000
0!
0%
#147775000000
1!
1%
#147780000000
0!
0%
#147785000000
1!
1%
#147790000000
0!
0%
#147795000000
1!
1%
#147800000000
0!
0%
#147805000000
1!
1%
#147810000000
0!
0%
#147815000000
1!
1%
#147820000000
0!
0%
#147825000000
1!
1%
#147830000000
0!
0%
#147835000000
1!
1%
#147840000000
0!
0%
#147845000000
1!
1%
#147850000000
0!
0%
#147855000000
1!
1%
#147860000000
0!
0%
#147865000000
1!
1%
#147870000000
0!
0%
#147875000000
1!
1%
#147880000000
0!
0%
#147885000000
1!
1%
#147890000000
0!
0%
#147895000000
1!
1%
#147900000000
0!
0%
#147905000000
1!
1%
#147910000000
0!
0%
#147915000000
1!
1%
#147920000000
0!
0%
#147925000000
1!
1%
#147930000000
0!
0%
#147935000000
1!
1%
#147940000000
0!
0%
#147945000000
1!
1%
#147950000000
0!
0%
#147955000000
1!
1%
#147960000000
0!
0%
#147965000000
1!
1%
#147970000000
0!
0%
#147975000000
1!
1%
#147980000000
0!
0%
#147985000000
1!
1%
#147990000000
0!
0%
#147995000000
1!
1%
#148000000000
0!
0%
#148005000000
1!
1%
#148010000000
0!
0%
#148015000000
1!
1%
#148020000000
0!
0%
#148025000000
1!
1%
#148030000000
0!
0%
#148035000000
1!
1%
#148040000000
0!
0%
#148045000000
1!
1%
#148050000000
0!
0%
#148055000000
1!
1%
#148060000000
0!
0%
#148065000000
1!
1%
#148070000000
0!
0%
#148075000000
1!
1%
#148080000000
0!
0%
#148085000000
1!
1%
#148090000000
0!
0%
#148095000000
1!
1%
#148100000000
0!
0%
#148105000000
1!
1%
#148110000000
0!
0%
#148115000000
1!
1%
#148120000000
0!
0%
#148125000000
1!
1%
#148130000000
0!
0%
#148135000000
1!
1%
#148140000000
0!
0%
#148145000000
1!
1%
#148150000000
0!
0%
#148155000000
1!
1%
#148160000000
0!
0%
#148165000000
1!
1%
#148170000000
0!
0%
#148175000000
1!
1%
#148180000000
0!
0%
#148185000000
1!
1%
#148190000000
0!
0%
#148195000000
1!
1%
#148200000000
0!
0%
#148205000000
1!
1%
#148210000000
0!
0%
#148215000000
1!
1%
#148220000000
0!
0%
#148225000000
1!
1%
#148230000000
0!
0%
#148235000000
1!
1%
#148240000000
0!
0%
#148245000000
1!
1%
#148250000000
0!
0%
#148255000000
1!
1%
#148260000000
0!
0%
#148265000000
1!
1%
#148270000000
0!
0%
#148275000000
1!
1%
#148280000000
0!
0%
#148285000000
1!
1%
#148290000000
0!
0%
#148295000000
1!
1%
#148300000000
0!
0%
#148305000000
1!
1%
#148310000000
0!
0%
#148315000000
1!
1%
#148320000000
0!
0%
#148325000000
1!
1%
#148330000000
0!
0%
#148335000000
1!
1%
#148340000000
0!
0%
#148345000000
1!
1%
#148350000000
0!
0%
#148355000000
1!
1%
#148360000000
0!
0%
#148365000000
1!
1%
#148370000000
0!
0%
#148375000000
1!
1%
#148380000000
0!
0%
#148385000000
1!
1%
#148390000000
0!
0%
#148395000000
1!
1%
#148400000000
0!
0%
#148405000000
1!
1%
#148410000000
0!
0%
#148415000000
1!
1%
#148420000000
0!
0%
#148425000000
1!
1%
#148430000000
0!
0%
#148435000000
1!
1%
#148440000000
0!
0%
#148445000000
1!
1%
#148450000000
0!
0%
#148455000000
1!
1%
#148460000000
0!
0%
#148465000000
1!
1%
#148470000000
0!
0%
#148475000000
1!
1%
#148480000000
0!
0%
#148485000000
1!
1%
#148490000000
0!
0%
#148495000000
1!
1%
#148500000000
0!
0%
#148505000000
1!
1%
#148510000000
0!
0%
#148515000000
1!
1%
#148520000000
0!
0%
#148525000000
1!
1%
#148530000000
0!
0%
#148535000000
1!
1%
#148540000000
0!
0%
#148545000000
1!
1%
#148550000000
0!
0%
#148555000000
1!
1%
#148560000000
0!
0%
#148565000000
1!
1%
#148570000000
0!
0%
#148575000000
1!
1%
#148580000000
0!
0%
#148585000000
1!
1%
#148590000000
0!
0%
#148595000000
1!
1%
#148600000000
0!
0%
#148605000000
1!
1%
#148610000000
0!
0%
#148615000000
1!
1%
#148620000000
0!
0%
#148625000000
1!
1%
#148630000000
0!
0%
#148635000000
1!
1%
#148640000000
0!
0%
#148645000000
1!
1%
#148650000000
0!
0%
#148655000000
1!
1%
#148660000000
0!
0%
#148665000000
1!
1%
#148670000000
0!
0%
#148675000000
1!
1%
#148680000000
0!
0%
#148685000000
1!
1%
#148690000000
0!
0%
#148695000000
1!
1%
#148700000000
0!
0%
#148705000000
1!
1%
#148710000000
0!
0%
#148715000000
1!
1%
#148720000000
0!
0%
#148725000000
1!
1%
#148730000000
0!
0%
#148735000000
1!
1%
#148740000000
0!
0%
#148745000000
1!
1%
#148750000000
0!
0%
#148755000000
1!
1%
#148760000000
0!
0%
#148765000000
1!
1%
#148770000000
0!
0%
#148775000000
1!
1%
#148780000000
0!
0%
#148785000000
1!
1%
#148790000000
0!
0%
#148795000000
1!
1%
#148800000000
0!
0%
#148805000000
1!
1%
#148810000000
0!
0%
#148815000000
1!
1%
#148820000000
0!
0%
#148825000000
1!
1%
#148830000000
0!
0%
#148835000000
1!
1%
#148840000000
0!
0%
#148845000000
1!
1%
#148850000000
0!
0%
#148855000000
1!
1%
#148860000000
0!
0%
#148865000000
1!
1%
#148870000000
0!
0%
#148875000000
1!
1%
#148880000000
0!
0%
#148885000000
1!
1%
#148890000000
0!
0%
#148895000000
1!
1%
#148900000000
0!
0%
#148905000000
1!
1%
#148910000000
0!
0%
#148915000000
1!
1%
#148920000000
0!
0%
#148925000000
1!
1%
#148930000000
0!
0%
#148935000000
1!
1%
#148940000000
0!
0%
#148945000000
1!
1%
#148950000000
0!
0%
#148955000000
1!
1%
#148960000000
0!
0%
#148965000000
1!
1%
#148970000000
0!
0%
#148975000000
1!
1%
#148980000000
0!
0%
#148985000000
1!
1%
#148990000000
0!
0%
#148995000000
1!
1%
#149000000000
0!
0%
#149005000000
1!
1%
#149010000000
0!
0%
#149015000000
1!
1%
#149020000000
0!
0%
#149025000000
1!
1%
#149030000000
0!
0%
#149035000000
1!
1%
#149040000000
0!
0%
#149045000000
1!
1%
#149050000000
0!
0%
#149055000000
1!
1%
#149060000000
0!
0%
#149065000000
1!
1%
#149070000000
0!
0%
#149075000000
1!
1%
#149080000000
0!
0%
#149085000000
1!
1%
#149090000000
0!
0%
#149095000000
1!
1%
#149100000000
0!
0%
#149105000000
1!
1%
#149110000000
0!
0%
#149115000000
1!
1%
#149120000000
0!
0%
#149125000000
1!
1%
#149130000000
0!
0%
#149135000000
1!
1%
#149140000000
0!
0%
#149145000000
1!
1%
#149150000000
0!
0%
#149155000000
1!
1%
#149160000000
0!
0%
#149165000000
1!
1%
#149170000000
0!
0%
#149175000000
1!
1%
#149180000000
0!
0%
#149185000000
1!
1%
#149190000000
0!
0%
#149195000000
1!
1%
#149200000000
0!
0%
#149205000000
1!
1%
#149210000000
0!
0%
#149215000000
1!
1%
#149220000000
0!
0%
#149225000000
1!
1%
#149230000000
0!
0%
#149235000000
1!
1%
#149240000000
0!
0%
#149245000000
1!
1%
#149250000000
0!
0%
#149255000000
1!
1%
#149260000000
0!
0%
#149265000000
1!
1%
#149270000000
0!
0%
#149275000000
1!
1%
#149280000000
0!
0%
#149285000000
1!
1%
#149290000000
0!
0%
#149295000000
1!
1%
#149300000000
0!
0%
#149305000000
1!
1%
#149310000000
0!
0%
#149315000000
1!
1%
#149320000000
0!
0%
#149325000000
1!
1%
#149330000000
0!
0%
#149335000000
1!
1%
#149340000000
0!
0%
#149345000000
1!
1%
#149350000000
0!
0%
#149355000000
1!
1%
#149360000000
0!
0%
#149365000000
1!
1%
#149370000000
0!
0%
#149375000000
1!
1%
#149380000000
0!
0%
#149385000000
1!
1%
#149390000000
0!
0%
#149395000000
1!
1%
#149400000000
0!
0%
#149405000000
1!
1%
#149410000000
0!
0%
#149415000000
1!
1%
#149420000000
0!
0%
#149425000000
1!
1%
#149430000000
0!
0%
#149435000000
1!
1%
#149440000000
0!
0%
#149445000000
1!
1%
#149450000000
0!
0%
#149455000000
1!
1%
#149460000000
0!
0%
#149465000000
1!
1%
#149470000000
0!
0%
#149475000000
1!
1%
#149480000000
0!
0%
#149485000000
1!
1%
#149490000000
0!
0%
#149495000000
1!
1%
#149500000000
0!
0%
#149505000000
1!
1%
#149510000000
0!
0%
#149515000000
1!
1%
#149520000000
0!
0%
#149525000000
1!
1%
#149530000000
0!
0%
#149535000000
1!
1%
#149540000000
0!
0%
#149545000000
1!
1%
#149550000000
0!
0%
#149555000000
1!
1%
#149560000000
0!
0%
#149565000000
1!
1%
#149570000000
0!
0%
#149575000000
1!
1%
#149580000000
0!
0%
#149585000000
1!
1%
#149590000000
0!
0%
#149595000000
1!
1%
#149600000000
0!
0%
#149605000000
1!
1%
#149610000000
0!
0%
#149615000000
1!
1%
#149620000000
0!
0%
#149625000000
1!
1%
#149630000000
0!
0%
#149635000000
1!
1%
#149640000000
0!
0%
#149645000000
1!
1%
#149650000000
0!
0%
#149655000000
1!
1%
#149660000000
0!
0%
#149665000000
1!
1%
#149670000000
0!
0%
#149675000000
1!
1%
#149680000000
0!
0%
#149685000000
1!
1%
#149690000000
0!
0%
#149695000000
1!
1%
#149700000000
0!
0%
#149705000000
1!
1%
#149710000000
0!
0%
#149715000000
1!
1%
#149720000000
0!
0%
#149725000000
1!
1%
#149730000000
0!
0%
#149735000000
1!
1%
#149740000000
0!
0%
#149745000000
1!
1%
#149750000000
0!
0%
#149755000000
1!
1%
#149760000000
0!
0%
#149765000000
1!
1%
#149770000000
0!
0%
#149775000000
1!
1%
#149780000000
0!
0%
#149785000000
1!
1%
#149790000000
0!
0%
#149795000000
1!
1%
#149800000000
0!
0%
#149805000000
1!
1%
#149810000000
0!
0%
#149815000000
1!
1%
#149820000000
0!
0%
#149825000000
1!
1%
#149830000000
0!
0%
#149835000000
1!
1%
#149840000000
0!
0%
#149845000000
1!
1%
#149850000000
0!
0%
#149855000000
1!
1%
#149860000000
0!
0%
#149865000000
1!
1%
#149870000000
0!
0%
#149875000000
1!
1%
#149880000000
0!
0%
#149885000000
1!
1%
#149890000000
0!
0%
#149895000000
1!
1%
#149900000000
0!
0%
#149905000000
1!
1%
#149910000000
0!
0%
#149915000000
1!
1%
#149920000000
0!
0%
#149925000000
1!
1%
#149930000000
0!
0%
#149935000000
1!
1%
#149940000000
0!
0%
#149945000000
1!
1%
#149950000000
0!
0%
#149955000000
1!
1%
#149960000000
0!
0%
#149965000000
1!
1%
#149970000000
0!
0%
#149975000000
1!
1%
#149980000000
0!
0%
#149985000000
1!
1%
#149990000000
0!
0%
#149995000000
1!
1%
#150000000000
0!
0%
#150005000000
1!
1%
#150010000000
0!
0%
#150015000000
1!
1%
#150020000000
0!
0%
#150025000000
1!
1%
#150030000000
0!
0%
#150035000000
1!
1%
#150040000000
0!
0%
#150045000000
1!
1%
#150050000000
0!
0%
#150055000000
1!
1%
#150060000000
0!
0%
#150065000000
1!
1%
#150070000000
0!
0%
#150075000000
1!
1%
#150080000000
0!
0%
#150085000000
1!
1%
#150090000000
0!
0%
#150095000000
1!
1%
#150100000000
0!
0%
#150105000000
1!
1%
#150110000000
0!
0%
#150115000000
1!
1%
#150120000000
0!
0%
#150125000000
1!
1%
#150130000000
0!
0%
#150135000000
1!
1%
#150140000000
0!
0%
#150145000000
1!
1%
#150150000000
0!
0%
#150155000000
1!
1%
#150160000000
0!
0%
#150165000000
1!
1%
#150170000000
0!
0%
#150175000000
1!
1%
#150180000000
0!
0%
#150185000000
1!
1%
#150190000000
0!
0%
#150195000000
1!
1%
#150200000000
0!
0%
#150205000000
1!
1%
#150210000000
0!
0%
#150215000000
1!
1%
#150220000000
0!
0%
#150225000000
1!
1%
#150230000000
0!
0%
#150235000000
1!
1%
#150240000000
0!
0%
#150245000000
1!
1%
#150250000000
0!
0%
#150255000000
1!
1%
#150260000000
0!
0%
#150265000000
1!
1%
#150270000000
0!
0%
#150275000000
1!
1%
#150280000000
0!
0%
#150285000000
1!
1%
#150290000000
0!
0%
#150295000000
1!
1%
#150300000000
0!
0%
#150305000000
1!
1%
#150310000000
0!
0%
#150315000000
1!
1%
#150320000000
0!
0%
#150325000000
1!
1%
#150330000000
0!
0%
#150335000000
1!
1%
#150340000000
0!
0%
#150345000000
1!
1%
#150350000000
0!
0%
#150355000000
1!
1%
#150360000000
0!
0%
#150365000000
1!
1%
#150370000000
0!
0%
#150375000000
1!
1%
#150380000000
0!
0%
#150385000000
1!
1%
#150390000000
0!
0%
#150395000000
1!
1%
#150400000000
0!
0%
#150405000000
1!
1%
#150410000000
0!
0%
#150415000000
1!
1%
#150420000000
0!
0%
#150425000000
1!
1%
#150430000000
0!
0%
#150435000000
1!
1%
#150440000000
0!
0%
#150445000000
1!
1%
#150450000000
0!
0%
#150455000000
1!
1%
#150460000000
0!
0%
#150465000000
1!
1%
#150470000000
0!
0%
#150475000000
1!
1%
#150480000000
0!
0%
#150485000000
1!
1%
#150490000000
0!
0%
#150495000000
1!
1%
#150500000000
0!
0%
#150505000000
1!
1%
#150510000000
0!
0%
#150515000000
1!
1%
#150520000000
0!
0%
#150525000000
1!
1%
#150530000000
0!
0%
#150535000000
1!
1%
#150540000000
0!
0%
#150545000000
1!
1%
#150550000000
0!
0%
#150555000000
1!
1%
#150560000000
0!
0%
#150565000000
1!
1%
#150570000000
0!
0%
#150575000000
1!
1%
#150580000000
0!
0%
#150585000000
1!
1%
#150590000000
0!
0%
#150595000000
1!
1%
#150600000000
0!
0%
#150605000000
1!
1%
#150610000000
0!
0%
#150615000000
1!
1%
#150620000000
0!
0%
#150625000000
1!
1%
#150630000000
0!
0%
#150635000000
1!
1%
#150640000000
0!
0%
#150645000000
1!
1%
#150650000000
0!
0%
#150655000000
1!
1%
#150660000000
0!
0%
#150665000000
1!
1%
#150670000000
0!
0%
#150675000000
1!
1%
#150680000000
0!
0%
#150685000000
1!
1%
#150690000000
0!
0%
#150695000000
1!
1%
#150700000000
0!
0%
#150705000000
1!
1%
#150710000000
0!
0%
#150715000000
1!
1%
#150720000000
0!
0%
#150725000000
1!
1%
#150730000000
0!
0%
#150735000000
1!
1%
#150740000000
0!
0%
#150745000000
1!
1%
#150750000000
0!
0%
#150755000000
1!
1%
#150760000000
0!
0%
#150765000000
1!
1%
#150770000000
0!
0%
#150775000000
1!
1%
#150780000000
0!
0%
#150785000000
1!
1%
#150790000000
0!
0%
#150795000000
1!
1%
#150800000000
0!
0%
#150805000000
1!
1%
#150810000000
0!
0%
#150815000000
1!
1%
#150820000000
0!
0%
#150825000000
1!
1%
#150830000000
0!
0%
#150835000000
1!
1%
#150840000000
0!
0%
#150845000000
1!
1%
#150850000000
0!
0%
#150855000000
1!
1%
#150860000000
0!
0%
#150865000000
1!
1%
#150870000000
0!
0%
#150875000000
1!
1%
#150880000000
0!
0%
#150885000000
1!
1%
#150890000000
0!
0%
#150895000000
1!
1%
#150900000000
0!
0%
#150905000000
1!
1%
#150910000000
0!
0%
#150915000000
1!
1%
#150920000000
0!
0%
#150925000000
1!
1%
#150930000000
0!
0%
#150935000000
1!
1%
#150940000000
0!
0%
#150945000000
1!
1%
#150950000000
0!
0%
#150955000000
1!
1%
#150960000000
0!
0%
#150965000000
1!
1%
#150970000000
0!
0%
#150975000000
1!
1%
#150980000000
0!
0%
#150985000000
1!
1%
#150990000000
0!
0%
#150995000000
1!
1%
#151000000000
0!
0%
#151005000000
1!
1%
#151010000000
0!
0%
#151015000000
1!
1%
#151020000000
0!
0%
#151025000000
1!
1%
#151030000000
0!
0%
#151035000000
1!
1%
#151040000000
0!
0%
#151045000000
1!
1%
#151050000000
0!
0%
#151055000000
1!
1%
#151060000000
0!
0%
#151065000000
1!
1%
#151070000000
0!
0%
#151075000000
1!
1%
#151080000000
0!
0%
#151085000000
1!
1%
#151090000000
0!
0%
#151095000000
1!
1%
#151100000000
0!
0%
#151105000000
1!
1%
#151110000000
0!
0%
#151115000000
1!
1%
#151120000000
0!
0%
#151125000000
1!
1%
#151130000000
0!
0%
#151135000000
1!
1%
#151140000000
0!
0%
#151145000000
1!
1%
#151150000000
0!
0%
#151155000000
1!
1%
#151160000000
0!
0%
#151165000000
1!
1%
#151170000000
0!
0%
#151175000000
1!
1%
#151180000000
0!
0%
#151185000000
1!
1%
#151190000000
0!
0%
#151195000000
1!
1%
#151200000000
0!
0%
#151205000000
1!
1%
#151210000000
0!
0%
#151215000000
1!
1%
#151220000000
0!
0%
#151225000000
1!
1%
#151230000000
0!
0%
#151235000000
1!
1%
#151240000000
0!
0%
#151245000000
1!
1%
#151250000000
0!
0%
#151255000000
1!
1%
#151260000000
0!
0%
#151265000000
1!
1%
#151270000000
0!
0%
#151275000000
1!
1%
#151280000000
0!
0%
#151285000000
1!
1%
#151290000000
0!
0%
#151295000000
1!
1%
#151300000000
0!
0%
#151305000000
1!
1%
#151310000000
0!
0%
#151315000000
1!
1%
#151320000000
0!
0%
#151325000000
1!
1%
#151330000000
0!
0%
#151335000000
1!
1%
#151340000000
0!
0%
#151345000000
1!
1%
#151350000000
0!
0%
#151355000000
1!
1%
#151360000000
0!
0%
#151365000000
1!
1%
#151370000000
0!
0%
#151375000000
1!
1%
#151380000000
0!
0%
#151385000000
1!
1%
#151390000000
0!
0%
#151395000000
1!
1%
#151400000000
0!
0%
#151405000000
1!
1%
#151410000000
0!
0%
#151415000000
1!
1%
#151420000000
0!
0%
#151425000000
1!
1%
#151430000000
0!
0%
#151435000000
1!
1%
#151440000000
0!
0%
#151445000000
1!
1%
#151450000000
0!
0%
#151455000000
1!
1%
#151460000000
0!
0%
#151465000000
1!
1%
#151470000000
0!
0%
#151475000000
1!
1%
#151480000000
0!
0%
#151485000000
1!
1%
#151490000000
0!
0%
#151495000000
1!
1%
#151500000000
0!
0%
#151505000000
1!
1%
#151510000000
0!
0%
#151515000000
1!
1%
#151520000000
0!
0%
#151525000000
1!
1%
#151530000000
0!
0%
#151535000000
1!
1%
#151540000000
0!
0%
#151545000000
1!
1%
#151550000000
0!
0%
#151555000000
1!
1%
#151560000000
0!
0%
#151565000000
1!
1%
#151570000000
0!
0%
#151575000000
1!
1%
#151580000000
0!
0%
#151585000000
1!
1%
#151590000000
0!
0%
#151595000000
1!
1%
#151600000000
0!
0%
#151605000000
1!
1%
#151610000000
0!
0%
#151615000000
1!
1%
#151620000000
0!
0%
#151625000000
1!
1%
#151630000000
0!
0%
#151635000000
1!
1%
#151640000000
0!
0%
#151645000000
1!
1%
#151650000000
0!
0%
#151655000000
1!
1%
#151660000000
0!
0%
#151665000000
1!
1%
#151670000000
0!
0%
#151675000000
1!
1%
#151680000000
0!
0%
#151685000000
1!
1%
#151690000000
0!
0%
#151695000000
1!
1%
#151700000000
0!
0%
#151705000000
1!
1%
#151710000000
0!
0%
#151715000000
1!
1%
#151720000000
0!
0%
#151725000000
1!
1%
#151730000000
0!
0%
#151735000000
1!
1%
#151740000000
0!
0%
#151745000000
1!
1%
#151750000000
0!
0%
#151755000000
1!
1%
#151760000000
0!
0%
#151765000000
1!
1%
#151770000000
0!
0%
#151775000000
1!
1%
#151780000000
0!
0%
#151785000000
1!
1%
#151790000000
0!
0%
#151795000000
1!
1%
#151800000000
0!
0%
#151805000000
1!
1%
#151810000000
0!
0%
#151815000000
1!
1%
#151820000000
0!
0%
#151825000000
1!
1%
#151830000000
0!
0%
#151835000000
1!
1%
#151840000000
0!
0%
#151845000000
1!
1%
#151850000000
0!
0%
#151855000000
1!
1%
#151860000000
0!
0%
#151865000000
1!
1%
#151870000000
0!
0%
#151875000000
1!
1%
#151880000000
0!
0%
#151885000000
1!
1%
#151890000000
0!
0%
#151895000000
1!
1%
#151900000000
0!
0%
#151905000000
1!
1%
#151910000000
0!
0%
#151915000000
1!
1%
#151920000000
0!
0%
#151925000000
1!
1%
#151930000000
0!
0%
#151935000000
1!
1%
#151940000000
0!
0%
#151945000000
1!
1%
#151950000000
0!
0%
#151955000000
1!
1%
#151960000000
0!
0%
#151965000000
1!
1%
#151970000000
0!
0%
#151975000000
1!
1%
#151980000000
0!
0%
#151985000000
1!
1%
#151990000000
0!
0%
#151995000000
1!
1%
#152000000000
0!
0%
#152005000000
1!
1%
#152010000000
0!
0%
#152015000000
1!
1%
#152020000000
0!
0%
#152025000000
1!
1%
#152030000000
0!
0%
#152035000000
1!
1%
#152040000000
0!
0%
#152045000000
1!
1%
#152050000000
0!
0%
#152055000000
1!
1%
#152060000000
0!
0%
#152065000000
1!
1%
#152070000000
0!
0%
#152075000000
1!
1%
#152080000000
0!
0%
#152085000000
1!
1%
#152090000000
0!
0%
#152095000000
1!
1%
#152100000000
0!
0%
#152105000000
1!
1%
#152110000000
0!
0%
#152115000000
1!
1%
#152120000000
0!
0%
#152125000000
1!
1%
#152130000000
0!
0%
#152135000000
1!
1%
#152140000000
0!
0%
#152145000000
1!
1%
#152150000000
0!
0%
#152155000000
1!
1%
#152160000000
0!
0%
#152165000000
1!
1%
#152170000000
0!
0%
#152175000000
1!
1%
#152180000000
0!
0%
#152185000000
1!
1%
#152190000000
0!
0%
#152195000000
1!
1%
#152200000000
0!
0%
#152205000000
1!
1%
#152210000000
0!
0%
#152215000000
1!
1%
#152220000000
0!
0%
#152225000000
1!
1%
#152230000000
0!
0%
#152235000000
1!
1%
#152240000000
0!
0%
#152245000000
1!
1%
#152250000000
0!
0%
#152255000000
1!
1%
#152260000000
0!
0%
#152265000000
1!
1%
#152270000000
0!
0%
#152275000000
1!
1%
#152280000000
0!
0%
#152285000000
1!
1%
#152290000000
0!
0%
#152295000000
1!
1%
#152300000000
0!
0%
#152305000000
1!
1%
#152310000000
0!
0%
#152315000000
1!
1%
#152320000000
0!
0%
#152325000000
1!
1%
#152330000000
0!
0%
#152335000000
1!
1%
#152340000000
0!
0%
#152345000000
1!
1%
#152350000000
0!
0%
#152355000000
1!
1%
#152360000000
0!
0%
#152365000000
1!
1%
#152370000000
0!
0%
#152375000000
1!
1%
#152380000000
0!
0%
#152385000000
1!
1%
#152390000000
0!
0%
#152395000000
1!
1%
#152400000000
0!
0%
#152405000000
1!
1%
#152410000000
0!
0%
#152415000000
1!
1%
#152420000000
0!
0%
#152425000000
1!
1%
#152430000000
0!
0%
#152435000000
1!
1%
#152440000000
0!
0%
#152445000000
1!
1%
#152450000000
0!
0%
#152455000000
1!
1%
#152460000000
0!
0%
#152465000000
1!
1%
#152470000000
0!
0%
#152475000000
1!
1%
#152480000000
0!
0%
#152485000000
1!
1%
#152490000000
0!
0%
#152495000000
1!
1%
#152500000000
0!
0%
#152505000000
1!
1%
#152510000000
0!
0%
#152515000000
1!
1%
#152520000000
0!
0%
#152525000000
1!
1%
#152530000000
0!
0%
#152535000000
1!
1%
#152540000000
0!
0%
#152545000000
1!
1%
#152550000000
0!
0%
#152555000000
1!
1%
#152560000000
0!
0%
#152565000000
1!
1%
#152570000000
0!
0%
#152575000000
1!
1%
#152580000000
0!
0%
#152585000000
1!
1%
#152590000000
0!
0%
#152595000000
1!
1%
#152600000000
0!
0%
#152605000000
1!
1%
#152610000000
0!
0%
#152615000000
1!
1%
#152620000000
0!
0%
#152625000000
1!
1%
#152630000000
0!
0%
#152635000000
1!
1%
#152640000000
0!
0%
#152645000000
1!
1%
#152650000000
0!
0%
#152655000000
1!
1%
#152660000000
0!
0%
#152665000000
1!
1%
#152670000000
0!
0%
#152675000000
1!
1%
#152680000000
0!
0%
#152685000000
1!
1%
#152690000000
0!
0%
#152695000000
1!
1%
#152700000000
0!
0%
#152705000000
1!
1%
#152710000000
0!
0%
#152715000000
1!
1%
#152720000000
0!
0%
#152725000000
1!
1%
#152730000000
0!
0%
#152735000000
1!
1%
#152740000000
0!
0%
#152745000000
1!
1%
#152750000000
0!
0%
#152755000000
1!
1%
#152760000000
0!
0%
#152765000000
1!
1%
#152770000000
0!
0%
#152775000000
1!
1%
#152780000000
0!
0%
#152785000000
1!
1%
#152790000000
0!
0%
#152795000000
1!
1%
#152800000000
0!
0%
#152805000000
1!
1%
#152810000000
0!
0%
#152815000000
1!
1%
#152820000000
0!
0%
#152825000000
1!
1%
#152830000000
0!
0%
#152835000000
1!
1%
#152840000000
0!
0%
#152845000000
1!
1%
#152850000000
0!
0%
#152855000000
1!
1%
#152860000000
0!
0%
#152865000000
1!
1%
#152870000000
0!
0%
#152875000000
1!
1%
#152880000000
0!
0%
#152885000000
1!
1%
#152890000000
0!
0%
#152895000000
1!
1%
#152900000000
0!
0%
#152905000000
1!
1%
#152910000000
0!
0%
#152915000000
1!
1%
#152920000000
0!
0%
#152925000000
1!
1%
#152930000000
0!
0%
#152935000000
1!
1%
#152940000000
0!
0%
#152945000000
1!
1%
#152950000000
0!
0%
#152955000000
1!
1%
#152960000000
0!
0%
#152965000000
1!
1%
#152970000000
0!
0%
#152975000000
1!
1%
#152980000000
0!
0%
#152985000000
1!
1%
#152990000000
0!
0%
#152995000000
1!
1%
#153000000000
0!
0%
#153005000000
1!
1%
#153010000000
0!
0%
#153015000000
1!
1%
#153020000000
0!
0%
#153025000000
1!
1%
#153030000000
0!
0%
#153035000000
1!
1%
#153040000000
0!
0%
#153045000000
1!
1%
#153050000000
0!
0%
#153055000000
1!
1%
#153060000000
0!
0%
#153065000000
1!
1%
#153070000000
0!
0%
#153075000000
1!
1%
#153080000000
0!
0%
#153085000000
1!
1%
#153090000000
0!
0%
#153095000000
1!
1%
#153100000000
0!
0%
#153105000000
1!
1%
#153110000000
0!
0%
#153115000000
1!
1%
#153120000000
0!
0%
#153125000000
1!
1%
#153130000000
0!
0%
#153135000000
1!
1%
#153140000000
0!
0%
#153145000000
1!
1%
#153150000000
0!
0%
#153155000000
1!
1%
#153160000000
0!
0%
#153165000000
1!
1%
#153170000000
0!
0%
#153175000000
1!
1%
#153180000000
0!
0%
#153185000000
1!
1%
#153190000000
0!
0%
#153195000000
1!
1%
#153200000000
0!
0%
#153205000000
1!
1%
#153210000000
0!
0%
#153215000000
1!
1%
#153220000000
0!
0%
#153225000000
1!
1%
#153230000000
0!
0%
#153235000000
1!
1%
#153240000000
0!
0%
#153245000000
1!
1%
#153250000000
0!
0%
#153255000000
1!
1%
#153260000000
0!
0%
#153265000000
1!
1%
#153270000000
0!
0%
#153275000000
1!
1%
#153280000000
0!
0%
#153285000000
1!
1%
#153290000000
0!
0%
#153295000000
1!
1%
#153300000000
0!
0%
#153305000000
1!
1%
#153310000000
0!
0%
#153315000000
1!
1%
#153320000000
0!
0%
#153325000000
1!
1%
#153330000000
0!
0%
#153335000000
1!
1%
#153340000000
0!
0%
#153345000000
1!
1%
#153350000000
0!
0%
#153355000000
1!
1%
#153360000000
0!
0%
#153365000000
1!
1%
#153370000000
0!
0%
#153375000000
1!
1%
#153380000000
0!
0%
#153385000000
1!
1%
#153390000000
0!
0%
#153395000000
1!
1%
#153400000000
0!
0%
#153405000000
1!
1%
#153410000000
0!
0%
#153415000000
1!
1%
#153420000000
0!
0%
#153425000000
1!
1%
#153430000000
0!
0%
#153435000000
1!
1%
#153440000000
0!
0%
#153445000000
1!
1%
#153450000000
0!
0%
#153455000000
1!
1%
#153460000000
0!
0%
#153465000000
1!
1%
#153470000000
0!
0%
#153475000000
1!
1%
#153480000000
0!
0%
#153485000000
1!
1%
#153490000000
0!
0%
#153495000000
1!
1%
#153500000000
0!
0%
#153505000000
1!
1%
#153510000000
0!
0%
#153515000000
1!
1%
#153520000000
0!
0%
#153525000000
1!
1%
#153530000000
0!
0%
#153535000000
1!
1%
#153540000000
0!
0%
#153545000000
1!
1%
#153550000000
0!
0%
#153555000000
1!
1%
#153560000000
0!
0%
#153565000000
1!
1%
#153570000000
0!
0%
#153575000000
1!
1%
#153580000000
0!
0%
#153585000000
1!
1%
#153590000000
0!
0%
#153595000000
1!
1%
#153600000000
0!
0%
#153605000000
1!
1%
#153610000000
0!
0%
#153615000000
1!
1%
#153620000000
0!
0%
#153625000000
1!
1%
#153630000000
0!
0%
#153635000000
1!
1%
#153640000000
0!
0%
#153645000000
1!
1%
#153650000000
0!
0%
#153655000000
1!
1%
#153660000000
0!
0%
#153665000000
1!
1%
#153670000000
0!
0%
#153675000000
1!
1%
#153680000000
0!
0%
#153685000000
1!
1%
#153690000000
0!
0%
#153695000000
1!
1%
#153700000000
0!
0%
#153705000000
1!
1%
#153710000000
0!
0%
#153715000000
1!
1%
#153720000000
0!
0%
#153725000000
1!
1%
#153730000000
0!
0%
#153735000000
1!
1%
#153740000000
0!
0%
#153745000000
1!
1%
#153750000000
0!
0%
#153755000000
1!
1%
#153760000000
0!
0%
#153765000000
1!
1%
#153770000000
0!
0%
#153775000000
1!
1%
#153780000000
0!
0%
#153785000000
1!
1%
#153790000000
0!
0%
#153795000000
1!
1%
#153800000000
0!
0%
#153805000000
1!
1%
#153810000000
0!
0%
#153815000000
1!
1%
#153820000000
0!
0%
#153825000000
1!
1%
#153830000000
0!
0%
#153835000000
1!
1%
#153840000000
0!
0%
#153845000000
1!
1%
#153850000000
0!
0%
#153855000000
1!
1%
#153860000000
0!
0%
#153865000000
1!
1%
#153870000000
0!
0%
#153875000000
1!
1%
#153880000000
0!
0%
#153885000000
1!
1%
#153890000000
0!
0%
#153895000000
1!
1%
#153900000000
0!
0%
#153905000000
1!
1%
#153910000000
0!
0%
#153915000000
1!
1%
#153920000000
0!
0%
#153925000000
1!
1%
#153930000000
0!
0%
#153935000000
1!
1%
#153940000000
0!
0%
#153945000000
1!
1%
#153950000000
0!
0%
#153955000000
1!
1%
#153960000000
0!
0%
#153965000000
1!
1%
#153970000000
0!
0%
#153975000000
1!
1%
#153980000000
0!
0%
#153985000000
1!
1%
#153990000000
0!
0%
#153995000000
1!
1%
#154000000000
0!
0%
#154005000000
1!
1%
#154010000000
0!
0%
#154015000000
1!
1%
#154020000000
0!
0%
#154025000000
1!
1%
#154030000000
0!
0%
#154035000000
1!
1%
#154040000000
0!
0%
#154045000000
1!
1%
#154050000000
0!
0%
#154055000000
1!
1%
#154060000000
0!
0%
#154065000000
1!
1%
#154070000000
0!
0%
#154075000000
1!
1%
#154080000000
0!
0%
#154085000000
1!
1%
#154090000000
0!
0%
#154095000000
1!
1%
#154100000000
0!
0%
#154105000000
1!
1%
#154110000000
0!
0%
#154115000000
1!
1%
#154120000000
0!
0%
#154125000000
1!
1%
#154130000000
0!
0%
#154135000000
1!
1%
#154140000000
0!
0%
#154145000000
1!
1%
#154150000000
0!
0%
#154155000000
1!
1%
#154160000000
0!
0%
#154165000000
1!
1%
#154170000000
0!
0%
#154175000000
1!
1%
#154180000000
0!
0%
#154185000000
1!
1%
#154190000000
0!
0%
#154195000000
1!
1%
#154200000000
0!
0%
#154205000000
1!
1%
#154210000000
0!
0%
#154215000000
1!
1%
#154220000000
0!
0%
#154225000000
1!
1%
#154230000000
0!
0%
#154235000000
1!
1%
#154240000000
0!
0%
#154245000000
1!
1%
#154250000000
0!
0%
#154255000000
1!
1%
#154260000000
0!
0%
#154265000000
1!
1%
#154270000000
0!
0%
#154275000000
1!
1%
#154280000000
0!
0%
#154285000000
1!
1%
#154290000000
0!
0%
#154295000000
1!
1%
#154300000000
0!
0%
#154305000000
1!
1%
#154310000000
0!
0%
#154315000000
1!
1%
#154320000000
0!
0%
#154325000000
1!
1%
#154330000000
0!
0%
#154335000000
1!
1%
#154340000000
0!
0%
#154345000000
1!
1%
#154350000000
0!
0%
#154355000000
1!
1%
#154360000000
0!
0%
#154365000000
1!
1%
#154370000000
0!
0%
#154375000000
1!
1%
#154380000000
0!
0%
#154385000000
1!
1%
#154390000000
0!
0%
#154395000000
1!
1%
#154400000000
0!
0%
#154405000000
1!
1%
#154410000000
0!
0%
#154415000000
1!
1%
#154420000000
0!
0%
#154425000000
1!
1%
#154430000000
0!
0%
#154435000000
1!
1%
#154440000000
0!
0%
#154445000000
1!
1%
#154450000000
0!
0%
#154455000000
1!
1%
#154460000000
0!
0%
#154465000000
1!
1%
#154470000000
0!
0%
#154475000000
1!
1%
#154480000000
0!
0%
#154485000000
1!
1%
#154490000000
0!
0%
#154495000000
1!
1%
#154500000000
0!
0%
#154505000000
1!
1%
#154510000000
0!
0%
#154515000000
1!
1%
#154520000000
0!
0%
#154525000000
1!
1%
#154530000000
0!
0%
#154535000000
1!
1%
#154540000000
0!
0%
#154545000000
1!
1%
#154550000000
0!
0%
#154555000000
1!
1%
#154560000000
0!
0%
#154565000000
1!
1%
#154570000000
0!
0%
#154575000000
1!
1%
#154580000000
0!
0%
#154585000000
1!
1%
#154590000000
0!
0%
#154595000000
1!
1%
#154600000000
0!
0%
#154605000000
1!
1%
#154610000000
0!
0%
#154615000000
1!
1%
#154620000000
0!
0%
#154625000000
1!
1%
#154630000000
0!
0%
#154635000000
1!
1%
#154640000000
0!
0%
#154645000000
1!
1%
#154650000000
0!
0%
#154655000000
1!
1%
#154660000000
0!
0%
#154665000000
1!
1%
#154670000000
0!
0%
#154675000000
1!
1%
#154680000000
0!
0%
#154685000000
1!
1%
#154690000000
0!
0%
#154695000000
1!
1%
#154700000000
0!
0%
#154705000000
1!
1%
#154710000000
0!
0%
#154715000000
1!
1%
#154720000000
0!
0%
#154725000000
1!
1%
#154730000000
0!
0%
#154735000000
1!
1%
#154740000000
0!
0%
#154745000000
1!
1%
#154750000000
0!
0%
#154755000000
1!
1%
#154760000000
0!
0%
#154765000000
1!
1%
#154770000000
0!
0%
#154775000000
1!
1%
#154780000000
0!
0%
#154785000000
1!
1%
#154790000000
0!
0%
#154795000000
1!
1%
#154800000000
0!
0%
#154805000000
1!
1%
#154810000000
0!
0%
#154815000000
1!
1%
#154820000000
0!
0%
#154825000000
1!
1%
#154830000000
0!
0%
#154835000000
1!
1%
#154840000000
0!
0%
#154845000000
1!
1%
#154850000000
0!
0%
#154855000000
1!
1%
#154860000000
0!
0%
#154865000000
1!
1%
#154870000000
0!
0%
#154875000000
1!
1%
#154880000000
0!
0%
#154885000000
1!
1%
#154890000000
0!
0%
#154895000000
1!
1%
#154900000000
0!
0%
#154905000000
1!
1%
#154910000000
0!
0%
#154915000000
1!
1%
#154920000000
0!
0%
#154925000000
1!
1%
#154930000000
0!
0%
#154935000000
1!
1%
#154940000000
0!
0%
#154945000000
1!
1%
#154950000000
0!
0%
#154955000000
1!
1%
#154960000000
0!
0%
#154965000000
1!
1%
#154970000000
0!
0%
#154975000000
1!
1%
#154980000000
0!
0%
#154985000000
1!
1%
#154990000000
0!
0%
#154995000000
1!
1%
#155000000000
0!
0%
#155005000000
1!
1%
#155010000000
0!
0%
#155015000000
1!
1%
#155020000000
0!
0%
#155025000000
1!
1%
#155030000000
0!
0%
#155035000000
1!
1%
#155040000000
0!
0%
#155045000000
1!
1%
#155050000000
0!
0%
#155055000000
1!
1%
#155060000000
0!
0%
#155065000000
1!
1%
#155070000000
0!
0%
#155075000000
1!
1%
#155080000000
0!
0%
#155085000000
1!
1%
#155090000000
0!
0%
#155095000000
1!
1%
#155100000000
0!
0%
#155105000000
1!
1%
#155110000000
0!
0%
#155115000000
1!
1%
#155120000000
0!
0%
#155125000000
1!
1%
#155130000000
0!
0%
#155135000000
1!
1%
#155140000000
0!
0%
#155145000000
1!
1%
#155150000000
0!
0%
#155155000000
1!
1%
#155160000000
0!
0%
#155165000000
1!
1%
#155170000000
0!
0%
#155175000000
1!
1%
#155180000000
0!
0%
#155185000000
1!
1%
#155190000000
0!
0%
#155195000000
1!
1%
#155200000000
0!
0%
#155205000000
1!
1%
#155210000000
0!
0%
#155215000000
1!
1%
#155220000000
0!
0%
#155225000000
1!
1%
#155230000000
0!
0%
#155235000000
1!
1%
#155240000000
0!
0%
#155245000000
1!
1%
#155250000000
0!
0%
#155255000000
1!
1%
#155260000000
0!
0%
#155265000000
1!
1%
#155270000000
0!
0%
#155275000000
1!
1%
#155280000000
0!
0%
#155285000000
1!
1%
#155290000000
0!
0%
#155295000000
1!
1%
#155300000000
0!
0%
#155305000000
1!
1%
#155310000000
0!
0%
#155315000000
1!
1%
#155320000000
0!
0%
#155325000000
1!
1%
#155330000000
0!
0%
#155335000000
1!
1%
#155340000000
0!
0%
#155345000000
1!
1%
#155350000000
0!
0%
#155355000000
1!
1%
#155360000000
0!
0%
#155365000000
1!
1%
#155370000000
0!
0%
#155375000000
1!
1%
#155380000000
0!
0%
#155385000000
1!
1%
#155390000000
0!
0%
#155395000000
1!
1%
#155400000000
0!
0%
#155405000000
1!
1%
#155410000000
0!
0%
#155415000000
1!
1%
#155420000000
0!
0%
#155425000000
1!
1%
#155430000000
0!
0%
#155435000000
1!
1%
#155440000000
0!
0%
#155445000000
1!
1%
#155450000000
0!
0%
#155455000000
1!
1%
#155460000000
0!
0%
#155465000000
1!
1%
#155470000000
0!
0%
#155475000000
1!
1%
#155480000000
0!
0%
#155485000000
1!
1%
#155490000000
0!
0%
#155495000000
1!
1%
#155500000000
0!
0%
#155505000000
1!
1%
#155510000000
0!
0%
#155515000000
1!
1%
#155520000000
0!
0%
#155525000000
1!
1%
#155530000000
0!
0%
#155535000000
1!
1%
#155540000000
0!
0%
#155545000000
1!
1%
#155550000000
0!
0%
#155555000000
1!
1%
#155560000000
0!
0%
#155565000000
1!
1%
#155570000000
0!
0%
#155575000000
1!
1%
#155580000000
0!
0%
#155585000000
1!
1%
#155590000000
0!
0%
#155595000000
1!
1%
#155600000000
0!
0%
#155605000000
1!
1%
#155610000000
0!
0%
#155615000000
1!
1%
#155620000000
0!
0%
#155625000000
1!
1%
#155630000000
0!
0%
#155635000000
1!
1%
#155640000000
0!
0%
#155645000000
1!
1%
#155650000000
0!
0%
#155655000000
1!
1%
#155660000000
0!
0%
#155665000000
1!
1%
#155670000000
0!
0%
#155675000000
1!
1%
#155680000000
0!
0%
#155685000000
1!
1%
#155690000000
0!
0%
#155695000000
1!
1%
#155700000000
0!
0%
#155705000000
1!
1%
#155710000000
0!
0%
#155715000000
1!
1%
#155720000000
0!
0%
#155725000000
1!
1%
#155730000000
0!
0%
#155735000000
1!
1%
#155740000000
0!
0%
#155745000000
1!
1%
#155750000000
0!
0%
#155755000000
1!
1%
#155760000000
0!
0%
#155765000000
1!
1%
#155770000000
0!
0%
#155775000000
1!
1%
#155780000000
0!
0%
#155785000000
1!
1%
#155790000000
0!
0%
#155795000000
1!
1%
#155800000000
0!
0%
#155805000000
1!
1%
#155810000000
0!
0%
#155815000000
1!
1%
#155820000000
0!
0%
#155825000000
1!
1%
#155830000000
0!
0%
#155835000000
1!
1%
#155840000000
0!
0%
#155845000000
1!
1%
#155850000000
0!
0%
#155855000000
1!
1%
#155860000000
0!
0%
#155865000000
1!
1%
#155870000000
0!
0%
#155875000000
1!
1%
#155880000000
0!
0%
#155885000000
1!
1%
#155890000000
0!
0%
#155895000000
1!
1%
#155900000000
0!
0%
#155905000000
1!
1%
#155910000000
0!
0%
#155915000000
1!
1%
#155920000000
0!
0%
#155925000000
1!
1%
#155930000000
0!
0%
#155935000000
1!
1%
#155940000000
0!
0%
#155945000000
1!
1%
#155950000000
0!
0%
#155955000000
1!
1%
#155960000000
0!
0%
#155965000000
1!
1%
#155970000000
0!
0%
#155975000000
1!
1%
#155980000000
0!
0%
#155985000000
1!
1%
#155990000000
0!
0%
#155995000000
1!
1%
#156000000000
0!
0%
#156005000000
1!
1%
#156010000000
0!
0%
#156015000000
1!
1%
#156020000000
0!
0%
#156025000000
1!
1%
#156030000000
0!
0%
#156035000000
1!
1%
#156040000000
0!
0%
#156045000000
1!
1%
#156050000000
0!
0%
#156055000000
1!
1%
#156060000000
0!
0%
#156065000000
1!
1%
#156070000000
0!
0%
#156075000000
1!
1%
#156080000000
0!
0%
#156085000000
1!
1%
#156090000000
0!
0%
#156095000000
1!
1%
#156100000000
0!
0%
#156105000000
1!
1%
#156110000000
0!
0%
#156115000000
1!
1%
#156120000000
0!
0%
#156125000000
1!
1%
#156130000000
0!
0%
#156135000000
1!
1%
#156140000000
0!
0%
#156145000000
1!
1%
#156150000000
0!
0%
#156155000000
1!
1%
#156160000000
0!
0%
#156165000000
1!
1%
#156170000000
0!
0%
#156175000000
1!
1%
#156180000000
0!
0%
#156185000000
1!
1%
#156190000000
0!
0%
#156195000000
1!
1%
#156200000000
0!
0%
#156205000000
1!
1%
#156210000000
0!
0%
#156215000000
1!
1%
#156220000000
0!
0%
#156225000000
1!
1%
#156230000000
0!
0%
#156235000000
1!
1%
#156240000000
0!
0%
#156245000000
1!
1%
#156250000000
0!
0%
#156255000000
1!
1%
#156260000000
0!
0%
#156265000000
1!
1%
#156270000000
0!
0%
#156275000000
1!
1%
#156280000000
0!
0%
#156285000000
1!
1%
#156290000000
0!
0%
#156295000000
1!
1%
#156300000000
0!
0%
#156305000000
1!
1%
#156310000000
0!
0%
#156315000000
1!
1%
#156320000000
0!
0%
#156325000000
1!
1%
#156330000000
0!
0%
#156335000000
1!
1%
#156340000000
0!
0%
#156345000000
1!
1%
#156350000000
0!
0%
#156355000000
1!
1%
#156360000000
0!
0%
#156365000000
1!
1%
#156370000000
0!
0%
#156375000000
1!
1%
#156380000000
0!
0%
#156385000000
1!
1%
#156390000000
0!
0%
#156395000000
1!
1%
#156400000000
0!
0%
#156405000000
1!
1%
#156410000000
0!
0%
#156415000000
1!
1%
#156420000000
0!
0%
#156425000000
1!
1%
#156430000000
0!
0%
#156435000000
1!
1%
#156440000000
0!
0%
#156445000000
1!
1%
#156450000000
0!
0%
#156455000000
1!
1%
#156460000000
0!
0%
#156465000000
1!
1%
#156470000000
0!
0%
#156475000000
1!
1%
#156480000000
0!
0%
#156485000000
1!
1%
#156490000000
0!
0%
#156495000000
1!
1%
#156500000000
0!
0%
#156505000000
1!
1%
#156510000000
0!
0%
#156515000000
1!
1%
#156520000000
0!
0%
#156525000000
1!
1%
#156530000000
0!
0%
#156535000000
1!
1%
#156540000000
0!
0%
#156545000000
1!
1%
#156550000000
0!
0%
#156555000000
1!
1%
#156560000000
0!
0%
#156565000000
1!
1%
#156570000000
0!
0%
#156575000000
1!
1%
#156580000000
0!
0%
#156585000000
1!
1%
#156590000000
0!
0%
#156595000000
1!
1%
#156600000000
0!
0%
#156605000000
1!
1%
#156610000000
0!
0%
#156615000000
1!
1%
#156620000000
0!
0%
#156625000000
1!
1%
#156630000000
0!
0%
#156635000000
1!
1%
#156640000000
0!
0%
#156645000000
1!
1%
#156650000000
0!
0%
#156655000000
1!
1%
#156660000000
0!
0%
#156665000000
1!
1%
#156670000000
0!
0%
#156675000000
1!
1%
#156680000000
0!
0%
#156685000000
1!
1%
#156690000000
0!
0%
#156695000000
1!
1%
#156700000000
0!
0%
#156705000000
1!
1%
#156710000000
0!
0%
#156715000000
1!
1%
#156720000000
0!
0%
#156725000000
1!
1%
#156730000000
0!
0%
#156735000000
1!
1%
#156740000000
0!
0%
#156745000000
1!
1%
#156750000000
0!
0%
#156755000000
1!
1%
#156760000000
0!
0%
#156765000000
1!
1%
#156770000000
0!
0%
#156775000000
1!
1%
#156780000000
0!
0%
#156785000000
1!
1%
#156790000000
0!
0%
#156795000000
1!
1%
#156800000000
0!
0%
#156805000000
1!
1%
#156810000000
0!
0%
#156815000000
1!
1%
#156820000000
0!
0%
#156825000000
1!
1%
#156830000000
0!
0%
#156835000000
1!
1%
#156840000000
0!
0%
#156845000000
1!
1%
#156850000000
0!
0%
#156855000000
1!
1%
#156860000000
0!
0%
#156865000000
1!
1%
#156870000000
0!
0%
#156875000000
1!
1%
#156880000000
0!
0%
#156885000000
1!
1%
#156890000000
0!
0%
#156895000000
1!
1%
#156900000000
0!
0%
#156905000000
1!
1%
#156910000000
0!
0%
#156915000000
1!
1%
#156920000000
0!
0%
#156925000000
1!
1%
#156930000000
0!
0%
#156935000000
1!
1%
#156940000000
0!
0%
#156945000000
1!
1%
#156950000000
0!
0%
#156955000000
1!
1%
#156960000000
0!
0%
#156965000000
1!
1%
#156970000000
0!
0%
#156975000000
1!
1%
#156980000000
0!
0%
#156985000000
1!
1%
#156990000000
0!
0%
#156995000000
1!
1%
#157000000000
0!
0%
#157005000000
1!
1%
#157010000000
0!
0%
#157015000000
1!
1%
#157020000000
0!
0%
#157025000000
1!
1%
#157030000000
0!
0%
#157035000000
1!
1%
#157040000000
0!
0%
#157045000000
1!
1%
#157050000000
0!
0%
#157055000000
1!
1%
#157060000000
0!
0%
#157065000000
1!
1%
#157070000000
0!
0%
#157075000000
1!
1%
#157080000000
0!
0%
#157085000000
1!
1%
#157090000000
0!
0%
#157095000000
1!
1%
#157100000000
0!
0%
#157105000000
1!
1%
#157110000000
0!
0%
#157115000000
1!
1%
#157120000000
0!
0%
#157125000000
1!
1%
#157130000000
0!
0%
#157135000000
1!
1%
#157140000000
0!
0%
#157145000000
1!
1%
#157150000000
0!
0%
#157155000000
1!
1%
#157160000000
0!
0%
#157165000000
1!
1%
#157170000000
0!
0%
#157175000000
1!
1%
#157180000000
0!
0%
#157185000000
1!
1%
#157190000000
0!
0%
#157195000000
1!
1%
#157200000000
0!
0%
#157205000000
1!
1%
#157210000000
0!
0%
#157215000000
1!
1%
#157220000000
0!
0%
#157225000000
1!
1%
#157230000000
0!
0%
#157235000000
1!
1%
#157240000000
0!
0%
#157245000000
1!
1%
#157250000000
0!
0%
#157255000000
1!
1%
#157260000000
0!
0%
#157265000000
1!
1%
#157270000000
0!
0%
#157275000000
1!
1%
#157280000000
0!
0%
#157285000000
1!
1%
#157290000000
0!
0%
#157295000000
1!
1%
#157300000000
0!
0%
#157305000000
1!
1%
#157310000000
0!
0%
#157315000000
1!
1%
#157320000000
0!
0%
#157325000000
1!
1%
#157330000000
0!
0%
#157335000000
1!
1%
#157340000000
0!
0%
#157345000000
1!
1%
#157350000000
0!
0%
#157355000000
1!
1%
#157360000000
0!
0%
#157365000000
1!
1%
#157370000000
0!
0%
#157375000000
1!
1%
#157380000000
0!
0%
#157385000000
1!
1%
#157390000000
0!
0%
#157395000000
1!
1%
#157400000000
0!
0%
#157405000000
1!
1%
#157410000000
0!
0%
#157415000000
1!
1%
#157420000000
0!
0%
#157425000000
1!
1%
#157430000000
0!
0%
#157435000000
1!
1%
#157440000000
0!
0%
#157445000000
1!
1%
#157450000000
0!
0%
#157455000000
1!
1%
#157460000000
0!
0%
#157465000000
1!
1%
#157470000000
0!
0%
#157475000000
1!
1%
#157480000000
0!
0%
#157485000000
1!
1%
#157490000000
0!
0%
#157495000000
1!
1%
#157500000000
0!
0%
#157505000000
1!
1%
#157510000000
0!
0%
#157515000000
1!
1%
#157520000000
0!
0%
#157525000000
1!
1%
#157530000000
0!
0%
#157535000000
1!
1%
#157540000000
0!
0%
#157545000000
1!
1%
#157550000000
0!
0%
#157555000000
1!
1%
#157560000000
0!
0%
#157565000000
1!
1%
#157570000000
0!
0%
#157575000000
1!
1%
#157580000000
0!
0%
#157585000000
1!
1%
#157590000000
0!
0%
#157595000000
1!
1%
#157600000000
0!
0%
#157605000000
1!
1%
#157610000000
0!
0%
#157615000000
1!
1%
#157620000000
0!
0%
#157625000000
1!
1%
#157630000000
0!
0%
#157635000000
1!
1%
#157640000000
0!
0%
#157645000000
1!
1%
#157650000000
0!
0%
#157655000000
1!
1%
#157660000000
0!
0%
#157665000000
1!
1%
#157670000000
0!
0%
#157675000000
1!
1%
#157680000000
0!
0%
#157685000000
1!
1%
#157690000000
0!
0%
#157695000000
1!
1%
#157700000000
0!
0%
#157705000000
1!
1%
#157710000000
0!
0%
#157715000000
1!
1%
#157720000000
0!
0%
#157725000000
1!
1%
#157730000000
0!
0%
#157735000000
1!
1%
#157740000000
0!
0%
#157745000000
1!
1%
#157750000000
0!
0%
#157755000000
1!
1%
#157760000000
0!
0%
#157765000000
1!
1%
#157770000000
0!
0%
#157775000000
1!
1%
#157780000000
0!
0%
#157785000000
1!
1%
#157790000000
0!
0%
#157795000000
1!
1%
#157800000000
0!
0%
#157805000000
1!
1%
#157810000000
0!
0%
#157815000000
1!
1%
#157820000000
0!
0%
#157825000000
1!
1%
#157830000000
0!
0%
#157835000000
1!
1%
#157840000000
0!
0%
#157845000000
1!
1%
#157850000000
0!
0%
#157855000000
1!
1%
#157860000000
0!
0%
#157865000000
1!
1%
#157870000000
0!
0%
#157875000000
1!
1%
#157880000000
0!
0%
#157885000000
1!
1%
#157890000000
0!
0%
#157895000000
1!
1%
#157900000000
0!
0%
#157905000000
1!
1%
#157910000000
0!
0%
#157915000000
1!
1%
#157920000000
0!
0%
#157925000000
1!
1%
#157930000000
0!
0%
#157935000000
1!
1%
#157940000000
0!
0%
#157945000000
1!
1%
#157950000000
0!
0%
#157955000000
1!
1%
#157960000000
0!
0%
#157965000000
1!
1%
#157970000000
0!
0%
#157975000000
1!
1%
#157980000000
0!
0%
#157985000000
1!
1%
#157990000000
0!
0%
#157995000000
1!
1%
#158000000000
0!
0%
#158005000000
1!
1%
#158010000000
0!
0%
#158015000000
1!
1%
#158020000000
0!
0%
#158025000000
1!
1%
#158030000000
0!
0%
#158035000000
1!
1%
#158040000000
0!
0%
#158045000000
1!
1%
#158050000000
0!
0%
#158055000000
1!
1%
#158060000000
0!
0%
#158065000000
1!
1%
#158070000000
0!
0%
#158075000000
1!
1%
#158080000000
0!
0%
#158085000000
1!
1%
#158090000000
0!
0%
#158095000000
1!
1%
#158100000000
0!
0%
#158105000000
1!
1%
#158110000000
0!
0%
#158115000000
1!
1%
#158120000000
0!
0%
#158125000000
1!
1%
#158130000000
0!
0%
#158135000000
1!
1%
#158140000000
0!
0%
#158145000000
1!
1%
#158150000000
0!
0%
#158155000000
1!
1%
#158160000000
0!
0%
#158165000000
1!
1%
#158170000000
0!
0%
#158175000000
1!
1%
#158180000000
0!
0%
#158185000000
1!
1%
#158190000000
0!
0%
#158195000000
1!
1%
#158200000000
0!
0%
#158205000000
1!
1%
#158210000000
0!
0%
#158215000000
1!
1%
#158220000000
0!
0%
#158225000000
1!
1%
#158230000000
0!
0%
#158235000000
1!
1%
#158240000000
0!
0%
#158245000000
1!
1%
#158250000000
0!
0%
#158255000000
1!
1%
#158260000000
0!
0%
#158265000000
1!
1%
#158270000000
0!
0%
#158275000000
1!
1%
#158280000000
0!
0%
#158285000000
1!
1%
#158290000000
0!
0%
#158295000000
1!
1%
#158300000000
0!
0%
#158305000000
1!
1%
#158310000000
0!
0%
#158315000000
1!
1%
#158320000000
0!
0%
#158325000000
1!
1%
#158330000000
0!
0%
#158335000000
1!
1%
#158340000000
0!
0%
#158345000000
1!
1%
#158350000000
0!
0%
#158355000000
1!
1%
#158360000000
0!
0%
#158365000000
1!
1%
#158370000000
0!
0%
#158375000000
1!
1%
#158380000000
0!
0%
#158385000000
1!
1%
#158390000000
0!
0%
#158395000000
1!
1%
#158400000000
0!
0%
#158405000000
1!
1%
#158410000000
0!
0%
#158415000000
1!
1%
#158420000000
0!
0%
#158425000000
1!
1%
#158430000000
0!
0%
#158435000000
1!
1%
#158440000000
0!
0%
#158445000000
1!
1%
#158450000000
0!
0%
#158455000000
1!
1%
#158460000000
0!
0%
#158465000000
1!
1%
#158470000000
0!
0%
#158475000000
1!
1%
#158480000000
0!
0%
#158485000000
1!
1%
#158490000000
0!
0%
#158495000000
1!
1%
#158500000000
0!
0%
#158505000000
1!
1%
#158510000000
0!
0%
#158515000000
1!
1%
#158520000000
0!
0%
#158525000000
1!
1%
#158530000000
0!
0%
#158535000000
1!
1%
#158540000000
0!
0%
#158545000000
1!
1%
#158550000000
0!
0%
#158555000000
1!
1%
#158560000000
0!
0%
#158565000000
1!
1%
#158570000000
0!
0%
#158575000000
1!
1%
#158580000000
0!
0%
#158585000000
1!
1%
#158590000000
0!
0%
#158595000000
1!
1%
#158600000000
0!
0%
#158605000000
1!
1%
#158610000000
0!
0%
#158615000000
1!
1%
#158620000000
0!
0%
#158625000000
1!
1%
#158630000000
0!
0%
#158635000000
1!
1%
#158640000000
0!
0%
#158645000000
1!
1%
#158650000000
0!
0%
#158655000000
1!
1%
#158660000000
0!
0%
#158665000000
1!
1%
#158670000000
0!
0%
#158675000000
1!
1%
#158680000000
0!
0%
#158685000000
1!
1%
#158690000000
0!
0%
#158695000000
1!
1%
#158700000000
0!
0%
#158705000000
1!
1%
#158710000000
0!
0%
#158715000000
1!
1%
#158720000000
0!
0%
#158725000000
1!
1%
#158730000000
0!
0%
#158735000000
1!
1%
#158740000000
0!
0%
#158745000000
1!
1%
#158750000000
0!
0%
#158755000000
1!
1%
#158760000000
0!
0%
#158765000000
1!
1%
#158770000000
0!
0%
#158775000000
1!
1%
#158780000000
0!
0%
#158785000000
1!
1%
#158790000000
0!
0%
#158795000000
1!
1%
#158800000000
0!
0%
#158805000000
1!
1%
#158810000000
0!
0%
#158815000000
1!
1%
#158820000000
0!
0%
#158825000000
1!
1%
#158830000000
0!
0%
#158835000000
1!
1%
#158840000000
0!
0%
#158845000000
1!
1%
#158850000000
0!
0%
#158855000000
1!
1%
#158860000000
0!
0%
#158865000000
1!
1%
#158870000000
0!
0%
#158875000000
1!
1%
#158880000000
0!
0%
#158885000000
1!
1%
#158890000000
0!
0%
#158895000000
1!
1%
#158900000000
0!
0%
#158905000000
1!
1%
#158910000000
0!
0%
#158915000000
1!
1%
#158920000000
0!
0%
#158925000000
1!
1%
#158930000000
0!
0%
#158935000000
1!
1%
#158940000000
0!
0%
#158945000000
1!
1%
#158950000000
0!
0%
#158955000000
1!
1%
#158960000000
0!
0%
#158965000000
1!
1%
#158970000000
0!
0%
#158975000000
1!
1%
#158980000000
0!
0%
#158985000000
1!
1%
#158990000000
0!
0%
#158995000000
1!
1%
#159000000000
0!
0%
#159005000000
1!
1%
#159010000000
0!
0%
#159015000000
1!
1%
#159020000000
0!
0%
#159025000000
1!
1%
#159030000000
0!
0%
#159035000000
1!
1%
#159040000000
0!
0%
#159045000000
1!
1%
#159050000000
0!
0%
#159055000000
1!
1%
#159060000000
0!
0%
#159065000000
1!
1%
#159070000000
0!
0%
#159075000000
1!
1%
#159080000000
0!
0%
#159085000000
1!
1%
#159090000000
0!
0%
#159095000000
1!
1%
#159100000000
0!
0%
#159105000000
1!
1%
#159110000000
0!
0%
#159115000000
1!
1%
#159120000000
0!
0%
#159125000000
1!
1%
#159130000000
0!
0%
#159135000000
1!
1%
#159140000000
0!
0%
#159145000000
1!
1%
#159150000000
0!
0%
#159155000000
1!
1%
#159160000000
0!
0%
#159165000000
1!
1%
#159170000000
0!
0%
#159175000000
1!
1%
#159180000000
0!
0%
#159185000000
1!
1%
#159190000000
0!
0%
#159195000000
1!
1%
#159200000000
0!
0%
#159205000000
1!
1%
#159210000000
0!
0%
#159215000000
1!
1%
#159220000000
0!
0%
#159225000000
1!
1%
#159230000000
0!
0%
#159235000000
1!
1%
#159240000000
0!
0%
#159245000000
1!
1%
#159250000000
0!
0%
#159255000000
1!
1%
#159260000000
0!
0%
#159265000000
1!
1%
#159270000000
0!
0%
#159275000000
1!
1%
#159280000000
0!
0%
#159285000000
1!
1%
#159290000000
0!
0%
#159295000000
1!
1%
#159300000000
0!
0%
#159305000000
1!
1%
#159310000000
0!
0%
#159315000000
1!
1%
#159320000000
0!
0%
#159325000000
1!
1%
#159330000000
0!
0%
#159335000000
1!
1%
#159340000000
0!
0%
#159345000000
1!
1%
#159350000000
0!
0%
#159355000000
1!
1%
#159360000000
0!
0%
#159365000000
1!
1%
#159370000000
0!
0%
#159375000000
1!
1%
#159380000000
0!
0%
#159385000000
1!
1%
#159390000000
0!
0%
#159395000000
1!
1%
#159400000000
0!
0%
#159405000000
1!
1%
#159410000000
0!
0%
#159415000000
1!
1%
#159420000000
0!
0%
#159425000000
1!
1%
#159430000000
0!
0%
#159435000000
1!
1%
#159440000000
0!
0%
#159445000000
1!
1%
#159450000000
0!
0%
#159455000000
1!
1%
#159460000000
0!
0%
#159465000000
1!
1%
#159470000000
0!
0%
#159475000000
1!
1%
#159480000000
0!
0%
#159485000000
1!
1%
#159490000000
0!
0%
#159495000000
1!
1%
#159500000000
0!
0%
#159505000000
1!
1%
#159510000000
0!
0%
#159515000000
1!
1%
#159520000000
0!
0%
#159525000000
1!
1%
#159530000000
0!
0%
#159535000000
1!
1%
#159540000000
0!
0%
#159545000000
1!
1%
#159550000000
0!
0%
#159555000000
1!
1%
#159560000000
0!
0%
#159565000000
1!
1%
#159570000000
0!
0%
#159575000000
1!
1%
#159580000000
0!
0%
#159585000000
1!
1%
#159590000000
0!
0%
#159595000000
1!
1%
#159600000000
0!
0%
#159605000000
1!
1%
#159610000000
0!
0%
#159615000000
1!
1%
#159620000000
0!
0%
#159625000000
1!
1%
#159630000000
0!
0%
#159635000000
1!
1%
#159640000000
0!
0%
#159645000000
1!
1%
#159650000000
0!
0%
#159655000000
1!
1%
#159660000000
0!
0%
#159665000000
1!
1%
#159670000000
0!
0%
#159675000000
1!
1%
#159680000000
0!
0%
#159685000000
1!
1%
#159690000000
0!
0%
#159695000000
1!
1%
#159700000000
0!
0%
#159705000000
1!
1%
#159710000000
0!
0%
#159715000000
1!
1%
#159720000000
0!
0%
#159725000000
1!
1%
#159730000000
0!
0%
#159735000000
1!
1%
#159740000000
0!
0%
#159745000000
1!
1%
#159750000000
0!
0%
#159755000000
1!
1%
#159760000000
0!
0%
#159765000000
1!
1%
#159770000000
0!
0%
#159775000000
1!
1%
#159780000000
0!
0%
#159785000000
1!
1%
#159790000000
0!
0%
#159795000000
1!
1%
#159800000000
0!
0%
#159805000000
1!
1%
#159810000000
0!
0%
#159815000000
1!
1%
#159820000000
0!
0%
#159825000000
1!
1%
#159830000000
0!
0%
#159835000000
1!
1%
#159840000000
0!
0%
#159845000000
1!
1%
#159850000000
0!
0%
#159855000000
1!
1%
#159860000000
0!
0%
#159865000000
1!
1%
#159870000000
0!
0%
#159875000000
1!
1%
#159880000000
0!
0%
#159885000000
1!
1%
#159890000000
0!
0%
#159895000000
1!
1%
#159900000000
0!
0%
#159905000000
1!
1%
#159910000000
0!
0%
#159915000000
1!
1%
#159920000000
0!
0%
#159925000000
1!
1%
#159930000000
0!
0%
#159935000000
1!
1%
#159940000000
0!
0%
#159945000000
1!
1%
#159950000000
0!
0%
#159955000000
1!
1%
#159960000000
0!
0%
#159965000000
1!
1%
#159970000000
0!
0%
#159975000000
1!
1%
#159980000000
0!
0%
#159985000000
1!
1%
#159990000000
0!
0%
#159995000000
1!
1%
#160000000000
0!
0%
#160005000000
1!
1%
#160010000000
0!
0%
#160015000000
1!
1%
#160020000000
0!
0%
#160025000000
1!
1%
#160030000000
0!
0%
#160035000000
1!
1%
#160040000000
0!
0%
#160045000000
1!
1%
#160050000000
0!
0%
#160055000000
1!
1%
#160060000000
0!
0%
#160065000000
1!
1%
#160070000000
0!
0%
#160075000000
1!
1%
#160080000000
0!
0%
#160085000000
1!
1%
#160090000000
0!
0%
#160095000000
1!
1%
#160100000000
0!
0%
#160105000000
1!
1%
#160110000000
0!
0%
#160115000000
1!
1%
#160120000000
0!
0%
#160125000000
1!
1%
#160130000000
0!
0%
#160135000000
1!
1%
#160140000000
0!
0%
#160145000000
1!
1%
#160150000000
0!
0%
#160155000000
1!
1%
#160160000000
0!
0%
#160165000000
1!
1%
#160170000000
0!
0%
#160175000000
1!
1%
#160180000000
0!
0%
#160185000000
1!
1%
#160190000000
0!
0%
#160195000000
1!
1%
#160200000000
0!
0%
#160205000000
1!
1%
#160210000000
0!
0%
#160215000000
1!
1%
#160220000000
0!
0%
#160225000000
1!
1%
#160230000000
0!
0%
#160235000000
1!
1%
#160240000000
0!
0%
#160245000000
1!
1%
#160250000000
0!
0%
#160255000000
1!
1%
#160260000000
0!
0%
#160265000000
1!
1%
#160270000000
0!
0%
#160275000000
1!
1%
#160280000000
0!
0%
#160285000000
1!
1%
#160290000000
0!
0%
#160295000000
1!
1%
#160300000000
0!
0%
#160305000000
1!
1%
#160310000000
0!
0%
#160315000000
1!
1%
#160320000000
0!
0%
#160325000000
1!
1%
#160330000000
0!
0%
#160335000000
1!
1%
#160340000000
0!
0%
#160345000000
1!
1%
#160350000000
0!
0%
#160355000000
1!
1%
#160360000000
0!
0%
#160365000000
1!
1%
#160370000000
0!
0%
#160375000000
1!
1%
#160380000000
0!
0%
#160385000000
1!
1%
#160390000000
0!
0%
#160395000000
1!
1%
#160400000000
0!
0%
#160405000000
1!
1%
#160410000000
0!
0%
#160415000000
1!
1%
#160420000000
0!
0%
#160425000000
1!
1%
#160430000000
0!
0%
#160435000000
1!
1%
#160440000000
0!
0%
#160445000000
1!
1%
#160450000000
0!
0%
#160455000000
1!
1%
#160460000000
0!
0%
#160465000000
1!
1%
#160470000000
0!
0%
#160475000000
1!
1%
#160480000000
0!
0%
#160485000000
1!
1%
#160490000000
0!
0%
#160495000000
1!
1%
#160500000000
0!
0%
#160505000000
1!
1%
#160510000000
0!
0%
#160515000000
1!
1%
#160520000000
0!
0%
#160525000000
1!
1%
#160530000000
0!
0%
#160535000000
1!
1%
#160540000000
0!
0%
#160545000000
1!
1%
#160550000000
0!
0%
#160555000000
1!
1%
#160560000000
0!
0%
#160565000000
1!
1%
#160570000000
0!
0%
#160575000000
1!
1%
#160580000000
0!
0%
#160585000000
1!
1%
#160590000000
0!
0%
#160595000000
1!
1%
#160600000000
0!
0%
#160605000000
1!
1%
#160610000000
0!
0%
#160615000000
1!
1%
#160620000000
0!
0%
#160625000000
1!
1%
#160630000000
0!
0%
#160635000000
1!
1%
#160640000000
0!
0%
#160645000000
1!
1%
#160650000000
0!
0%
#160655000000
1!
1%
#160660000000
0!
0%
#160665000000
1!
1%
#160670000000
0!
0%
#160675000000
1!
1%
#160680000000
0!
0%
#160685000000
1!
1%
#160690000000
0!
0%
#160695000000
1!
1%
#160700000000
0!
0%
#160705000000
1!
1%
#160710000000
0!
0%
#160715000000
1!
1%
#160720000000
0!
0%
#160725000000
1!
1%
#160730000000
0!
0%
#160735000000
1!
1%
#160740000000
0!
0%
#160745000000
1!
1%
#160750000000
0!
0%
#160755000000
1!
1%
#160760000000
0!
0%
#160765000000
1!
1%
#160770000000
0!
0%
#160775000000
1!
1%
#160780000000
0!
0%
#160785000000
1!
1%
#160790000000
0!
0%
#160795000000
1!
1%
#160800000000
0!
0%
#160805000000
1!
1%
#160810000000
0!
0%
#160815000000
1!
1%
#160820000000
0!
0%
#160825000000
1!
1%
#160830000000
0!
0%
#160835000000
1!
1%
#160840000000
0!
0%
#160845000000
1!
1%
#160850000000
0!
0%
#160855000000
1!
1%
#160860000000
0!
0%
#160865000000
1!
1%
#160870000000
0!
0%
#160875000000
1!
1%
#160880000000
0!
0%
#160885000000
1!
1%
#160890000000
0!
0%
#160895000000
1!
1%
#160900000000
0!
0%
#160905000000
1!
1%
#160910000000
0!
0%
#160915000000
1!
1%
#160920000000
0!
0%
#160925000000
1!
1%
#160930000000
0!
0%
#160935000000
1!
1%
#160940000000
0!
0%
#160945000000
1!
1%
#160950000000
0!
0%
#160955000000
1!
1%
#160960000000
0!
0%
#160965000000
1!
1%
#160970000000
0!
0%
#160975000000
1!
1%
#160980000000
0!
0%
#160985000000
1!
1%
#160990000000
0!
0%
#160995000000
1!
1%
#161000000000
0!
0%
#161005000000
1!
1%
#161010000000
0!
0%
#161015000000
1!
1%
#161020000000
0!
0%
#161025000000
1!
1%
#161030000000
0!
0%
#161035000000
1!
1%
#161040000000
0!
0%
#161045000000
1!
1%
#161050000000
0!
0%
#161055000000
1!
1%
#161060000000
0!
0%
#161065000000
1!
1%
#161070000000
0!
0%
#161075000000
1!
1%
#161080000000
0!
0%
#161085000000
1!
1%
#161090000000
0!
0%
#161095000000
1!
1%
#161100000000
0!
0%
#161105000000
1!
1%
#161110000000
0!
0%
#161115000000
1!
1%
#161120000000
0!
0%
#161125000000
1!
1%
#161130000000
0!
0%
#161135000000
1!
1%
#161140000000
0!
0%
#161145000000
1!
1%
#161150000000
0!
0%
#161155000000
1!
1%
#161160000000
0!
0%
#161165000000
1!
1%
#161170000000
0!
0%
#161175000000
1!
1%
#161180000000
0!
0%
#161185000000
1!
1%
#161190000000
0!
0%
#161195000000
1!
1%
#161200000000
0!
0%
#161205000000
1!
1%
#161210000000
0!
0%
#161215000000
1!
1%
#161220000000
0!
0%
#161225000000
1!
1%
#161230000000
0!
0%
#161235000000
1!
1%
#161240000000
0!
0%
#161245000000
1!
1%
#161250000000
0!
0%
#161255000000
1!
1%
#161260000000
0!
0%
#161265000000
1!
1%
#161270000000
0!
0%
#161275000000
1!
1%
#161280000000
0!
0%
#161285000000
1!
1%
#161290000000
0!
0%
#161295000000
1!
1%
#161300000000
0!
0%
#161305000000
1!
1%
#161310000000
0!
0%
#161315000000
1!
1%
#161320000000
0!
0%
#161325000000
1!
1%
#161330000000
0!
0%
#161335000000
1!
1%
#161340000000
0!
0%
#161345000000
1!
1%
#161350000000
0!
0%
#161355000000
1!
1%
#161360000000
0!
0%
#161365000000
1!
1%
#161370000000
0!
0%
#161375000000
1!
1%
#161380000000
0!
0%
#161385000000
1!
1%
#161390000000
0!
0%
#161395000000
1!
1%
#161400000000
0!
0%
#161405000000
1!
1%
#161410000000
0!
0%
#161415000000
1!
1%
#161420000000
0!
0%
#161425000000
1!
1%
#161430000000
0!
0%
#161435000000
1!
1%
#161440000000
0!
0%
#161445000000
1!
1%
#161450000000
0!
0%
#161455000000
1!
1%
#161460000000
0!
0%
#161465000000
1!
1%
#161470000000
0!
0%
#161475000000
1!
1%
#161480000000
0!
0%
#161485000000
1!
1%
#161490000000
0!
0%
#161495000000
1!
1%
#161500000000
0!
0%
#161505000000
1!
1%
#161510000000
0!
0%
#161515000000
1!
1%
#161520000000
0!
0%
#161525000000
1!
1%
#161530000000
0!
0%
#161535000000
1!
1%
#161540000000
0!
0%
#161545000000
1!
1%
#161550000000
0!
0%
#161555000000
1!
1%
#161560000000
0!
0%
#161565000000
1!
1%
#161570000000
0!
0%
#161575000000
1!
1%
#161580000000
0!
0%
#161585000000
1!
1%
#161590000000
0!
0%
#161595000000
1!
1%
#161600000000
0!
0%
#161605000000
1!
1%
#161610000000
0!
0%
#161615000000
1!
1%
#161620000000
0!
0%
#161625000000
1!
1%
#161630000000
0!
0%
#161635000000
1!
1%
#161640000000
0!
0%
#161645000000
1!
1%
#161650000000
0!
0%
#161655000000
1!
1%
#161660000000
0!
0%
#161665000000
1!
1%
#161670000000
0!
0%
#161675000000
1!
1%
#161680000000
0!
0%
#161685000000
1!
1%
#161690000000
0!
0%
#161695000000
1!
1%
#161700000000
0!
0%
#161705000000
1!
1%
#161710000000
0!
0%
#161715000000
1!
1%
#161720000000
0!
0%
#161725000000
1!
1%
#161730000000
0!
0%
#161735000000
1!
1%
#161740000000
0!
0%
#161745000000
1!
1%
#161750000000
0!
0%
#161755000000
1!
1%
#161760000000
0!
0%
#161765000000
1!
1%
#161770000000
0!
0%
#161775000000
1!
1%
#161780000000
0!
0%
#161785000000
1!
1%
#161790000000
0!
0%
#161795000000
1!
1%
#161800000000
0!
0%
#161805000000
1!
1%
#161810000000
0!
0%
#161815000000
1!
1%
#161820000000
0!
0%
#161825000000
1!
1%
#161830000000
0!
0%
#161835000000
1!
1%
#161840000000
0!
0%
#161845000000
1!
1%
#161850000000
0!
0%
#161855000000
1!
1%
#161860000000
0!
0%
#161865000000
1!
1%
#161870000000
0!
0%
#161875000000
1!
1%
#161880000000
0!
0%
#161885000000
1!
1%
#161890000000
0!
0%
#161895000000
1!
1%
#161900000000
0!
0%
#161905000000
1!
1%
#161910000000
0!
0%
#161915000000
1!
1%
#161920000000
0!
0%
#161925000000
1!
1%
#161930000000
0!
0%
#161935000000
1!
1%
#161940000000
0!
0%
#161945000000
1!
1%
#161950000000
0!
0%
#161955000000
1!
1%
#161960000000
0!
0%
#161965000000
1!
1%
#161970000000
0!
0%
#161975000000
1!
1%
#161980000000
0!
0%
#161985000000
1!
1%
#161990000000
0!
0%
#161995000000
1!
1%
#162000000000
0!
0%
#162005000000
1!
1%
#162010000000
0!
0%
#162015000000
1!
1%
#162020000000
0!
0%
#162025000000
1!
1%
#162030000000
0!
0%
#162035000000
1!
1%
#162040000000
0!
0%
#162045000000
1!
1%
#162050000000
0!
0%
#162055000000
1!
1%
#162060000000
0!
0%
#162065000000
1!
1%
#162070000000
0!
0%
#162075000000
1!
1%
#162080000000
0!
0%
#162085000000
1!
1%
#162090000000
0!
0%
#162095000000
1!
1%
#162100000000
0!
0%
#162105000000
1!
1%
#162110000000
0!
0%
#162115000000
1!
1%
#162120000000
0!
0%
#162125000000
1!
1%
#162130000000
0!
0%
#162135000000
1!
1%
#162140000000
0!
0%
#162145000000
1!
1%
#162150000000
0!
0%
#162155000000
1!
1%
#162160000000
0!
0%
#162165000000
1!
1%
#162170000000
0!
0%
#162175000000
1!
1%
#162180000000
0!
0%
#162185000000
1!
1%
#162190000000
0!
0%
#162195000000
1!
1%
#162200000000
0!
0%
#162205000000
1!
1%
#162210000000
0!
0%
#162215000000
1!
1%
#162220000000
0!
0%
#162225000000
1!
1%
#162230000000
0!
0%
#162235000000
1!
1%
#162240000000
0!
0%
#162245000000
1!
1%
#162250000000
0!
0%
#162255000000
1!
1%
#162260000000
0!
0%
#162265000000
1!
1%
#162270000000
0!
0%
#162275000000
1!
1%
#162280000000
0!
0%
#162285000000
1!
1%
#162290000000
0!
0%
#162295000000
1!
1%
#162300000000
0!
0%
#162305000000
1!
1%
#162310000000
0!
0%
#162315000000
1!
1%
#162320000000
0!
0%
#162325000000
1!
1%
#162330000000
0!
0%
#162335000000
1!
1%
#162340000000
0!
0%
#162345000000
1!
1%
#162350000000
0!
0%
#162355000000
1!
1%
#162360000000
0!
0%
#162365000000
1!
1%
#162370000000
0!
0%
#162375000000
1!
1%
#162380000000
0!
0%
#162385000000
1!
1%
#162390000000
0!
0%
#162395000000
1!
1%
#162400000000
0!
0%
#162405000000
1!
1%
#162410000000
0!
0%
#162415000000
1!
1%
#162420000000
0!
0%
#162425000000
1!
1%
#162430000000
0!
0%
#162435000000
1!
1%
#162440000000
0!
0%
#162445000000
1!
1%
#162450000000
0!
0%
#162455000000
1!
1%
#162460000000
0!
0%
#162465000000
1!
1%
#162470000000
0!
0%
#162475000000
1!
1%
#162480000000
0!
0%
#162485000000
1!
1%
#162490000000
0!
0%
#162495000000
1!
1%
#162500000000
0!
0%
#162505000000
1!
1%
#162510000000
0!
0%
#162515000000
1!
1%
#162520000000
0!
0%
#162525000000
1!
1%
#162530000000
0!
0%
#162535000000
1!
1%
#162540000000
0!
0%
#162545000000
1!
1%
#162550000000
0!
0%
#162555000000
1!
1%
#162560000000
0!
0%
#162565000000
1!
1%
#162570000000
0!
0%
#162575000000
1!
1%
#162580000000
0!
0%
#162585000000
1!
1%
#162590000000
0!
0%
#162595000000
1!
1%
#162600000000
0!
0%
#162605000000
1!
1%
#162610000000
0!
0%
#162615000000
1!
1%
#162620000000
0!
0%
#162625000000
1!
1%
#162630000000
0!
0%
#162635000000
1!
1%
#162640000000
0!
0%
#162645000000
1!
1%
#162650000000
0!
0%
#162655000000
1!
1%
#162660000000
0!
0%
#162665000000
1!
1%
#162670000000
0!
0%
#162675000000
1!
1%
#162680000000
0!
0%
#162685000000
1!
1%
#162690000000
0!
0%
#162695000000
1!
1%
#162700000000
0!
0%
#162705000000
1!
1%
#162710000000
0!
0%
#162715000000
1!
1%
#162720000000
0!
0%
#162725000000
1!
1%
#162730000000
0!
0%
#162735000000
1!
1%
#162740000000
0!
0%
#162745000000
1!
1%
#162750000000
0!
0%
#162755000000
1!
1%
#162760000000
0!
0%
#162765000000
1!
1%
#162770000000
0!
0%
#162775000000
1!
1%
#162780000000
0!
0%
#162785000000
1!
1%
#162790000000
0!
0%
#162795000000
1!
1%
#162800000000
0!
0%
#162805000000
1!
1%
#162810000000
0!
0%
#162815000000
1!
1%
#162820000000
0!
0%
#162825000000
1!
1%
#162830000000
0!
0%
#162835000000
1!
1%
#162840000000
0!
0%
#162845000000
1!
1%
#162850000000
0!
0%
#162855000000
1!
1%
#162860000000
0!
0%
#162865000000
1!
1%
#162870000000
0!
0%
#162875000000
1!
1%
#162880000000
0!
0%
#162885000000
1!
1%
#162890000000
0!
0%
#162895000000
1!
1%
#162900000000
0!
0%
#162905000000
1!
1%
#162910000000
0!
0%
#162915000000
1!
1%
#162920000000
0!
0%
#162925000000
1!
1%
#162930000000
0!
0%
#162935000000
1!
1%
#162940000000
0!
0%
#162945000000
1!
1%
#162950000000
0!
0%
#162955000000
1!
1%
#162960000000
0!
0%
#162965000000
1!
1%
#162970000000
0!
0%
#162975000000
1!
1%
#162980000000
0!
0%
#162985000000
1!
1%
#162990000000
0!
0%
#162995000000
1!
1%
#163000000000
0!
0%
#163005000000
1!
1%
#163010000000
0!
0%
#163015000000
1!
1%
#163020000000
0!
0%
#163025000000
1!
1%
#163030000000
0!
0%
#163035000000
1!
1%
#163040000000
0!
0%
#163045000000
1!
1%
#163050000000
0!
0%
#163055000000
1!
1%
#163060000000
0!
0%
#163065000000
1!
1%
#163070000000
0!
0%
#163075000000
1!
1%
#163080000000
0!
0%
#163085000000
1!
1%
#163090000000
0!
0%
#163095000000
1!
1%
#163100000000
0!
0%
#163105000000
1!
1%
#163110000000
0!
0%
#163115000000
1!
1%
#163120000000
0!
0%
#163125000000
1!
1%
#163130000000
0!
0%
#163135000000
1!
1%
#163140000000
0!
0%
#163145000000
1!
1%
#163150000000
0!
0%
#163155000000
1!
1%
#163160000000
0!
0%
#163165000000
1!
1%
#163170000000
0!
0%
#163175000000
1!
1%
#163180000000
0!
0%
#163185000000
1!
1%
#163190000000
0!
0%
#163195000000
1!
1%
#163200000000
0!
0%
#163205000000
1!
1%
#163210000000
0!
0%
#163215000000
1!
1%
#163220000000
0!
0%
#163225000000
1!
1%
#163230000000
0!
0%
#163235000000
1!
1%
#163240000000
0!
0%
#163245000000
1!
1%
#163250000000
0!
0%
#163255000000
1!
1%
#163260000000
0!
0%
#163265000000
1!
1%
#163270000000
0!
0%
#163275000000
1!
1%
#163280000000
0!
0%
#163285000000
1!
1%
#163290000000
0!
0%
#163295000000
1!
1%
#163300000000
0!
0%
#163305000000
1!
1%
#163310000000
0!
0%
#163315000000
1!
1%
#163320000000
0!
0%
#163325000000
1!
1%
#163330000000
0!
0%
#163335000000
1!
1%
#163340000000
0!
0%
#163345000000
1!
1%
#163350000000
0!
0%
#163355000000
1!
1%
#163360000000
0!
0%
#163365000000
1!
1%
#163370000000
0!
0%
#163375000000
1!
1%
#163380000000
0!
0%
#163385000000
1!
1%
#163390000000
0!
0%
#163395000000
1!
1%
#163400000000
0!
0%
#163405000000
1!
1%
#163410000000
0!
0%
#163415000000
1!
1%
#163420000000
0!
0%
#163425000000
1!
1%
#163430000000
0!
0%
#163435000000
1!
1%
#163440000000
0!
0%
#163445000000
1!
1%
#163450000000
0!
0%
#163455000000
1!
1%
#163460000000
0!
0%
#163465000000
1!
1%
#163470000000
0!
0%
#163475000000
1!
1%
#163480000000
0!
0%
#163485000000
1!
1%
#163490000000
0!
0%
#163495000000
1!
1%
#163500000000
0!
0%
#163505000000
1!
1%
#163510000000
0!
0%
#163515000000
1!
1%
#163520000000
0!
0%
#163525000000
1!
1%
#163530000000
0!
0%
#163535000000
1!
1%
#163540000000
0!
0%
#163545000000
1!
1%
#163550000000
0!
0%
#163555000000
1!
1%
#163560000000
0!
0%
#163565000000
1!
1%
#163570000000
0!
0%
#163575000000
1!
1%
#163580000000
0!
0%
#163585000000
1!
1%
#163590000000
0!
0%
#163595000000
1!
1%
#163600000000
0!
0%
#163605000000
1!
1%
#163610000000
0!
0%
#163615000000
1!
1%
#163620000000
0!
0%
#163625000000
1!
1%
#163630000000
0!
0%
#163635000000
1!
1%
#163640000000
0!
0%
#163645000000
1!
1%
#163650000000
0!
0%
#163655000000
1!
1%
#163660000000
0!
0%
#163665000000
1!
1%
#163670000000
0!
0%
#163675000000
1!
1%
#163680000000
0!
0%
#163685000000
1!
1%
#163690000000
0!
0%
#163695000000
1!
1%
#163700000000
0!
0%
#163705000000
1!
1%
#163710000000
0!
0%
#163715000000
1!
1%
#163720000000
0!
0%
#163725000000
1!
1%
#163730000000
0!
0%
#163735000000
1!
1%
#163740000000
0!
0%
#163745000000
1!
1%
#163750000000
0!
0%
#163755000000
1!
1%
#163760000000
0!
0%
#163765000000
1!
1%
#163770000000
0!
0%
#163775000000
1!
1%
#163780000000
0!
0%
#163785000000
1!
1%
#163790000000
0!
0%
#163795000000
1!
1%
#163800000000
0!
0%
#163805000000
1!
1%
#163810000000
0!
0%
#163815000000
1!
1%
#163820000000
0!
0%
#163825000000
1!
1%
#163830000000
0!
0%
#163835000000
1!
1%
#163840000000
0!
0%
#163845000000
1!
1%
#163850000000
0!
0%
#163855000000
1!
1%
#163860000000
0!
0%
#163865000000
1!
1%
#163870000000
0!
0%
#163875000000
1!
1%
#163880000000
0!
0%
#163885000000
1!
1%
#163890000000
0!
0%
#163895000000
1!
1%
#163900000000
0!
0%
#163905000000
1!
1%
#163910000000
0!
0%
#163915000000
1!
1%
#163920000000
0!
0%
#163925000000
1!
1%
#163930000000
0!
0%
#163935000000
1!
1%
#163940000000
0!
0%
#163945000000
1!
1%
#163950000000
0!
0%
#163955000000
1!
1%
#163960000000
0!
0%
#163965000000
1!
1%
#163970000000
0!
0%
#163975000000
1!
1%
#163980000000
0!
0%
#163985000000
1!
1%
#163990000000
0!
0%
#163995000000
1!
1%
#164000000000
0!
0%
#164005000000
1!
1%
#164010000000
0!
0%
#164015000000
1!
1%
#164020000000
0!
0%
#164025000000
1!
1%
#164030000000
0!
0%
#164035000000
1!
1%
#164040000000
0!
0%
#164045000000
1!
1%
#164050000000
0!
0%
#164055000000
1!
1%
#164060000000
0!
0%
#164065000000
1!
1%
#164070000000
0!
0%
#164075000000
1!
1%
#164080000000
0!
0%
#164085000000
1!
1%
#164090000000
0!
0%
#164095000000
1!
1%
#164100000000
0!
0%
#164105000000
1!
1%
#164110000000
0!
0%
#164115000000
1!
1%
#164120000000
0!
0%
#164125000000
1!
1%
#164130000000
0!
0%
#164135000000
1!
1%
#164140000000
0!
0%
#164145000000
1!
1%
#164150000000
0!
0%
#164155000000
1!
1%
#164160000000
0!
0%
#164165000000
1!
1%
#164170000000
0!
0%
#164175000000
1!
1%
#164180000000
0!
0%
#164185000000
1!
1%
#164190000000
0!
0%
#164195000000
1!
1%
#164200000000
0!
0%
#164205000000
1!
1%
#164210000000
0!
0%
#164215000000
1!
1%
#164220000000
0!
0%
#164225000000
1!
1%
#164230000000
0!
0%
#164235000000
1!
1%
#164240000000
0!
0%
#164245000000
1!
1%
#164250000000
0!
0%
#164255000000
1!
1%
#164260000000
0!
0%
#164265000000
1!
1%
#164270000000
0!
0%
#164275000000
1!
1%
#164280000000
0!
0%
#164285000000
1!
1%
#164290000000
0!
0%
#164295000000
1!
1%
#164300000000
0!
0%
#164305000000
1!
1%
#164310000000
0!
0%
#164315000000
1!
1%
#164320000000
0!
0%
#164325000000
1!
1%
#164330000000
0!
0%
#164335000000
1!
1%
#164340000000
0!
0%
#164345000000
1!
1%
#164350000000
0!
0%
#164355000000
1!
1%
#164360000000
0!
0%
#164365000000
1!
1%
#164370000000
0!
0%
#164375000000
1!
1%
#164380000000
0!
0%
#164385000000
1!
1%
#164390000000
0!
0%
#164395000000
1!
1%
#164400000000
0!
0%
#164405000000
1!
1%
#164410000000
0!
0%
#164415000000
1!
1%
#164420000000
0!
0%
#164425000000
1!
1%
#164430000000
0!
0%
#164435000000
1!
1%
#164440000000
0!
0%
#164445000000
1!
1%
#164450000000
0!
0%
#164455000000
1!
1%
#164460000000
0!
0%
#164465000000
1!
1%
#164470000000
0!
0%
#164475000000
1!
1%
#164480000000
0!
0%
#164485000000
1!
1%
#164490000000
0!
0%
#164495000000
1!
1%
#164500000000
0!
0%
#164505000000
1!
1%
#164510000000
0!
0%
#164515000000
1!
1%
#164520000000
0!
0%
#164525000000
1!
1%
#164530000000
0!
0%
#164535000000
1!
1%
#164540000000
0!
0%
#164545000000
1!
1%
#164550000000
0!
0%
#164555000000
1!
1%
#164560000000
0!
0%
#164565000000
1!
1%
#164570000000
0!
0%
#164575000000
1!
1%
#164580000000
0!
0%
#164585000000
1!
1%
#164590000000
0!
0%
#164595000000
1!
1%
#164600000000
0!
0%
#164605000000
1!
1%
#164610000000
0!
0%
#164615000000
1!
1%
#164620000000
0!
0%
#164625000000
1!
1%
#164630000000
0!
0%
#164635000000
1!
1%
#164640000000
0!
0%
#164645000000
1!
1%
#164650000000
0!
0%
#164655000000
1!
1%
#164660000000
0!
0%
#164665000000
1!
1%
#164670000000
0!
0%
#164675000000
1!
1%
#164680000000
0!
0%
#164685000000
1!
1%
#164690000000
0!
0%
#164695000000
1!
1%
#164700000000
0!
0%
#164705000000
1!
1%
#164710000000
0!
0%
#164715000000
1!
1%
#164720000000
0!
0%
#164725000000
1!
1%
#164730000000
0!
0%
#164735000000
1!
1%
#164740000000
0!
0%
#164745000000
1!
1%
#164750000000
0!
0%
#164755000000
1!
1%
#164760000000
0!
0%
#164765000000
1!
1%
#164770000000
0!
0%
#164775000000
1!
1%
#164780000000
0!
0%
#164785000000
1!
1%
#164790000000
0!
0%
#164795000000
1!
1%
#164800000000
0!
0%
#164805000000
1!
1%
#164810000000
0!
0%
#164815000000
1!
1%
#164820000000
0!
0%
#164825000000
1!
1%
#164830000000
0!
0%
#164835000000
1!
1%
#164840000000
0!
0%
#164845000000
1!
1%
#164850000000
0!
0%
#164855000000
1!
1%
#164860000000
0!
0%
#164865000000
1!
1%
#164870000000
0!
0%
#164875000000
1!
1%
#164880000000
0!
0%
#164885000000
1!
1%
#164890000000
0!
0%
#164895000000
1!
1%
#164900000000
0!
0%
#164905000000
1!
1%
#164910000000
0!
0%
#164915000000
1!
1%
#164920000000
0!
0%
#164925000000
1!
1%
#164930000000
0!
0%
#164935000000
1!
1%
#164940000000
0!
0%
#164945000000
1!
1%
#164950000000
0!
0%
#164955000000
1!
1%
#164960000000
0!
0%
#164965000000
1!
1%
#164970000000
0!
0%
#164975000000
1!
1%
#164980000000
0!
0%
#164985000000
1!
1%
#164990000000
0!
0%
#164995000000
1!
1%
#165000000000
0!
0%
#165005000000
1!
1%
#165010000000
0!
0%
#165015000000
1!
1%
#165020000000
0!
0%
#165025000000
1!
1%
#165030000000
0!
0%
#165035000000
1!
1%
#165040000000
0!
0%
#165045000000
1!
1%
#165050000000
0!
0%
#165055000000
1!
1%
#165060000000
0!
0%
#165065000000
1!
1%
#165070000000
0!
0%
#165075000000
1!
1%
#165080000000
0!
0%
#165085000000
1!
1%
#165090000000
0!
0%
#165095000000
1!
1%
#165100000000
0!
0%
#165105000000
1!
1%
#165110000000
0!
0%
#165115000000
1!
1%
#165120000000
0!
0%
#165125000000
1!
1%
#165130000000
0!
0%
#165135000000
1!
1%
#165140000000
0!
0%
#165145000000
1!
1%
#165150000000
0!
0%
#165155000000
1!
1%
#165160000000
0!
0%
#165165000000
1!
1%
#165170000000
0!
0%
#165175000000
1!
1%
#165180000000
0!
0%
#165185000000
1!
1%
#165190000000
0!
0%
#165195000000
1!
1%
#165200000000
0!
0%
#165205000000
1!
1%
#165210000000
0!
0%
#165215000000
1!
1%
#165220000000
0!
0%
#165225000000
1!
1%
#165230000000
0!
0%
#165235000000
1!
1%
#165240000000
0!
0%
#165245000000
1!
1%
#165250000000
0!
0%
#165255000000
1!
1%
#165260000000
0!
0%
#165265000000
1!
1%
#165270000000
0!
0%
#165275000000
1!
1%
#165280000000
0!
0%
#165285000000
1!
1%
#165290000000
0!
0%
#165295000000
1!
1%
#165300000000
0!
0%
#165305000000
1!
1%
#165310000000
0!
0%
#165315000000
1!
1%
#165320000000
0!
0%
#165325000000
1!
1%
#165330000000
0!
0%
#165335000000
1!
1%
#165340000000
0!
0%
#165345000000
1!
1%
#165350000000
0!
0%
#165355000000
1!
1%
#165360000000
0!
0%
#165365000000
1!
1%
#165370000000
0!
0%
#165375000000
1!
1%
#165380000000
0!
0%
#165385000000
1!
1%
#165390000000
0!
0%
#165395000000
1!
1%
#165400000000
0!
0%
#165405000000
1!
1%
#165410000000
0!
0%
#165415000000
1!
1%
#165420000000
0!
0%
#165425000000
1!
1%
#165430000000
0!
0%
#165435000000
1!
1%
#165440000000
0!
0%
#165445000000
1!
1%
#165450000000
0!
0%
#165455000000
1!
1%
#165460000000
0!
0%
#165465000000
1!
1%
#165470000000
0!
0%
#165475000000
1!
1%
#165480000000
0!
0%
#165485000000
1!
1%
#165490000000
0!
0%
#165495000000
1!
1%
#165500000000
0!
0%
#165505000000
1!
1%
#165510000000
0!
0%
#165515000000
1!
1%
#165520000000
0!
0%
#165525000000
1!
1%
#165530000000
0!
0%
#165535000000
1!
1%
#165540000000
0!
0%
#165545000000
1!
1%
#165550000000
0!
0%
#165555000000
1!
1%
#165560000000
0!
0%
#165565000000
1!
1%
#165570000000
0!
0%
#165575000000
1!
1%
#165580000000
0!
0%
#165585000000
1!
1%
#165590000000
0!
0%
#165595000000
1!
1%
#165600000000
0!
0%
#165605000000
1!
1%
#165610000000
0!
0%
#165615000000
1!
1%
#165620000000
0!
0%
#165625000000
1!
1%
#165630000000
0!
0%
#165635000000
1!
1%
#165640000000
0!
0%
#165645000000
1!
1%
#165650000000
0!
0%
#165655000000
1!
1%
#165660000000
0!
0%
#165665000000
1!
1%
#165670000000
0!
0%
#165675000000
1!
1%
#165680000000
0!
0%
#165685000000
1!
1%
#165690000000
0!
0%
#165695000000
1!
1%
#165700000000
0!
0%
#165705000000
1!
1%
#165710000000
0!
0%
#165715000000
1!
1%
#165720000000
0!
0%
#165725000000
1!
1%
#165730000000
0!
0%
#165735000000
1!
1%
#165740000000
0!
0%
#165745000000
1!
1%
#165750000000
0!
0%
#165755000000
1!
1%
#165760000000
0!
0%
#165765000000
1!
1%
#165770000000
0!
0%
#165775000000
1!
1%
#165780000000
0!
0%
#165785000000
1!
1%
#165790000000
0!
0%
#165795000000
1!
1%
#165800000000
0!
0%
#165805000000
1!
1%
#165810000000
0!
0%
#165815000000
1!
1%
#165820000000
0!
0%
#165825000000
1!
1%
#165830000000
0!
0%
#165835000000
1!
1%
#165840000000
0!
0%
#165845000000
1!
1%
#165850000000
0!
0%
#165855000000
1!
1%
#165860000000
0!
0%
#165865000000
1!
1%
#165870000000
0!
0%
#165875000000
1!
1%
#165880000000
0!
0%
#165885000000
1!
1%
#165890000000
0!
0%
#165895000000
1!
1%
#165900000000
0!
0%
#165905000000
1!
1%
#165910000000
0!
0%
#165915000000
1!
1%
#165920000000
0!
0%
#165925000000
1!
1%
#165930000000
0!
0%
#165935000000
1!
1%
#165940000000
0!
0%
#165945000000
1!
1%
#165950000000
0!
0%
#165955000000
1!
1%
#165960000000
0!
0%
#165965000000
1!
1%
#165970000000
0!
0%
#165975000000
1!
1%
#165980000000
0!
0%
#165985000000
1!
1%
#165990000000
0!
0%
#165995000000
1!
1%
#166000000000
0!
0%
#166005000000
1!
1%
#166010000000
0!
0%
#166015000000
1!
1%
#166020000000
0!
0%
#166025000000
1!
1%
#166030000000
0!
0%
#166035000000
1!
1%
#166040000000
0!
0%
#166045000000
1!
1%
#166050000000
0!
0%
#166055000000
1!
1%
#166060000000
0!
0%
#166065000000
1!
1%
#166070000000
0!
0%
#166075000000
1!
1%
#166080000000
0!
0%
#166085000000
1!
1%
#166090000000
0!
0%
#166095000000
1!
1%
#166100000000
0!
0%
#166105000000
1!
1%
#166110000000
0!
0%
#166115000000
1!
1%
#166120000000
0!
0%
#166125000000
1!
1%
#166130000000
0!
0%
#166135000000
1!
1%
#166140000000
0!
0%
#166145000000
1!
1%
#166150000000
0!
0%
#166155000000
1!
1%
#166160000000
0!
0%
#166165000000
1!
1%
#166170000000
0!
0%
#166175000000
1!
1%
#166180000000
0!
0%
#166185000000
1!
1%
#166190000000
0!
0%
#166195000000
1!
1%
#166200000000
0!
0%
#166205000000
1!
1%
#166210000000
0!
0%
#166215000000
1!
1%
#166220000000
0!
0%
#166225000000
1!
1%
#166230000000
0!
0%
#166235000000
1!
1%
#166240000000
0!
0%
#166245000000
1!
1%
#166250000000
0!
0%
#166255000000
1!
1%
#166260000000
0!
0%
#166265000000
1!
1%
#166270000000
0!
0%
#166275000000
1!
1%
#166280000000
0!
0%
#166285000000
1!
1%
#166290000000
0!
0%
#166295000000
1!
1%
#166300000000
0!
0%
#166305000000
1!
1%
#166310000000
0!
0%
#166315000000
1!
1%
#166320000000
0!
0%
#166325000000
1!
1%
#166330000000
0!
0%
#166335000000
1!
1%
#166340000000
0!
0%
#166345000000
1!
1%
#166350000000
0!
0%
#166355000000
1!
1%
#166360000000
0!
0%
#166365000000
1!
1%
#166370000000
0!
0%
#166375000000
1!
1%
#166380000000
0!
0%
#166385000000
1!
1%
#166390000000
0!
0%
#166395000000
1!
1%
#166400000000
0!
0%
#166405000000
1!
1%
#166410000000
0!
0%
#166415000000
1!
1%
#166420000000
0!
0%
#166425000000
1!
1%
#166430000000
0!
0%
#166435000000
1!
1%
#166440000000
0!
0%
#166445000000
1!
1%
#166450000000
0!
0%
#166455000000
1!
1%
#166460000000
0!
0%
#166465000000
1!
1%
#166470000000
0!
0%
#166475000000
1!
1%
#166480000000
0!
0%
#166485000000
1!
1%
#166490000000
0!
0%
#166495000000
1!
1%
#166500000000
0!
0%
#166505000000
1!
1%
#166510000000
0!
0%
#166515000000
1!
1%
#166520000000
0!
0%
#166525000000
1!
1%
#166530000000
0!
0%
#166535000000
1!
1%
#166540000000
0!
0%
#166545000000
1!
1%
#166550000000
0!
0%
#166555000000
1!
1%
#166560000000
0!
0%
#166565000000
1!
1%
#166570000000
0!
0%
#166575000000
1!
1%
#166580000000
0!
0%
#166585000000
1!
1%
#166590000000
0!
0%
#166595000000
1!
1%
#166600000000
0!
0%
#166605000000
1!
1%
#166610000000
0!
0%
#166615000000
1!
1%
#166620000000
0!
0%
#166625000000
1!
1%
#166630000000
0!
0%
#166635000000
1!
1%
#166640000000
0!
0%
#166645000000
1!
1%
#166650000000
0!
0%
#166655000000
1!
1%
#166660000000
0!
0%
#166665000000
1!
1%
#166670000000
0!
0%
#166675000000
1!
1%
#166680000000
0!
0%
#166685000000
1!
1%
#166690000000
0!
0%
#166695000000
1!
1%
#166700000000
0!
0%
#166705000000
1!
1%
#166710000000
0!
0%
#166715000000
1!
1%
#166720000000
0!
0%
#166725000000
1!
1%
#166730000000
0!
0%
#166735000000
1!
1%
#166740000000
0!
0%
#166745000000
1!
1%
#166750000000
0!
0%
#166755000000
1!
1%
#166760000000
0!
0%
#166765000000
1!
1%
#166770000000
0!
0%
#166775000000
1!
1%
#166780000000
0!
0%
#166785000000
1!
1%
#166790000000
0!
0%
#166795000000
1!
1%
#166800000000
0!
0%
#166805000000
1!
1%
#166810000000
0!
0%
#166815000000
1!
1%
#166820000000
0!
0%
#166825000000
1!
1%
#166830000000
0!
0%
#166835000000
1!
1%
#166840000000
0!
0%
#166845000000
1!
1%
#166850000000
0!
0%
#166855000000
1!
1%
#166860000000
0!
0%
#166865000000
1!
1%
#166870000000
0!
0%
#166875000000
1!
1%
#166880000000
0!
0%
#166885000000
1!
1%
#166890000000
0!
0%
#166895000000
1!
1%
#166900000000
0!
0%
#166905000000
1!
1%
#166910000000
0!
0%
#166915000000
1!
1%
#166920000000
0!
0%
#166925000000
1!
1%
#166930000000
0!
0%
#166935000000
1!
1%
#166940000000
0!
0%
#166945000000
1!
1%
#166950000000
0!
0%
#166955000000
1!
1%
#166960000000
0!
0%
#166965000000
1!
1%
#166970000000
0!
0%
#166975000000
1!
1%
#166980000000
0!
0%
#166985000000
1!
1%
#166990000000
0!
0%
#166995000000
1!
1%
#167000000000
0!
0%
#167005000000
1!
1%
#167010000000
0!
0%
#167015000000
1!
1%
#167020000000
0!
0%
#167025000000
1!
1%
#167030000000
0!
0%
#167035000000
1!
1%
#167040000000
0!
0%
#167045000000
1!
1%
#167050000000
0!
0%
#167055000000
1!
1%
#167060000000
0!
0%
#167065000000
1!
1%
#167070000000
0!
0%
#167075000000
1!
1%
#167080000000
0!
0%
#167085000000
1!
1%
#167090000000
0!
0%
#167095000000
1!
1%
#167100000000
0!
0%
#167105000000
1!
1%
#167110000000
0!
0%
#167115000000
1!
1%
#167120000000
0!
0%
#167125000000
1!
1%
#167130000000
0!
0%
#167135000000
1!
1%
#167140000000
0!
0%
#167145000000
1!
1%
#167150000000
0!
0%
#167155000000
1!
1%
#167160000000
0!
0%
#167165000000
1!
1%
#167170000000
0!
0%
#167175000000
1!
1%
#167180000000
0!
0%
#167185000000
1!
1%
#167190000000
0!
0%
#167195000000
1!
1%
#167200000000
0!
0%
#167205000000
1!
1%
#167210000000
0!
0%
#167215000000
1!
1%
#167220000000
0!
0%
#167225000000
1!
1%
#167230000000
0!
0%
#167235000000
1!
1%
#167240000000
0!
0%
#167245000000
1!
1%
#167250000000
0!
0%
#167255000000
1!
1%
#167260000000
0!
0%
#167265000000
1!
1%
#167270000000
0!
0%
#167275000000
1!
1%
#167280000000
0!
0%
#167285000000
1!
1%
#167290000000
0!
0%
#167295000000
1!
1%
#167300000000
0!
0%
#167305000000
1!
1%
#167310000000
0!
0%
#167315000000
1!
1%
#167320000000
0!
0%
#167325000000
1!
1%
#167330000000
0!
0%
#167335000000
1!
1%
#167340000000
0!
0%
#167345000000
1!
1%
#167350000000
0!
0%
#167355000000
1!
1%
#167360000000
0!
0%
#167365000000
1!
1%
#167370000000
0!
0%
#167375000000
1!
1%
#167380000000
0!
0%
#167385000000
1!
1%
#167390000000
0!
0%
#167395000000
1!
1%
#167400000000
0!
0%
#167405000000
1!
1%
#167410000000
0!
0%
#167415000000
1!
1%
#167420000000
0!
0%
#167425000000
1!
1%
#167430000000
0!
0%
#167435000000
1!
1%
#167440000000
0!
0%
#167445000000
1!
1%
#167450000000
0!
0%
#167455000000
1!
1%
#167460000000
0!
0%
#167465000000
1!
1%
#167470000000
0!
0%
#167475000000
1!
1%
#167480000000
0!
0%
#167485000000
1!
1%
#167490000000
0!
0%
#167495000000
1!
1%
#167500000000
0!
0%
#167505000000
1!
1%
#167510000000
0!
0%
#167515000000
1!
1%
#167520000000
0!
0%
#167525000000
1!
1%
#167530000000
0!
0%
#167535000000
1!
1%
#167540000000
0!
0%
#167545000000
1!
1%
#167550000000
0!
0%
#167555000000
1!
1%
#167560000000
0!
0%
#167565000000
1!
1%
#167570000000
0!
0%
#167575000000
1!
1%
#167580000000
0!
0%
#167585000000
1!
1%
#167590000000
0!
0%
#167595000000
1!
1%
#167600000000
0!
0%
#167605000000
1!
1%
#167610000000
0!
0%
#167615000000
1!
1%
#167620000000
0!
0%
#167625000000
1!
1%
#167630000000
0!
0%
#167635000000
1!
1%
#167640000000
0!
0%
#167645000000
1!
1%
#167650000000
0!
0%
#167655000000
1!
1%
#167660000000
0!
0%
#167665000000
1!
1%
#167670000000
0!
0%
#167675000000
1!
1%
#167680000000
0!
0%
#167685000000
1!
1%
#167690000000
0!
0%
#167695000000
1!
1%
#167700000000
0!
0%
#167705000000
1!
1%
#167710000000
0!
0%
#167715000000
1!
1%
#167720000000
0!
0%
#167725000000
1!
1%
#167730000000
0!
0%
#167735000000
1!
1%
#167740000000
0!
0%
#167745000000
1!
1%
#167750000000
0!
0%
#167755000000
1!
1%
#167760000000
0!
0%
#167765000000
1!
1%
#167770000000
0!
0%
#167775000000
1!
1%
#167780000000
0!
0%
#167785000000
1!
1%
#167790000000
0!
0%
#167795000000
1!
1%
#167800000000
0!
0%
#167805000000
1!
1%
#167810000000
0!
0%
#167815000000
1!
1%
#167820000000
0!
0%
#167825000000
1!
1%
#167830000000
0!
0%
#167835000000
1!
1%
#167840000000
0!
0%
#167845000000
1!
1%
#167850000000
0!
0%
#167855000000
1!
1%
#167860000000
0!
0%
#167865000000
1!
1%
#167870000000
0!
0%
#167875000000
1!
1%
#167880000000
0!
0%
#167885000000
1!
1%
#167890000000
0!
0%
#167895000000
1!
1%
#167900000000
0!
0%
#167905000000
1!
1%
#167910000000
0!
0%
#167915000000
1!
1%
#167920000000
0!
0%
#167925000000
1!
1%
#167930000000
0!
0%
#167935000000
1!
1%
#167940000000
0!
0%
#167945000000
1!
1%
#167950000000
0!
0%
#167955000000
1!
1%
#167960000000
0!
0%
#167965000000
1!
1%
#167970000000
0!
0%
#167975000000
1!
1%
#167980000000
0!
0%
#167985000000
1!
1%
#167990000000
0!
0%
#167995000000
1!
1%
#168000000000
0!
0%
#168005000000
1!
1%
#168010000000
0!
0%
#168015000000
1!
1%
#168020000000
0!
0%
#168025000000
1!
1%
#168030000000
0!
0%
#168035000000
1!
1%
#168040000000
0!
0%
#168045000000
1!
1%
#168050000000
0!
0%
#168055000000
1!
1%
#168060000000
0!
0%
#168065000000
1!
1%
#168070000000
0!
0%
#168075000000
1!
1%
#168080000000
0!
0%
#168085000000
1!
1%
#168090000000
0!
0%
#168095000000
1!
1%
#168100000000
0!
0%
#168105000000
1!
1%
#168110000000
0!
0%
#168115000000
1!
1%
#168120000000
0!
0%
#168125000000
1!
1%
#168130000000
0!
0%
#168135000000
1!
1%
#168140000000
0!
0%
#168145000000
1!
1%
#168150000000
0!
0%
#168155000000
1!
1%
#168160000000
0!
0%
#168165000000
1!
1%
#168170000000
0!
0%
#168175000000
1!
1%
#168180000000
0!
0%
#168185000000
1!
1%
#168190000000
0!
0%
#168195000000
1!
1%
#168200000000
0!
0%
#168205000000
1!
1%
#168210000000
0!
0%
#168215000000
1!
1%
#168220000000
0!
0%
#168225000000
1!
1%
#168230000000
0!
0%
#168235000000
1!
1%
#168240000000
0!
0%
#168245000000
1!
1%
#168250000000
0!
0%
#168255000000
1!
1%
#168260000000
0!
0%
#168265000000
1!
1%
#168270000000
0!
0%
#168275000000
1!
1%
#168280000000
0!
0%
#168285000000
1!
1%
#168290000000
0!
0%
#168295000000
1!
1%
#168300000000
0!
0%
#168305000000
1!
1%
#168310000000
0!
0%
#168315000000
1!
1%
#168320000000
0!
0%
#168325000000
1!
1%
#168330000000
0!
0%
#168335000000
1!
1%
#168340000000
0!
0%
#168345000000
1!
1%
#168350000000
0!
0%
#168355000000
1!
1%
#168360000000
0!
0%
#168365000000
1!
1%
#168370000000
0!
0%
#168375000000
1!
1%
#168380000000
0!
0%
#168385000000
1!
1%
#168390000000
0!
0%
#168395000000
1!
1%
#168400000000
0!
0%
#168405000000
1!
1%
#168410000000
0!
0%
#168415000000
1!
1%
#168420000000
0!
0%
#168425000000
1!
1%
#168430000000
0!
0%
#168435000000
1!
1%
#168440000000
0!
0%
#168445000000
1!
1%
#168450000000
0!
0%
#168455000000
1!
1%
#168460000000
0!
0%
#168465000000
1!
1%
#168470000000
0!
0%
#168475000000
1!
1%
#168480000000
0!
0%
#168485000000
1!
1%
#168490000000
0!
0%
#168495000000
1!
1%
#168500000000
0!
0%
#168505000000
1!
1%
#168510000000
0!
0%
#168515000000
1!
1%
#168520000000
0!
0%
#168525000000
1!
1%
#168530000000
0!
0%
#168535000000
1!
1%
#168540000000
0!
0%
#168545000000
1!
1%
#168550000000
0!
0%
#168555000000
1!
1%
#168560000000
0!
0%
#168565000000
1!
1%
#168570000000
0!
0%
#168575000000
1!
1%
#168580000000
0!
0%
#168585000000
1!
1%
#168590000000
0!
0%
#168595000000
1!
1%
#168600000000
0!
0%
#168605000000
1!
1%
#168610000000
0!
0%
#168615000000
1!
1%
#168620000000
0!
0%
#168625000000
1!
1%
#168630000000
0!
0%
#168635000000
1!
1%
#168640000000
0!
0%
#168645000000
1!
1%
#168650000000
0!
0%
#168655000000
1!
1%
#168660000000
0!
0%
#168665000000
1!
1%
#168670000000
0!
0%
#168675000000
1!
1%
#168680000000
0!
0%
#168685000000
1!
1%
#168690000000
0!
0%
#168695000000
1!
1%
#168700000000
0!
0%
#168705000000
1!
1%
#168710000000
0!
0%
#168715000000
1!
1%
#168720000000
0!
0%
#168725000000
1!
1%
#168730000000
0!
0%
#168735000000
1!
1%
#168740000000
0!
0%
#168745000000
1!
1%
#168750000000
0!
0%
#168755000000
1!
1%
#168760000000
0!
0%
#168765000000
1!
1%
#168770000000
0!
0%
#168775000000
1!
1%
#168780000000
0!
0%
#168785000000
1!
1%
#168790000000
0!
0%
#168795000000
1!
1%
#168800000000
0!
0%
#168805000000
1!
1%
#168810000000
0!
0%
#168815000000
1!
1%
#168820000000
0!
0%
#168825000000
1!
1%
#168830000000
0!
0%
#168835000000
1!
1%
#168840000000
0!
0%
#168845000000
1!
1%
#168850000000
0!
0%
#168855000000
1!
1%
#168860000000
0!
0%
#168865000000
1!
1%
#168870000000
0!
0%
#168875000000
1!
1%
#168880000000
0!
0%
#168885000000
1!
1%
#168890000000
0!
0%
#168895000000
1!
1%
#168900000000
0!
0%
#168905000000
1!
1%
#168910000000
0!
0%
#168915000000
1!
1%
#168920000000
0!
0%
#168925000000
1!
1%
#168930000000
0!
0%
#168935000000
1!
1%
#168940000000
0!
0%
#168945000000
1!
1%
#168950000000
0!
0%
#168955000000
1!
1%
#168960000000
0!
0%
#168965000000
1!
1%
#168970000000
0!
0%
#168975000000
1!
1%
#168980000000
0!
0%
#168985000000
1!
1%
#168990000000
0!
0%
#168995000000
1!
1%
#169000000000
0!
0%
#169005000000
1!
1%
#169010000000
0!
0%
#169015000000
1!
1%
#169020000000
0!
0%
#169025000000
1!
1%
#169030000000
0!
0%
#169035000000
1!
1%
#169040000000
0!
0%
#169045000000
1!
1%
#169050000000
0!
0%
#169055000000
1!
1%
#169060000000
0!
0%
#169065000000
1!
1%
#169070000000
0!
0%
#169075000000
1!
1%
#169080000000
0!
0%
#169085000000
1!
1%
#169090000000
0!
0%
#169095000000
1!
1%
#169100000000
0!
0%
#169105000000
1!
1%
#169110000000
0!
0%
#169115000000
1!
1%
#169120000000
0!
0%
#169125000000
1!
1%
#169130000000
0!
0%
#169135000000
1!
1%
#169140000000
0!
0%
#169145000000
1!
1%
#169150000000
0!
0%
#169155000000
1!
1%
#169160000000
0!
0%
#169165000000
1!
1%
#169170000000
0!
0%
#169175000000
1!
1%
#169180000000
0!
0%
#169185000000
1!
1%
#169190000000
0!
0%
#169195000000
1!
1%
#169200000000
0!
0%
#169205000000
1!
1%
#169210000000
0!
0%
#169215000000
1!
1%
#169220000000
0!
0%
#169225000000
1!
1%
#169230000000
0!
0%
#169235000000
1!
1%
#169240000000
0!
0%
#169245000000
1!
1%
#169250000000
0!
0%
#169255000000
1!
1%
#169260000000
0!
0%
#169265000000
1!
1%
#169270000000
0!
0%
#169275000000
1!
1%
#169280000000
0!
0%
#169285000000
1!
1%
#169290000000
0!
0%
#169295000000
1!
1%
#169300000000
0!
0%
#169305000000
1!
1%
#169310000000
0!
0%
#169315000000
1!
1%
#169320000000
0!
0%
#169325000000
1!
1%
#169330000000
0!
0%
#169335000000
1!
1%
#169340000000
0!
0%
#169345000000
1!
1%
#169350000000
0!
0%
#169355000000
1!
1%
#169360000000
0!
0%
#169365000000
1!
1%
#169370000000
0!
0%
#169375000000
1!
1%
#169380000000
0!
0%
#169385000000
1!
1%
#169390000000
0!
0%
#169395000000
1!
1%
#169400000000
0!
0%
#169405000000
1!
1%
#169410000000
0!
0%
#169415000000
1!
1%
#169420000000
0!
0%
#169425000000
1!
1%
#169430000000
0!
0%
#169435000000
1!
1%
#169440000000
0!
0%
#169445000000
1!
1%
#169450000000
0!
0%
#169455000000
1!
1%
#169460000000
0!
0%
#169465000000
1!
1%
#169470000000
0!
0%
#169475000000
1!
1%
#169480000000
0!
0%
#169485000000
1!
1%
#169490000000
0!
0%
#169495000000
1!
1%
#169500000000
0!
0%
#169505000000
1!
1%
#169510000000
0!
0%
#169515000000
1!
1%
#169520000000
0!
0%
#169525000000
1!
1%
#169530000000
0!
0%
#169535000000
1!
1%
#169540000000
0!
0%
#169545000000
1!
1%
#169550000000
0!
0%
#169555000000
1!
1%
#169560000000
0!
0%
#169565000000
1!
1%
#169570000000
0!
0%
#169575000000
1!
1%
#169580000000
0!
0%
#169585000000
1!
1%
#169590000000
0!
0%
#169595000000
1!
1%
#169600000000
0!
0%
#169605000000
1!
1%
#169610000000
0!
0%
#169615000000
1!
1%
#169620000000
0!
0%
#169625000000
1!
1%
#169630000000
0!
0%
#169635000000
1!
1%
#169640000000
0!
0%
#169645000000
1!
1%
#169650000000
0!
0%
#169655000000
1!
1%
#169660000000
0!
0%
#169665000000
1!
1%
#169670000000
0!
0%
#169675000000
1!
1%
#169680000000
0!
0%
#169685000000
1!
1%
#169690000000
0!
0%
#169695000000
1!
1%
#169700000000
0!
0%
#169705000000
1!
1%
#169710000000
0!
0%
#169715000000
1!
1%
#169720000000
0!
0%
#169725000000
1!
1%
#169730000000
0!
0%
#169735000000
1!
1%
#169740000000
0!
0%
#169745000000
1!
1%
#169750000000
0!
0%
#169755000000
1!
1%
#169760000000
0!
0%
#169765000000
1!
1%
#169770000000
0!
0%
#169775000000
1!
1%
#169780000000
0!
0%
#169785000000
1!
1%
#169790000000
0!
0%
#169795000000
1!
1%
#169800000000
0!
0%
#169805000000
1!
1%
#169810000000
0!
0%
#169815000000
1!
1%
#169820000000
0!
0%
#169825000000
1!
1%
#169830000000
0!
0%
#169835000000
1!
1%
#169840000000
0!
0%
#169845000000
1!
1%
#169850000000
0!
0%
#169855000000
1!
1%
#169860000000
0!
0%
#169865000000
1!
1%
#169870000000
0!
0%
#169875000000
1!
1%
#169880000000
0!
0%
#169885000000
1!
1%
#169890000000
0!
0%
#169895000000
1!
1%
#169900000000
0!
0%
#169905000000
1!
1%
#169910000000
0!
0%
#169915000000
1!
1%
#169920000000
0!
0%
#169925000000
1!
1%
#169930000000
0!
0%
#169935000000
1!
1%
#169940000000
0!
0%
#169945000000
1!
1%
#169950000000
0!
0%
#169955000000
1!
1%
#169960000000
0!
0%
#169965000000
1!
1%
#169970000000
0!
0%
#169975000000
1!
1%
#169980000000
0!
0%
#169985000000
1!
1%
#169990000000
0!
0%
#169995000000
1!
1%
#170000000000
0!
0%
#170005000000
1!
1%
#170010000000
0!
0%
#170015000000
1!
1%
#170020000000
0!
0%
#170025000000
1!
1%
#170030000000
0!
0%
#170035000000
1!
1%
#170040000000
0!
0%
#170045000000
1!
1%
#170050000000
0!
0%
#170055000000
1!
1%
#170060000000
0!
0%
#170065000000
1!
1%
#170070000000
0!
0%
#170075000000
1!
1%
#170080000000
0!
0%
#170085000000
1!
1%
#170090000000
0!
0%
#170095000000
1!
1%
#170100000000
0!
0%
#170105000000
1!
1%
#170110000000
0!
0%
#170115000000
1!
1%
#170120000000
0!
0%
#170125000000
1!
1%
#170130000000
0!
0%
#170135000000
1!
1%
#170140000000
0!
0%
#170145000000
1!
1%
#170150000000
0!
0%
#170155000000
1!
1%
#170160000000
0!
0%
#170165000000
1!
1%
#170170000000
0!
0%
#170175000000
1!
1%
#170180000000
0!
0%
#170185000000
1!
1%
#170190000000
0!
0%
#170195000000
1!
1%
#170200000000
0!
0%
#170205000000
1!
1%
#170210000000
0!
0%
#170215000000
1!
1%
#170220000000
0!
0%
#170225000000
1!
1%
#170230000000
0!
0%
#170235000000
1!
1%
#170240000000
0!
0%
#170245000000
1!
1%
#170250000000
0!
0%
#170255000000
1!
1%
#170260000000
0!
0%
#170265000000
1!
1%
#170270000000
0!
0%
#170275000000
1!
1%
#170280000000
0!
0%
#170285000000
1!
1%
#170290000000
0!
0%
#170295000000
1!
1%
#170300000000
0!
0%
#170305000000
1!
1%
#170310000000
0!
0%
#170315000000
1!
1%
#170320000000
0!
0%
#170325000000
1!
1%
#170330000000
0!
0%
#170335000000
1!
1%
#170340000000
0!
0%
#170345000000
1!
1%
#170350000000
0!
0%
#170355000000
1!
1%
#170360000000
0!
0%
#170365000000
1!
1%
#170370000000
0!
0%
#170375000000
1!
1%
#170380000000
0!
0%
#170385000000
1!
1%
#170390000000
0!
0%
#170395000000
1!
1%
#170400000000
0!
0%
#170405000000
1!
1%
#170410000000
0!
0%
#170415000000
1!
1%
#170420000000
0!
0%
#170425000000
1!
1%
#170430000000
0!
0%
#170435000000
1!
1%
#170440000000
0!
0%
#170445000000
1!
1%
#170450000000
0!
0%
#170455000000
1!
1%
#170460000000
0!
0%
#170465000000
1!
1%
#170470000000
0!
0%
#170475000000
1!
1%
#170480000000
0!
0%
#170485000000
1!
1%
#170490000000
0!
0%
#170495000000
1!
1%
#170500000000
0!
0%
#170505000000
1!
1%
#170510000000
0!
0%
#170515000000
1!
1%
#170520000000
0!
0%
#170525000000
1!
1%
#170530000000
0!
0%
#170535000000
1!
1%
#170540000000
0!
0%
#170545000000
1!
1%
#170550000000
0!
0%
#170555000000
1!
1%
#170560000000
0!
0%
#170565000000
1!
1%
#170570000000
0!
0%
#170575000000
1!
1%
#170580000000
0!
0%
#170585000000
1!
1%
#170590000000
0!
0%
#170595000000
1!
1%
#170600000000
0!
0%
#170605000000
1!
1%
#170610000000
0!
0%
#170615000000
1!
1%
#170620000000
0!
0%
#170625000000
1!
1%
#170630000000
0!
0%
#170635000000
1!
1%
#170640000000
0!
0%
#170645000000
1!
1%
#170650000000
0!
0%
#170655000000
1!
1%
#170660000000
0!
0%
#170665000000
1!
1%
#170670000000
0!
0%
#170675000000
1!
1%
#170680000000
0!
0%
#170685000000
1!
1%
#170690000000
0!
0%
#170695000000
1!
1%
#170700000000
0!
0%
#170705000000
1!
1%
#170710000000
0!
0%
#170715000000
1!
1%
#170720000000
0!
0%
#170725000000
1!
1%
#170730000000
0!
0%
#170735000000
1!
1%
#170740000000
0!
0%
#170745000000
1!
1%
#170750000000
0!
0%
#170755000000
1!
1%
#170760000000
0!
0%
#170765000000
1!
1%
#170770000000
0!
0%
#170775000000
1!
1%
#170780000000
0!
0%
#170785000000
1!
1%
#170790000000
0!
0%
#170795000000
1!
1%
#170800000000
0!
0%
#170805000000
1!
1%
#170810000000
0!
0%
#170815000000
1!
1%
#170820000000
0!
0%
#170825000000
1!
1%
#170830000000
0!
0%
#170835000000
1!
1%
#170840000000
0!
0%
#170845000000
1!
1%
#170850000000
0!
0%
#170855000000
1!
1%
#170860000000
0!
0%
#170865000000
1!
1%
#170870000000
0!
0%
#170875000000
1!
1%
#170880000000
0!
0%
#170885000000
1!
1%
#170890000000
0!
0%
#170895000000
1!
1%
#170900000000
0!
0%
#170905000000
1!
1%
#170910000000
0!
0%
#170915000000
1!
1%
#170920000000
0!
0%
#170925000000
1!
1%
#170930000000
0!
0%
#170935000000
1!
1%
#170940000000
0!
0%
#170945000000
1!
1%
#170950000000
0!
0%
#170955000000
1!
1%
#170960000000
0!
0%
#170965000000
1!
1%
#170970000000
0!
0%
#170975000000
1!
1%
#170980000000
0!
0%
#170985000000
1!
1%
#170990000000
0!
0%
#170995000000
1!
1%
#171000000000
0!
0%
#171005000000
1!
1%
#171010000000
0!
0%
#171015000000
1!
1%
#171020000000
0!
0%
#171025000000
1!
1%
#171030000000
0!
0%
#171035000000
1!
1%
#171040000000
0!
0%
#171045000000
1!
1%
#171050000000
0!
0%
#171055000000
1!
1%
#171060000000
0!
0%
#171065000000
1!
1%
#171070000000
0!
0%
#171075000000
1!
1%
#171080000000
0!
0%
#171085000000
1!
1%
#171090000000
0!
0%
#171095000000
1!
1%
#171100000000
0!
0%
#171105000000
1!
1%
#171110000000
0!
0%
#171115000000
1!
1%
#171120000000
0!
0%
#171125000000
1!
1%
#171130000000
0!
0%
#171135000000
1!
1%
#171140000000
0!
0%
#171145000000
1!
1%
#171150000000
0!
0%
#171155000000
1!
1%
#171160000000
0!
0%
#171165000000
1!
1%
#171170000000
0!
0%
#171175000000
1!
1%
#171180000000
0!
0%
#171185000000
1!
1%
#171190000000
0!
0%
#171195000000
1!
1%
#171200000000
0!
0%
#171205000000
1!
1%
#171210000000
0!
0%
#171215000000
1!
1%
#171220000000
0!
0%
#171225000000
1!
1%
#171230000000
0!
0%
#171235000000
1!
1%
#171240000000
0!
0%
#171245000000
1!
1%
#171250000000
0!
0%
#171255000000
1!
1%
#171260000000
0!
0%
#171265000000
1!
1%
#171270000000
0!
0%
#171275000000
1!
1%
#171280000000
0!
0%
#171285000000
1!
1%
#171290000000
0!
0%
#171295000000
1!
1%
#171300000000
0!
0%
#171305000000
1!
1%
#171310000000
0!
0%
#171315000000
1!
1%
#171320000000
0!
0%
#171325000000
1!
1%
#171330000000
0!
0%
#171335000000
1!
1%
#171340000000
0!
0%
#171345000000
1!
1%
#171350000000
0!
0%
#171355000000
1!
1%
#171360000000
0!
0%
#171365000000
1!
1%
#171370000000
0!
0%
#171375000000
1!
1%
#171380000000
0!
0%
#171385000000
1!
1%
#171390000000
0!
0%
#171395000000
1!
1%
#171400000000
0!
0%
#171405000000
1!
1%
#171410000000
0!
0%
#171415000000
1!
1%
#171420000000
0!
0%
#171425000000
1!
1%
#171430000000
0!
0%
#171435000000
1!
1%
#171440000000
0!
0%
#171445000000
1!
1%
#171450000000
0!
0%
#171455000000
1!
1%
#171460000000
0!
0%
#171465000000
1!
1%
#171470000000
0!
0%
#171475000000
1!
1%
#171480000000
0!
0%
#171485000000
1!
1%
#171490000000
0!
0%
#171495000000
1!
1%
#171500000000
0!
0%
#171505000000
1!
1%
#171510000000
0!
0%
#171515000000
1!
1%
#171520000000
0!
0%
#171525000000
1!
1%
#171530000000
0!
0%
#171535000000
1!
1%
#171540000000
0!
0%
#171545000000
1!
1%
#171550000000
0!
0%
#171555000000
1!
1%
#171560000000
0!
0%
#171565000000
1!
1%
#171570000000
0!
0%
#171575000000
1!
1%
#171580000000
0!
0%
#171585000000
1!
1%
#171590000000
0!
0%
#171595000000
1!
1%
#171600000000
0!
0%
#171605000000
1!
1%
#171610000000
0!
0%
#171615000000
1!
1%
#171620000000
0!
0%
#171625000000
1!
1%
#171630000000
0!
0%
#171635000000
1!
1%
#171640000000
0!
0%
#171645000000
1!
1%
#171650000000
0!
0%
#171655000000
1!
1%
#171660000000
0!
0%
#171665000000
1!
1%
#171670000000
0!
0%
#171675000000
1!
1%
#171680000000
0!
0%
#171685000000
1!
1%
#171690000000
0!
0%
#171695000000
1!
1%
#171700000000
0!
0%
#171705000000
1!
1%
#171710000000
0!
0%
#171715000000
1!
1%
#171720000000
0!
0%
#171725000000
1!
1%
#171730000000
0!
0%
#171735000000
1!
1%
#171740000000
0!
0%
#171745000000
1!
1%
#171750000000
0!
0%
#171755000000
1!
1%
#171760000000
0!
0%
#171765000000
1!
1%
#171770000000
0!
0%
#171775000000
1!
1%
#171780000000
0!
0%
#171785000000
1!
1%
#171790000000
0!
0%
#171795000000
1!
1%
#171800000000
0!
0%
#171805000000
1!
1%
#171810000000
0!
0%
#171815000000
1!
1%
#171820000000
0!
0%
#171825000000
1!
1%
#171830000000
0!
0%
#171835000000
1!
1%
#171840000000
0!
0%
#171845000000
1!
1%
#171850000000
0!
0%
#171855000000
1!
1%
#171860000000
0!
0%
#171865000000
1!
1%
#171870000000
0!
0%
#171875000000
1!
1%
#171880000000
0!
0%
#171885000000
1!
1%
#171890000000
0!
0%
#171895000000
1!
1%
#171900000000
0!
0%
#171905000000
1!
1%
#171910000000
0!
0%
#171915000000
1!
1%
#171920000000
0!
0%
#171925000000
1!
1%
#171930000000
0!
0%
#171935000000
1!
1%
#171940000000
0!
0%
#171945000000
1!
1%
#171950000000
0!
0%
#171955000000
1!
1%
#171960000000
0!
0%
#171965000000
1!
1%
#171970000000
0!
0%
#171975000000
1!
1%
#171980000000
0!
0%
#171985000000
1!
1%
#171990000000
0!
0%
#171995000000
1!
1%
#172000000000
0!
0%
#172005000000
1!
1%
#172010000000
0!
0%
#172015000000
1!
1%
#172020000000
0!
0%
#172025000000
1!
1%
#172030000000
0!
0%
#172035000000
1!
1%
#172040000000
0!
0%
#172045000000
1!
1%
#172050000000
0!
0%
#172055000000
1!
1%
#172060000000
0!
0%
#172065000000
1!
1%
#172070000000
0!
0%
#172075000000
1!
1%
#172080000000
0!
0%
#172085000000
1!
1%
#172090000000
0!
0%
#172095000000
1!
1%
#172100000000
0!
0%
#172105000000
1!
1%
#172110000000
0!
0%
#172115000000
1!
1%
#172120000000
0!
0%
#172125000000
1!
1%
#172130000000
0!
0%
#172135000000
1!
1%
#172140000000
0!
0%
#172145000000
1!
1%
#172150000000
0!
0%
#172155000000
1!
1%
#172160000000
0!
0%
#172165000000
1!
1%
#172170000000
0!
0%
#172175000000
1!
1%
#172180000000
0!
0%
#172185000000
1!
1%
#172190000000
0!
0%
#172195000000
1!
1%
#172200000000
0!
0%
#172205000000
1!
1%
#172210000000
0!
0%
#172215000000
1!
1%
#172220000000
0!
0%
#172225000000
1!
1%
#172230000000
0!
0%
#172235000000
1!
1%
#172240000000
0!
0%
#172245000000
1!
1%
#172250000000
0!
0%
#172255000000
1!
1%
#172260000000
0!
0%
#172265000000
1!
1%
#172270000000
0!
0%
#172275000000
1!
1%
#172280000000
0!
0%
#172285000000
1!
1%
#172290000000
0!
0%
#172295000000
1!
1%
#172300000000
0!
0%
#172305000000
1!
1%
#172310000000
0!
0%
#172315000000
1!
1%
#172320000000
0!
0%
#172325000000
1!
1%
#172330000000
0!
0%
#172335000000
1!
1%
#172340000000
0!
0%
#172345000000
1!
1%
#172350000000
0!
0%
#172355000000
1!
1%
#172360000000
0!
0%
#172365000000
1!
1%
#172370000000
0!
0%
#172375000000
1!
1%
#172380000000
0!
0%
#172385000000
1!
1%
#172390000000
0!
0%
#172395000000
1!
1%
#172400000000
0!
0%
#172405000000
1!
1%
#172410000000
0!
0%
#172415000000
1!
1%
#172420000000
0!
0%
#172425000000
1!
1%
#172430000000
0!
0%
#172435000000
1!
1%
#172440000000
0!
0%
#172445000000
1!
1%
#172450000000
0!
0%
#172455000000
1!
1%
#172460000000
0!
0%
#172465000000
1!
1%
#172470000000
0!
0%
#172475000000
1!
1%
#172480000000
0!
0%
#172485000000
1!
1%
#172490000000
0!
0%
#172495000000
1!
1%
#172500000000
0!
0%
#172505000000
1!
1%
#172510000000
0!
0%
#172515000000
1!
1%
#172520000000
0!
0%
#172525000000
1!
1%
#172530000000
0!
0%
#172535000000
1!
1%
#172540000000
0!
0%
#172545000000
1!
1%
#172550000000
0!
0%
#172555000000
1!
1%
#172560000000
0!
0%
#172565000000
1!
1%
#172570000000
0!
0%
#172575000000
1!
1%
#172580000000
0!
0%
#172585000000
1!
1%
#172590000000
0!
0%
#172595000000
1!
1%
#172600000000
0!
0%
#172605000000
1!
1%
#172610000000
0!
0%
#172615000000
1!
1%
#172620000000
0!
0%
#172625000000
1!
1%
#172630000000
0!
0%
#172635000000
1!
1%
#172640000000
0!
0%
#172645000000
1!
1%
#172650000000
0!
0%
#172655000000
1!
1%
#172660000000
0!
0%
#172665000000
1!
1%
#172670000000
0!
0%
#172675000000
1!
1%
#172680000000
0!
0%
#172685000000
1!
1%
#172690000000
0!
0%
#172695000000
1!
1%
#172700000000
0!
0%
#172705000000
1!
1%
#172710000000
0!
0%
#172715000000
1!
1%
#172720000000
0!
0%
#172725000000
1!
1%
#172730000000
0!
0%
#172735000000
1!
1%
#172740000000
0!
0%
#172745000000
1!
1%
#172750000000
0!
0%
#172755000000
1!
1%
#172760000000
0!
0%
#172765000000
1!
1%
#172770000000
0!
0%
#172775000000
1!
1%
#172780000000
0!
0%
#172785000000
1!
1%
#172790000000
0!
0%
#172795000000
1!
1%
#172800000000
0!
0%
#172805000000
1!
1%
#172810000000
0!
0%
#172815000000
1!
1%
#172820000000
0!
0%
#172825000000
1!
1%
#172830000000
0!
0%
#172835000000
1!
1%
#172840000000
0!
0%
#172845000000
1!
1%
#172850000000
0!
0%
#172855000000
1!
1%
#172860000000
0!
0%
#172865000000
1!
1%
#172870000000
0!
0%
#172875000000
1!
1%
#172880000000
0!
0%
#172885000000
1!
1%
#172890000000
0!
0%
#172895000000
1!
1%
#172900000000
0!
0%
#172905000000
1!
1%
#172910000000
0!
0%
#172915000000
1!
1%
#172920000000
0!
0%
#172925000000
1!
1%
#172930000000
0!
0%
#172935000000
1!
1%
#172940000000
0!
0%
#172945000000
1!
1%
#172950000000
0!
0%
#172955000000
1!
1%
#172960000000
0!
0%
#172965000000
1!
1%
#172970000000
0!
0%
#172975000000
1!
1%
#172980000000
0!
0%
#172985000000
1!
1%
#172990000000
0!
0%
#172995000000
1!
1%
#173000000000
0!
0%
#173005000000
1!
1%
#173010000000
0!
0%
#173015000000
1!
1%
#173020000000
0!
0%
#173025000000
1!
1%
#173030000000
0!
0%
#173035000000
1!
1%
#173040000000
0!
0%
#173045000000
1!
1%
#173050000000
0!
0%
#173055000000
1!
1%
#173060000000
0!
0%
#173065000000
1!
1%
#173070000000
0!
0%
#173075000000
1!
1%
#173080000000
0!
0%
#173085000000
1!
1%
#173090000000
0!
0%
#173095000000
1!
1%
#173100000000
0!
0%
#173105000000
1!
1%
#173110000000
0!
0%
#173115000000
1!
1%
#173120000000
0!
0%
#173125000000
1!
1%
#173130000000
0!
0%
#173135000000
1!
1%
#173140000000
0!
0%
#173145000000
1!
1%
#173150000000
0!
0%
#173155000000
1!
1%
#173160000000
0!
0%
#173165000000
1!
1%
#173170000000
0!
0%
#173175000000
1!
1%
#173180000000
0!
0%
#173185000000
1!
1%
#173190000000
0!
0%
#173195000000
1!
1%
#173200000000
0!
0%
#173205000000
1!
1%
#173210000000
0!
0%
#173215000000
1!
1%
#173220000000
0!
0%
#173225000000
1!
1%
#173230000000
0!
0%
#173235000000
1!
1%
#173240000000
0!
0%
#173245000000
1!
1%
#173250000000
0!
0%
#173255000000
1!
1%
#173260000000
0!
0%
#173265000000
1!
1%
#173270000000
0!
0%
#173275000000
1!
1%
#173280000000
0!
0%
#173285000000
1!
1%
#173290000000
0!
0%
#173295000000
1!
1%
#173300000000
0!
0%
#173305000000
1!
1%
#173310000000
0!
0%
#173315000000
1!
1%
#173320000000
0!
0%
#173325000000
1!
1%
#173330000000
0!
0%
#173335000000
1!
1%
#173340000000
0!
0%
#173345000000
1!
1%
#173350000000
0!
0%
#173355000000
1!
1%
#173360000000
0!
0%
#173365000000
1!
1%
#173370000000
0!
0%
#173375000000
1!
1%
#173380000000
0!
0%
#173385000000
1!
1%
#173390000000
0!
0%
#173395000000
1!
1%
#173400000000
0!
0%
#173405000000
1!
1%
#173410000000
0!
0%
#173415000000
1!
1%
#173420000000
0!
0%
#173425000000
1!
1%
#173430000000
0!
0%
#173435000000
1!
1%
#173440000000
0!
0%
#173445000000
1!
1%
#173450000000
0!
0%
#173455000000
1!
1%
#173460000000
0!
0%
#173465000000
1!
1%
#173470000000
0!
0%
#173475000000
1!
1%
#173480000000
0!
0%
#173485000000
1!
1%
#173490000000
0!
0%
#173495000000
1!
1%
#173500000000
0!
0%
#173505000000
1!
1%
#173510000000
0!
0%
#173515000000
1!
1%
#173520000000
0!
0%
#173525000000
1!
1%
#173530000000
0!
0%
#173535000000
1!
1%
#173540000000
0!
0%
#173545000000
1!
1%
#173550000000
0!
0%
#173555000000
1!
1%
#173560000000
0!
0%
#173565000000
1!
1%
#173570000000
0!
0%
#173575000000
1!
1%
#173580000000
0!
0%
#173585000000
1!
1%
#173590000000
0!
0%
#173595000000
1!
1%
#173600000000
0!
0%
#173605000000
1!
1%
#173610000000
0!
0%
#173615000000
1!
1%
#173620000000
0!
0%
#173625000000
1!
1%
#173630000000
0!
0%
#173635000000
1!
1%
#173640000000
0!
0%
#173645000000
1!
1%
#173650000000
0!
0%
#173655000000
1!
1%
#173660000000
0!
0%
#173665000000
1!
1%
#173670000000
0!
0%
#173675000000
1!
1%
#173680000000
0!
0%
#173685000000
1!
1%
#173690000000
0!
0%
#173695000000
1!
1%
#173700000000
0!
0%
#173705000000
1!
1%
#173710000000
0!
0%
#173715000000
1!
1%
#173720000000
0!
0%
#173725000000
1!
1%
#173730000000
0!
0%
#173735000000
1!
1%
#173740000000
0!
0%
#173745000000
1!
1%
#173750000000
0!
0%
#173755000000
1!
1%
#173760000000
0!
0%
#173765000000
1!
1%
#173770000000
0!
0%
#173775000000
1!
1%
#173780000000
0!
0%
#173785000000
1!
1%
#173790000000
0!
0%
#173795000000
1!
1%
#173800000000
0!
0%
#173805000000
1!
1%
#173810000000
0!
0%
#173815000000
1!
1%
#173820000000
0!
0%
#173825000000
1!
1%
#173830000000
0!
0%
#173835000000
1!
1%
#173840000000
0!
0%
#173845000000
1!
1%
#173850000000
0!
0%
#173855000000
1!
1%
#173860000000
0!
0%
#173865000000
1!
1%
#173870000000
0!
0%
#173875000000
1!
1%
#173880000000
0!
0%
#173885000000
1!
1%
#173890000000
0!
0%
#173895000000
1!
1%
#173900000000
0!
0%
#173905000000
1!
1%
#173910000000
0!
0%
#173915000000
1!
1%
#173920000000
0!
0%
#173925000000
1!
1%
#173930000000
0!
0%
#173935000000
1!
1%
#173940000000
0!
0%
#173945000000
1!
1%
#173950000000
0!
0%
#173955000000
1!
1%
#173960000000
0!
0%
#173965000000
1!
1%
#173970000000
0!
0%
#173975000000
1!
1%
#173980000000
0!
0%
#173985000000
1!
1%
#173990000000
0!
0%
#173995000000
1!
1%
#174000000000
0!
0%
#174005000000
1!
1%
#174010000000
0!
0%
#174015000000
1!
1%
#174020000000
0!
0%
#174025000000
1!
1%
#174030000000
0!
0%
#174035000000
1!
1%
#174040000000
0!
0%
#174045000000
1!
1%
#174050000000
0!
0%
#174055000000
1!
1%
#174060000000
0!
0%
#174065000000
1!
1%
#174070000000
0!
0%
#174075000000
1!
1%
#174080000000
0!
0%
#174085000000
1!
1%
#174090000000
0!
0%
#174095000000
1!
1%
#174100000000
0!
0%
#174105000000
1!
1%
#174110000000
0!
0%
#174115000000
1!
1%
#174120000000
0!
0%
#174125000000
1!
1%
#174130000000
0!
0%
#174135000000
1!
1%
#174140000000
0!
0%
#174145000000
1!
1%
#174150000000
0!
0%
#174155000000
1!
1%
#174160000000
0!
0%
#174165000000
1!
1%
#174170000000
0!
0%
#174175000000
1!
1%
#174180000000
0!
0%
#174185000000
1!
1%
#174190000000
0!
0%
#174195000000
1!
1%
#174200000000
0!
0%
#174205000000
1!
1%
#174210000000
0!
0%
#174215000000
1!
1%
#174220000000
0!
0%
#174225000000
1!
1%
#174230000000
0!
0%
#174235000000
1!
1%
#174240000000
0!
0%
#174245000000
1!
1%
#174250000000
0!
0%
#174255000000
1!
1%
#174260000000
0!
0%
#174265000000
1!
1%
#174270000000
0!
0%
#174275000000
1!
1%
#174280000000
0!
0%
#174285000000
1!
1%
#174290000000
0!
0%
#174295000000
1!
1%
#174300000000
0!
0%
#174305000000
1!
1%
#174310000000
0!
0%
#174315000000
1!
1%
#174320000000
0!
0%
#174325000000
1!
1%
#174330000000
0!
0%
#174335000000
1!
1%
#174340000000
0!
0%
#174345000000
1!
1%
#174350000000
0!
0%
#174355000000
1!
1%
#174360000000
0!
0%
#174365000000
1!
1%
#174370000000
0!
0%
#174375000000
1!
1%
#174380000000
0!
0%
#174385000000
1!
1%
#174390000000
0!
0%
#174395000000
1!
1%
#174400000000
0!
0%
#174405000000
1!
1%
#174410000000
0!
0%
#174415000000
1!
1%
#174420000000
0!
0%
#174425000000
1!
1%
#174430000000
0!
0%
#174435000000
1!
1%
#174440000000
0!
0%
#174445000000
1!
1%
#174450000000
0!
0%
#174455000000
1!
1%
#174460000000
0!
0%
#174465000000
1!
1%
#174470000000
0!
0%
#174475000000
1!
1%
#174480000000
0!
0%
#174485000000
1!
1%
#174490000000
0!
0%
#174495000000
1!
1%
#174500000000
0!
0%
#174505000000
1!
1%
#174510000000
0!
0%
#174515000000
1!
1%
#174520000000
0!
0%
#174525000000
1!
1%
#174530000000
0!
0%
#174535000000
1!
1%
#174540000000
0!
0%
#174545000000
1!
1%
#174550000000
0!
0%
#174555000000
1!
1%
#174560000000
0!
0%
#174565000000
1!
1%
#174570000000
0!
0%
#174575000000
1!
1%
#174580000000
0!
0%
#174585000000
1!
1%
#174590000000
0!
0%
#174595000000
1!
1%
#174600000000
0!
0%
#174605000000
1!
1%
#174610000000
0!
0%
#174615000000
1!
1%
#174620000000
0!
0%
#174625000000
1!
1%
#174630000000
0!
0%
#174635000000
1!
1%
#174640000000
0!
0%
#174645000000
1!
1%
#174650000000
0!
0%
#174655000000
1!
1%
#174660000000
0!
0%
#174665000000
1!
1%
#174670000000
0!
0%
#174675000000
1!
1%
#174680000000
0!
0%
#174685000000
1!
1%
#174690000000
0!
0%
#174695000000
1!
1%
#174700000000
0!
0%
#174705000000
1!
1%
#174710000000
0!
0%
#174715000000
1!
1%
#174720000000
0!
0%
#174725000000
1!
1%
#174730000000
0!
0%
#174735000000
1!
1%
#174740000000
0!
0%
#174745000000
1!
1%
#174750000000
0!
0%
#174755000000
1!
1%
#174760000000
0!
0%
#174765000000
1!
1%
#174770000000
0!
0%
#174775000000
1!
1%
#174780000000
0!
0%
#174785000000
1!
1%
#174790000000
0!
0%
#174795000000
1!
1%
#174800000000
0!
0%
#174805000000
1!
1%
#174810000000
0!
0%
#174815000000
1!
1%
#174820000000
0!
0%
#174825000000
1!
1%
#174830000000
0!
0%
#174835000000
1!
1%
#174840000000
0!
0%
#174845000000
1!
1%
#174850000000
0!
0%
#174855000000
1!
1%
#174860000000
0!
0%
#174865000000
1!
1%
#174870000000
0!
0%
#174875000000
1!
1%
#174880000000
0!
0%
#174885000000
1!
1%
#174890000000
0!
0%
#174895000000
1!
1%
#174900000000
0!
0%
#174905000000
1!
1%
#174910000000
0!
0%
#174915000000
1!
1%
#174920000000
0!
0%
#174925000000
1!
1%
#174930000000
0!
0%
#174935000000
1!
1%
#174940000000
0!
0%
#174945000000
1!
1%
#174950000000
0!
0%
#174955000000
1!
1%
#174960000000
0!
0%
#174965000000
1!
1%
#174970000000
0!
0%
#174975000000
1!
1%
#174980000000
0!
0%
#174985000000
1!
1%
#174990000000
0!
0%
#174995000000
1!
1%
#175000000000
0!
0%
#175005000000
1!
1%
#175010000000
0!
0%
#175015000000
1!
1%
#175020000000
0!
0%
#175025000000
1!
1%
#175030000000
0!
0%
#175035000000
1!
1%
#175040000000
0!
0%
#175045000000
1!
1%
#175050000000
0!
0%
#175055000000
1!
1%
#175060000000
0!
0%
#175065000000
1!
1%
#175070000000
0!
0%
#175075000000
1!
1%
#175080000000
0!
0%
#175085000000
1!
1%
#175090000000
0!
0%
#175095000000
1!
1%
#175100000000
0!
0%
#175105000000
1!
1%
#175110000000
0!
0%
#175115000000
1!
1%
#175120000000
0!
0%
#175125000000
1!
1%
#175130000000
0!
0%
#175135000000
1!
1%
#175140000000
0!
0%
#175145000000
1!
1%
#175150000000
0!
0%
#175155000000
1!
1%
#175160000000
0!
0%
#175165000000
1!
1%
#175170000000
0!
0%
#175175000000
1!
1%
#175180000000
0!
0%
#175185000000
1!
1%
#175190000000
0!
0%
#175195000000
1!
1%
#175200000000
0!
0%
#175205000000
1!
1%
#175210000000
0!
0%
#175215000000
1!
1%
#175220000000
0!
0%
#175225000000
1!
1%
#175230000000
0!
0%
#175235000000
1!
1%
#175240000000
0!
0%
#175245000000
1!
1%
#175250000000
0!
0%
#175255000000
1!
1%
#175260000000
0!
0%
#175265000000
1!
1%
#175270000000
0!
0%
#175275000000
1!
1%
#175280000000
0!
0%
#175285000000
1!
1%
#175290000000
0!
0%
#175295000000
1!
1%
#175300000000
0!
0%
#175305000000
1!
1%
#175310000000
0!
0%
#175315000000
1!
1%
#175320000000
0!
0%
#175325000000
1!
1%
#175330000000
0!
0%
#175335000000
1!
1%
#175340000000
0!
0%
#175345000000
1!
1%
#175350000000
0!
0%
#175355000000
1!
1%
#175360000000
0!
0%
#175365000000
1!
1%
#175370000000
0!
0%
#175375000000
1!
1%
#175380000000
0!
0%
#175385000000
1!
1%
#175390000000
0!
0%
#175395000000
1!
1%
#175400000000
0!
0%
#175405000000
1!
1%
#175410000000
0!
0%
#175415000000
1!
1%
#175420000000
0!
0%
#175425000000
1!
1%
#175430000000
0!
0%
#175435000000
1!
1%
#175440000000
0!
0%
#175445000000
1!
1%
#175450000000
0!
0%
#175455000000
1!
1%
#175460000000
0!
0%
#175465000000
1!
1%
#175470000000
0!
0%
#175475000000
1!
1%
#175480000000
0!
0%
#175485000000
1!
1%
#175490000000
0!
0%
#175495000000
1!
1%
#175500000000
0!
0%
#175505000000
1!
1%
#175510000000
0!
0%
#175515000000
1!
1%
#175520000000
0!
0%
#175525000000
1!
1%
#175530000000
0!
0%
#175535000000
1!
1%
#175540000000
0!
0%
#175545000000
1!
1%
#175550000000
0!
0%
#175555000000
1!
1%
#175560000000
0!
0%
#175565000000
1!
1%
#175570000000
0!
0%
#175575000000
1!
1%
#175580000000
0!
0%
#175585000000
1!
1%
#175590000000
0!
0%
#175595000000
1!
1%
#175600000000
0!
0%
#175605000000
1!
1%
#175610000000
0!
0%
#175615000000
1!
1%
#175620000000
0!
0%
#175625000000
1!
1%
#175630000000
0!
0%
#175635000000
1!
1%
#175640000000
0!
0%
#175645000000
1!
1%
#175650000000
0!
0%
#175655000000
1!
1%
#175660000000
0!
0%
#175665000000
1!
1%
#175670000000
0!
0%
#175675000000
1!
1%
#175680000000
0!
0%
#175685000000
1!
1%
#175690000000
0!
0%
#175695000000
1!
1%
#175700000000
0!
0%
#175705000000
1!
1%
#175710000000
0!
0%
#175715000000
1!
1%
#175720000000
0!
0%
#175725000000
1!
1%
#175730000000
0!
0%
#175735000000
1!
1%
#175740000000
0!
0%
#175745000000
1!
1%
#175750000000
0!
0%
#175755000000
1!
1%
#175760000000
0!
0%
#175765000000
1!
1%
#175770000000
0!
0%
#175775000000
1!
1%
#175780000000
0!
0%
#175785000000
1!
1%
#175790000000
0!
0%
#175795000000
1!
1%
#175800000000
0!
0%
#175805000000
1!
1%
#175810000000
0!
0%
#175815000000
1!
1%
#175820000000
0!
0%
#175825000000
1!
1%
#175830000000
0!
0%
#175835000000
1!
1%
#175840000000
0!
0%
#175845000000
1!
1%
#175850000000
0!
0%
#175855000000
1!
1%
#175860000000
0!
0%
#175865000000
1!
1%
#175870000000
0!
0%
#175875000000
1!
1%
#175880000000
0!
0%
#175885000000
1!
1%
#175890000000
0!
0%
#175895000000
1!
1%
#175900000000
0!
0%
#175905000000
1!
1%
#175910000000
0!
0%
#175915000000
1!
1%
#175920000000
0!
0%
#175925000000
1!
1%
#175930000000
0!
0%
#175935000000
1!
1%
#175940000000
0!
0%
#175945000000
1!
1%
#175950000000
0!
0%
#175955000000
1!
1%
#175960000000
0!
0%
#175965000000
1!
1%
#175970000000
0!
0%
#175975000000
1!
1%
#175980000000
0!
0%
#175985000000
1!
1%
#175990000000
0!
0%
#175995000000
1!
1%
#176000000000
0!
0%
#176005000000
1!
1%
#176010000000
0!
0%
#176015000000
1!
1%
#176020000000
0!
0%
#176025000000
1!
1%
#176030000000
0!
0%
#176035000000
1!
1%
#176040000000
0!
0%
#176045000000
1!
1%
#176050000000
0!
0%
#176055000000
1!
1%
#176060000000
0!
0%
#176065000000
1!
1%
#176070000000
0!
0%
#176075000000
1!
1%
#176080000000
0!
0%
#176085000000
1!
1%
#176090000000
0!
0%
#176095000000
1!
1%
#176100000000
0!
0%
#176105000000
1!
1%
#176110000000
0!
0%
#176115000000
1!
1%
#176120000000
0!
0%
#176125000000
1!
1%
#176130000000
0!
0%
#176135000000
1!
1%
#176140000000
0!
0%
#176145000000
1!
1%
#176150000000
0!
0%
#176155000000
1!
1%
#176160000000
0!
0%
#176165000000
1!
1%
#176170000000
0!
0%
#176175000000
1!
1%
#176180000000
0!
0%
#176185000000
1!
1%
#176190000000
0!
0%
#176195000000
1!
1%
#176200000000
0!
0%
#176205000000
1!
1%
#176210000000
0!
0%
#176215000000
1!
1%
#176220000000
0!
0%
#176225000000
1!
1%
#176230000000
0!
0%
#176235000000
1!
1%
#176240000000
0!
0%
#176245000000
1!
1%
#176250000000
0!
0%
#176255000000
1!
1%
#176260000000
0!
0%
#176265000000
1!
1%
#176270000000
0!
0%
#176275000000
1!
1%
#176280000000
0!
0%
#176285000000
1!
1%
#176290000000
0!
0%
#176295000000
1!
1%
#176300000000
0!
0%
#176305000000
1!
1%
#176310000000
0!
0%
#176315000000
1!
1%
#176320000000
0!
0%
#176325000000
1!
1%
#176330000000
0!
0%
#176335000000
1!
1%
#176340000000
0!
0%
#176345000000
1!
1%
#176350000000
0!
0%
#176355000000
1!
1%
#176360000000
0!
0%
#176365000000
1!
1%
#176370000000
0!
0%
#176375000000
1!
1%
#176380000000
0!
0%
#176385000000
1!
1%
#176390000000
0!
0%
#176395000000
1!
1%
#176400000000
0!
0%
#176405000000
1!
1%
#176410000000
0!
0%
#176415000000
1!
1%
#176420000000
0!
0%
#176425000000
1!
1%
#176430000000
0!
0%
#176435000000
1!
1%
#176440000000
0!
0%
#176445000000
1!
1%
#176450000000
0!
0%
#176455000000
1!
1%
#176460000000
0!
0%
#176465000000
1!
1%
#176470000000
0!
0%
#176475000000
1!
1%
#176480000000
0!
0%
#176485000000
1!
1%
#176490000000
0!
0%
#176495000000
1!
1%
#176500000000
0!
0%
#176505000000
1!
1%
#176510000000
0!
0%
#176515000000
1!
1%
#176520000000
0!
0%
#176525000000
1!
1%
#176530000000
0!
0%
#176535000000
1!
1%
#176540000000
0!
0%
#176545000000
1!
1%
#176550000000
0!
0%
#176555000000
1!
1%
#176560000000
0!
0%
#176565000000
1!
1%
#176570000000
0!
0%
#176575000000
1!
1%
#176580000000
0!
0%
#176585000000
1!
1%
#176590000000
0!
0%
#176595000000
1!
1%
#176600000000
0!
0%
#176605000000
1!
1%
#176610000000
0!
0%
#176615000000
1!
1%
#176620000000
0!
0%
#176625000000
1!
1%
#176630000000
0!
0%
#176635000000
1!
1%
#176640000000
0!
0%
#176645000000
1!
1%
#176650000000
0!
0%
#176655000000
1!
1%
#176660000000
0!
0%
#176665000000
1!
1%
#176670000000
0!
0%
#176675000000
1!
1%
#176680000000
0!
0%
#176685000000
1!
1%
#176690000000
0!
0%
#176695000000
1!
1%
#176700000000
0!
0%
#176705000000
1!
1%
#176710000000
0!
0%
#176715000000
1!
1%
#176720000000
0!
0%
#176725000000
1!
1%
#176730000000
0!
0%
#176735000000
1!
1%
#176740000000
0!
0%
#176745000000
1!
1%
#176750000000
0!
0%
#176755000000
1!
1%
#176760000000
0!
0%
#176765000000
1!
1%
#176770000000
0!
0%
#176775000000
1!
1%
#176780000000
0!
0%
#176785000000
1!
1%
#176790000000
0!
0%
#176795000000
1!
1%
#176800000000
0!
0%
#176805000000
1!
1%
#176810000000
0!
0%
#176815000000
1!
1%
#176820000000
0!
0%
#176825000000
1!
1%
#176830000000
0!
0%
#176835000000
1!
1%
#176840000000
0!
0%
#176845000000
1!
1%
#176850000000
0!
0%
#176855000000
1!
1%
#176860000000
0!
0%
#176865000000
1!
1%
#176870000000
0!
0%
#176875000000
1!
1%
#176880000000
0!
0%
#176885000000
1!
1%
#176890000000
0!
0%
#176895000000
1!
1%
#176900000000
0!
0%
#176905000000
1!
1%
#176910000000
0!
0%
#176915000000
1!
1%
#176920000000
0!
0%
#176925000000
1!
1%
#176930000000
0!
0%
#176935000000
1!
1%
#176940000000
0!
0%
#176945000000
1!
1%
#176950000000
0!
0%
#176955000000
1!
1%
#176960000000
0!
0%
#176965000000
1!
1%
#176970000000
0!
0%
#176975000000
1!
1%
#176980000000
0!
0%
#176985000000
1!
1%
#176990000000
0!
0%
#176995000000
1!
1%
#177000000000
0!
0%
#177005000000
1!
1%
#177010000000
0!
0%
#177015000000
1!
1%
#177020000000
0!
0%
#177025000000
1!
1%
#177030000000
0!
0%
#177035000000
1!
1%
#177040000000
0!
0%
#177045000000
1!
1%
#177050000000
0!
0%
#177055000000
1!
1%
#177060000000
0!
0%
#177065000000
1!
1%
#177070000000
0!
0%
#177075000000
1!
1%
#177080000000
0!
0%
#177085000000
1!
1%
#177090000000
0!
0%
#177095000000
1!
1%
#177100000000
0!
0%
#177105000000
1!
1%
#177110000000
0!
0%
#177115000000
1!
1%
#177120000000
0!
0%
#177125000000
1!
1%
#177130000000
0!
0%
#177135000000
1!
1%
#177140000000
0!
0%
#177145000000
1!
1%
#177150000000
0!
0%
#177155000000
1!
1%
#177160000000
0!
0%
#177165000000
1!
1%
#177170000000
0!
0%
#177175000000
1!
1%
#177180000000
0!
0%
#177185000000
1!
1%
#177190000000
0!
0%
#177195000000
1!
1%
#177200000000
0!
0%
#177205000000
1!
1%
#177210000000
0!
0%
#177215000000
1!
1%
#177220000000
0!
0%
#177225000000
1!
1%
#177230000000
0!
0%
#177235000000
1!
1%
#177240000000
0!
0%
#177245000000
1!
1%
#177250000000
0!
0%
#177255000000
1!
1%
#177260000000
0!
0%
#177265000000
1!
1%
#177270000000
0!
0%
#177275000000
1!
1%
#177280000000
0!
0%
#177285000000
1!
1%
#177290000000
0!
0%
#177295000000
1!
1%
#177300000000
0!
0%
#177305000000
1!
1%
#177310000000
0!
0%
#177315000000
1!
1%
#177320000000
0!
0%
#177325000000
1!
1%
#177330000000
0!
0%
#177335000000
1!
1%
#177340000000
0!
0%
#177345000000
1!
1%
#177350000000
0!
0%
#177355000000
1!
1%
#177360000000
0!
0%
#177365000000
1!
1%
#177370000000
0!
0%
#177375000000
1!
1%
#177380000000
0!
0%
#177385000000
1!
1%
#177390000000
0!
0%
#177395000000
1!
1%
#177400000000
0!
0%
#177405000000
1!
1%
#177410000000
0!
0%
#177415000000
1!
1%
#177420000000
0!
0%
#177425000000
1!
1%
#177430000000
0!
0%
#177435000000
1!
1%
#177440000000
0!
0%
#177445000000
1!
1%
#177450000000
0!
0%
#177455000000
1!
1%
#177460000000
0!
0%
#177465000000
1!
1%
#177470000000
0!
0%
#177475000000
1!
1%
#177480000000
0!
0%
#177485000000
1!
1%
#177490000000
0!
0%
#177495000000
1!
1%
#177500000000
0!
0%
#177505000000
1!
1%
#177510000000
0!
0%
#177515000000
1!
1%
#177520000000
0!
0%
#177525000000
1!
1%
#177530000000
0!
0%
#177535000000
1!
1%
#177540000000
0!
0%
#177545000000
1!
1%
#177550000000
0!
0%
#177555000000
1!
1%
#177560000000
0!
0%
#177565000000
1!
1%
#177570000000
0!
0%
#177575000000
1!
1%
#177580000000
0!
0%
#177585000000
1!
1%
#177590000000
0!
0%
#177595000000
1!
1%
#177600000000
0!
0%
#177605000000
1!
1%
#177610000000
0!
0%
#177615000000
1!
1%
#177620000000
0!
0%
#177625000000
1!
1%
#177630000000
0!
0%
#177635000000
1!
1%
#177640000000
0!
0%
#177645000000
1!
1%
#177650000000
0!
0%
#177655000000
1!
1%
#177660000000
0!
0%
#177665000000
1!
1%
#177670000000
0!
0%
#177675000000
1!
1%
#177680000000
0!
0%
#177685000000
1!
1%
#177690000000
0!
0%
#177695000000
1!
1%
#177700000000
0!
0%
#177705000000
1!
1%
#177710000000
0!
0%
#177715000000
1!
1%
#177720000000
0!
0%
#177725000000
1!
1%
#177730000000
0!
0%
#177735000000
1!
1%
#177740000000
0!
0%
#177745000000
1!
1%
#177750000000
0!
0%
#177755000000
1!
1%
#177760000000
0!
0%
#177765000000
1!
1%
#177770000000
0!
0%
#177775000000
1!
1%
#177780000000
0!
0%
#177785000000
1!
1%
#177790000000
0!
0%
#177795000000
1!
1%
#177800000000
0!
0%
#177805000000
1!
1%
#177810000000
0!
0%
#177815000000
1!
1%
#177820000000
0!
0%
#177825000000
1!
1%
#177830000000
0!
0%
#177835000000
1!
1%
#177840000000
0!
0%
#177845000000
1!
1%
#177850000000
0!
0%
#177855000000
1!
1%
#177860000000
0!
0%
#177865000000
1!
1%
#177870000000
0!
0%
#177875000000
1!
1%
#177880000000
0!
0%
#177885000000
1!
1%
#177890000000
0!
0%
#177895000000
1!
1%
#177900000000
0!
0%
#177905000000
1!
1%
#177910000000
0!
0%
#177915000000
1!
1%
#177920000000
0!
0%
#177925000000
1!
1%
#177930000000
0!
0%
#177935000000
1!
1%
#177940000000
0!
0%
#177945000000
1!
1%
#177950000000
0!
0%
#177955000000
1!
1%
#177960000000
0!
0%
#177965000000
1!
1%
#177970000000
0!
0%
#177975000000
1!
1%
#177980000000
0!
0%
#177985000000
1!
1%
#177990000000
0!
0%
#177995000000
1!
1%
#178000000000
0!
0%
#178005000000
1!
1%
#178010000000
0!
0%
#178015000000
1!
1%
#178020000000
0!
0%
#178025000000
1!
1%
#178030000000
0!
0%
#178035000000
1!
1%
#178040000000
0!
0%
#178045000000
1!
1%
#178050000000
0!
0%
#178055000000
1!
1%
#178060000000
0!
0%
#178065000000
1!
1%
#178070000000
0!
0%
#178075000000
1!
1%
#178080000000
0!
0%
#178085000000
1!
1%
#178090000000
0!
0%
#178095000000
1!
1%
#178100000000
0!
0%
#178105000000
1!
1%
#178110000000
0!
0%
#178115000000
1!
1%
#178120000000
0!
0%
#178125000000
1!
1%
#178130000000
0!
0%
#178135000000
1!
1%
#178140000000
0!
0%
#178145000000
1!
1%
#178150000000
0!
0%
#178155000000
1!
1%
#178160000000
0!
0%
#178165000000
1!
1%
#178170000000
0!
0%
#178175000000
1!
1%
#178180000000
0!
0%
#178185000000
1!
1%
#178190000000
0!
0%
#178195000000
1!
1%
#178200000000
0!
0%
#178205000000
1!
1%
#178210000000
0!
0%
#178215000000
1!
1%
#178220000000
0!
0%
#178225000000
1!
1%
#178230000000
0!
0%
#178235000000
1!
1%
#178240000000
0!
0%
#178245000000
1!
1%
#178250000000
0!
0%
#178255000000
1!
1%
#178260000000
0!
0%
#178265000000
1!
1%
#178270000000
0!
0%
#178275000000
1!
1%
#178280000000
0!
0%
#178285000000
1!
1%
#178290000000
0!
0%
#178295000000
1!
1%
#178300000000
0!
0%
#178305000000
1!
1%
#178310000000
0!
0%
#178315000000
1!
1%
#178320000000
0!
0%
#178325000000
1!
1%
#178330000000
0!
0%
#178335000000
1!
1%
#178340000000
0!
0%
#178345000000
1!
1%
#178350000000
0!
0%
#178355000000
1!
1%
#178360000000
0!
0%
#178365000000
1!
1%
#178370000000
0!
0%
#178375000000
1!
1%
#178380000000
0!
0%
#178385000000
1!
1%
#178390000000
0!
0%
#178395000000
1!
1%
#178400000000
0!
0%
#178405000000
1!
1%
#178410000000
0!
0%
#178415000000
1!
1%
#178420000000
0!
0%
#178425000000
1!
1%
#178430000000
0!
0%
#178435000000
1!
1%
#178440000000
0!
0%
#178445000000
1!
1%
#178450000000
0!
0%
#178455000000
1!
1%
#178460000000
0!
0%
#178465000000
1!
1%
#178470000000
0!
0%
#178475000000
1!
1%
#178480000000
0!
0%
#178485000000
1!
1%
#178490000000
0!
0%
#178495000000
1!
1%
#178500000000
0!
0%
#178505000000
1!
1%
#178510000000
0!
0%
#178515000000
1!
1%
#178520000000
0!
0%
#178525000000
1!
1%
#178530000000
0!
0%
#178535000000
1!
1%
#178540000000
0!
0%
#178545000000
1!
1%
#178550000000
0!
0%
#178555000000
1!
1%
#178560000000
0!
0%
#178565000000
1!
1%
#178570000000
0!
0%
#178575000000
1!
1%
#178580000000
0!
0%
#178585000000
1!
1%
#178590000000
0!
0%
#178595000000
1!
1%
#178600000000
0!
0%
#178605000000
1!
1%
#178610000000
0!
0%
#178615000000
1!
1%
#178620000000
0!
0%
#178625000000
1!
1%
#178630000000
0!
0%
#178635000000
1!
1%
#178640000000
0!
0%
#178645000000
1!
1%
#178650000000
0!
0%
#178655000000
1!
1%
#178660000000
0!
0%
#178665000000
1!
1%
#178670000000
0!
0%
#178675000000
1!
1%
#178680000000
0!
0%
#178685000000
1!
1%
#178690000000
0!
0%
#178695000000
1!
1%
#178700000000
0!
0%
#178705000000
1!
1%
#178710000000
0!
0%
#178715000000
1!
1%
#178720000000
0!
0%
#178725000000
1!
1%
#178730000000
0!
0%
#178735000000
1!
1%
#178740000000
0!
0%
#178745000000
1!
1%
#178750000000
0!
0%
#178755000000
1!
1%
#178760000000
0!
0%
#178765000000
1!
1%
#178770000000
0!
0%
#178775000000
1!
1%
#178780000000
0!
0%
#178785000000
1!
1%
#178790000000
0!
0%
#178795000000
1!
1%
#178800000000
0!
0%
#178805000000
1!
1%
#178810000000
0!
0%
#178815000000
1!
1%
#178820000000
0!
0%
#178825000000
1!
1%
#178830000000
0!
0%
#178835000000
1!
1%
#178840000000
0!
0%
#178845000000
1!
1%
#178850000000
0!
0%
#178855000000
1!
1%
#178860000000
0!
0%
#178865000000
1!
1%
#178870000000
0!
0%
#178875000000
1!
1%
#178880000000
0!
0%
#178885000000
1!
1%
#178890000000
0!
0%
#178895000000
1!
1%
#178900000000
0!
0%
#178905000000
1!
1%
#178910000000
0!
0%
#178915000000
1!
1%
#178920000000
0!
0%
#178925000000
1!
1%
#178930000000
0!
0%
#178935000000
1!
1%
#178940000000
0!
0%
#178945000000
1!
1%
#178950000000
0!
0%
#178955000000
1!
1%
#178960000000
0!
0%
#178965000000
1!
1%
#178970000000
0!
0%
#178975000000
1!
1%
#178980000000
0!
0%
#178985000000
1!
1%
#178990000000
0!
0%
#178995000000
1!
1%
#179000000000
0!
0%
#179005000000
1!
1%
#179010000000
0!
0%
#179015000000
1!
1%
#179020000000
0!
0%
#179025000000
1!
1%
#179030000000
0!
0%
#179035000000
1!
1%
#179040000000
0!
0%
#179045000000
1!
1%
#179050000000
0!
0%
#179055000000
1!
1%
#179060000000
0!
0%
#179065000000
1!
1%
#179070000000
0!
0%
#179075000000
1!
1%
#179080000000
0!
0%
#179085000000
1!
1%
#179090000000
0!
0%
#179095000000
1!
1%
#179100000000
0!
0%
#179105000000
1!
1%
#179110000000
0!
0%
#179115000000
1!
1%
#179120000000
0!
0%
#179125000000
1!
1%
#179130000000
0!
0%
#179135000000
1!
1%
#179140000000
0!
0%
#179145000000
1!
1%
#179150000000
0!
0%
#179155000000
1!
1%
#179160000000
0!
0%
#179165000000
1!
1%
#179170000000
0!
0%
#179175000000
1!
1%
#179180000000
0!
0%
#179185000000
1!
1%
#179190000000
0!
0%
#179195000000
1!
1%
#179200000000
0!
0%
#179205000000
1!
1%
#179210000000
0!
0%
#179215000000
1!
1%
#179220000000
0!
0%
#179225000000
1!
1%
#179230000000
0!
0%
#179235000000
1!
1%
#179240000000
0!
0%
#179245000000
1!
1%
#179250000000
0!
0%
#179255000000
1!
1%
#179260000000
0!
0%
#179265000000
1!
1%
#179270000000
0!
0%
#179275000000
1!
1%
#179280000000
0!
0%
#179285000000
1!
1%
#179290000000
0!
0%
#179295000000
1!
1%
#179300000000
0!
0%
#179305000000
1!
1%
#179310000000
0!
0%
#179315000000
1!
1%
#179320000000
0!
0%
#179325000000
1!
1%
#179330000000
0!
0%
#179335000000
1!
1%
#179340000000
0!
0%
#179345000000
1!
1%
#179350000000
0!
0%
#179355000000
1!
1%
#179360000000
0!
0%
#179365000000
1!
1%
#179370000000
0!
0%
#179375000000
1!
1%
#179380000000
0!
0%
#179385000000
1!
1%
#179390000000
0!
0%
#179395000000
1!
1%
#179400000000
0!
0%
#179405000000
1!
1%
#179410000000
0!
0%
#179415000000
1!
1%
#179420000000
0!
0%
#179425000000
1!
1%
#179430000000
0!
0%
#179435000000
1!
1%
#179440000000
0!
0%
#179445000000
1!
1%
#179450000000
0!
0%
#179455000000
1!
1%
#179460000000
0!
0%
#179465000000
1!
1%
#179470000000
0!
0%
#179475000000
1!
1%
#179480000000
0!
0%
#179485000000
1!
1%
#179490000000
0!
0%
#179495000000
1!
1%
#179500000000
0!
0%
#179505000000
1!
1%
#179510000000
0!
0%
#179515000000
1!
1%
#179520000000
0!
0%
#179525000000
1!
1%
#179530000000
0!
0%
#179535000000
1!
1%
#179540000000
0!
0%
#179545000000
1!
1%
#179550000000
0!
0%
#179555000000
1!
1%
#179560000000
0!
0%
#179565000000
1!
1%
#179570000000
0!
0%
#179575000000
1!
1%
#179580000000
0!
0%
#179585000000
1!
1%
#179590000000
0!
0%
#179595000000
1!
1%
#179600000000
0!
0%
#179605000000
1!
1%
#179610000000
0!
0%
#179615000000
1!
1%
#179620000000
0!
0%
#179625000000
1!
1%
#179630000000
0!
0%
#179635000000
1!
1%
#179640000000
0!
0%
#179645000000
1!
1%
#179650000000
0!
0%
#179655000000
1!
1%
#179660000000
0!
0%
#179665000000
1!
1%
#179670000000
0!
0%
#179675000000
1!
1%
#179680000000
0!
0%
#179685000000
1!
1%
#179690000000
0!
0%
#179695000000
1!
1%
#179700000000
0!
0%
#179705000000
1!
1%
#179710000000
0!
0%
#179715000000
1!
1%
#179720000000
0!
0%
#179725000000
1!
1%
#179730000000
0!
0%
#179735000000
1!
1%
#179740000000
0!
0%
#179745000000
1!
1%
#179750000000
0!
0%
#179755000000
1!
1%
#179760000000
0!
0%
#179765000000
1!
1%
#179770000000
0!
0%
#179775000000
1!
1%
#179780000000
0!
0%
#179785000000
1!
1%
#179790000000
0!
0%
#179795000000
1!
1%
#179800000000
0!
0%
#179805000000
1!
1%
#179810000000
0!
0%
#179815000000
1!
1%
#179820000000
0!
0%
#179825000000
1!
1%
#179830000000
0!
0%
#179835000000
1!
1%
#179840000000
0!
0%
#179845000000
1!
1%
#179850000000
0!
0%
#179855000000
1!
1%
#179860000000
0!
0%
#179865000000
1!
1%
#179870000000
0!
0%
#179875000000
1!
1%
#179880000000
0!
0%
#179885000000
1!
1%
#179890000000
0!
0%
#179895000000
1!
1%
#179900000000
0!
0%
#179905000000
1!
1%
#179910000000
0!
0%
#179915000000
1!
1%
#179920000000
0!
0%
#179925000000
1!
1%
#179930000000
0!
0%
#179935000000
1!
1%
#179940000000
0!
0%
#179945000000
1!
1%
#179950000000
0!
0%
#179955000000
1!
1%
#179960000000
0!
0%
#179965000000
1!
1%
#179970000000
0!
0%
#179975000000
1!
1%
#179980000000
0!
0%
#179985000000
1!
1%
#179990000000
0!
0%
#179995000000
1!
1%
#180000000000
0!
0%
#180005000000
1!
1%
#180010000000
0!
0%
#180015000000
1!
1%
#180020000000
0!
0%
#180025000000
1!
1%
#180030000000
0!
0%
#180035000000
1!
1%
#180040000000
0!
0%
#180045000000
1!
1%
#180050000000
0!
0%
#180055000000
1!
1%
#180060000000
0!
0%
#180065000000
1!
1%
#180070000000
0!
0%
#180075000000
1!
1%
#180080000000
0!
0%
#180085000000
1!
1%
#180090000000
0!
0%
#180095000000
1!
1%
#180100000000
0!
0%
#180105000000
1!
1%
#180110000000
0!
0%
#180115000000
1!
1%
#180120000000
0!
0%
#180125000000
1!
1%
#180130000000
0!
0%
#180135000000
1!
1%
#180140000000
0!
0%
#180145000000
1!
1%
#180150000000
0!
0%
#180155000000
1!
1%
#180160000000
0!
0%
#180165000000
1!
1%
#180170000000
0!
0%
#180175000000
1!
1%
#180180000000
0!
0%
#180185000000
1!
1%
#180190000000
0!
0%
#180195000000
1!
1%
#180200000000
0!
0%
#180205000000
1!
1%
#180210000000
0!
0%
#180215000000
1!
1%
#180220000000
0!
0%
#180225000000
1!
1%
#180230000000
0!
0%
#180235000000
1!
1%
#180240000000
0!
0%
#180245000000
1!
1%
#180250000000
0!
0%
#180255000000
1!
1%
#180260000000
0!
0%
#180265000000
1!
1%
#180270000000
0!
0%
#180275000000
1!
1%
#180280000000
0!
0%
#180285000000
1!
1%
#180290000000
0!
0%
#180295000000
1!
1%
#180300000000
0!
0%
#180305000000
1!
1%
#180310000000
0!
0%
#180315000000
1!
1%
#180320000000
0!
0%
#180325000000
1!
1%
#180330000000
0!
0%
#180335000000
1!
1%
#180340000000
0!
0%
#180345000000
1!
1%
#180350000000
0!
0%
#180355000000
1!
1%
#180360000000
0!
0%
#180365000000
1!
1%
#180370000000
0!
0%
#180375000000
1!
1%
#180380000000
0!
0%
#180385000000
1!
1%
#180390000000
0!
0%
#180395000000
1!
1%
#180400000000
0!
0%
#180405000000
1!
1%
#180410000000
0!
0%
#180415000000
1!
1%
#180420000000
0!
0%
#180425000000
1!
1%
#180430000000
0!
0%
#180435000000
1!
1%
#180440000000
0!
0%
#180445000000
1!
1%
#180450000000
0!
0%
#180455000000
1!
1%
#180460000000
0!
0%
#180465000000
1!
1%
#180470000000
0!
0%
#180475000000
1!
1%
#180480000000
0!
0%
#180485000000
1!
1%
#180490000000
0!
0%
#180495000000
1!
1%
#180500000000
0!
0%
#180505000000
1!
1%
#180510000000
0!
0%
#180515000000
1!
1%
#180520000000
0!
0%
#180525000000
1!
1%
#180530000000
0!
0%
#180535000000
1!
1%
#180540000000
0!
0%
#180545000000
1!
1%
#180550000000
0!
0%
#180555000000
1!
1%
#180560000000
0!
0%
#180565000000
1!
1%
#180570000000
0!
0%
#180575000000
1!
1%
#180580000000
0!
0%
#180585000000
1!
1%
#180590000000
0!
0%
#180595000000
1!
1%
#180600000000
0!
0%
#180605000000
1!
1%
#180610000000
0!
0%
#180615000000
1!
1%
#180620000000
0!
0%
#180625000000
1!
1%
#180630000000
0!
0%
#180635000000
1!
1%
#180640000000
0!
0%
#180645000000
1!
1%
#180650000000
0!
0%
#180655000000
1!
1%
#180660000000
0!
0%
#180665000000
1!
1%
#180670000000
0!
0%
#180675000000
1!
1%
#180680000000
0!
0%
#180685000000
1!
1%
#180690000000
0!
0%
#180695000000
1!
1%
#180700000000
0!
0%
#180705000000
1!
1%
#180710000000
0!
0%
#180715000000
1!
1%
#180720000000
0!
0%
#180725000000
1!
1%
#180730000000
0!
0%
#180735000000
1!
1%
#180740000000
0!
0%
#180745000000
1!
1%
#180750000000
0!
0%
#180755000000
1!
1%
#180760000000
0!
0%
#180765000000
1!
1%
#180770000000
0!
0%
#180775000000
1!
1%
#180780000000
0!
0%
#180785000000
1!
1%
#180790000000
0!
0%
#180795000000
1!
1%
#180800000000
0!
0%
#180805000000
1!
1%
#180810000000
0!
0%
#180815000000
1!
1%
#180820000000
0!
0%
#180825000000
1!
1%
#180830000000
0!
0%
#180835000000
1!
1%
#180840000000
0!
0%
#180845000000
1!
1%
#180850000000
0!
0%
#180855000000
1!
1%
#180860000000
0!
0%
#180865000000
1!
1%
#180870000000
0!
0%
#180875000000
1!
1%
#180880000000
0!
0%
#180885000000
1!
1%
#180890000000
0!
0%
#180895000000
1!
1%
#180900000000
0!
0%
#180905000000
1!
1%
#180910000000
0!
0%
#180915000000
1!
1%
#180920000000
0!
0%
#180925000000
1!
1%
#180930000000
0!
0%
#180935000000
1!
1%
#180940000000
0!
0%
#180945000000
1!
1%
#180950000000
0!
0%
#180955000000
1!
1%
#180960000000
0!
0%
#180965000000
1!
1%
#180970000000
0!
0%
#180975000000
1!
1%
#180980000000
0!
0%
#180985000000
1!
1%
#180990000000
0!
0%
#180995000000
1!
1%
#181000000000
0!
0%
#181005000000
1!
1%
#181010000000
0!
0%
#181015000000
1!
1%
#181020000000
0!
0%
#181025000000
1!
1%
#181030000000
0!
0%
#181035000000
1!
1%
#181040000000
0!
0%
#181045000000
1!
1%
#181050000000
0!
0%
#181055000000
1!
1%
#181060000000
0!
0%
#181065000000
1!
1%
#181070000000
0!
0%
#181075000000
1!
1%
#181080000000
0!
0%
#181085000000
1!
1%
#181090000000
0!
0%
#181095000000
1!
1%
#181100000000
0!
0%
#181105000000
1!
1%
#181110000000
0!
0%
#181115000000
1!
1%
#181120000000
0!
0%
#181125000000
1!
1%
#181130000000
0!
0%
#181135000000
1!
1%
#181140000000
0!
0%
#181145000000
1!
1%
#181150000000
0!
0%
#181155000000
1!
1%
#181160000000
0!
0%
#181165000000
1!
1%
#181170000000
0!
0%
#181175000000
1!
1%
#181180000000
0!
0%
#181185000000
1!
1%
#181190000000
0!
0%
#181195000000
1!
1%
#181200000000
0!
0%
#181205000000
1!
1%
#181210000000
0!
0%
#181215000000
1!
1%
#181220000000
0!
0%
#181225000000
1!
1%
#181230000000
0!
0%
#181235000000
1!
1%
#181240000000
0!
0%
#181245000000
1!
1%
#181250000000
0!
0%
#181255000000
1!
1%
#181260000000
0!
0%
#181265000000
1!
1%
#181270000000
0!
0%
#181275000000
1!
1%
#181280000000
0!
0%
#181285000000
1!
1%
#181290000000
0!
0%
#181295000000
1!
1%
#181300000000
0!
0%
#181305000000
1!
1%
#181310000000
0!
0%
#181315000000
1!
1%
#181320000000
0!
0%
#181325000000
1!
1%
#181330000000
0!
0%
#181335000000
1!
1%
#181340000000
0!
0%
#181345000000
1!
1%
#181350000000
0!
0%
#181355000000
1!
1%
#181360000000
0!
0%
#181365000000
1!
1%
#181370000000
0!
0%
#181375000000
1!
1%
#181380000000
0!
0%
#181385000000
1!
1%
#181390000000
0!
0%
#181395000000
1!
1%
#181400000000
0!
0%
#181405000000
1!
1%
#181410000000
0!
0%
#181415000000
1!
1%
#181420000000
0!
0%
#181425000000
1!
1%
#181430000000
0!
0%
#181435000000
1!
1%
#181440000000
0!
0%
#181445000000
1!
1%
#181450000000
0!
0%
#181455000000
1!
1%
#181460000000
0!
0%
#181465000000
1!
1%
#181470000000
0!
0%
#181475000000
1!
1%
#181480000000
0!
0%
#181485000000
1!
1%
#181490000000
0!
0%
#181495000000
1!
1%
#181500000000
0!
0%
#181505000000
1!
1%
#181510000000
0!
0%
#181515000000
1!
1%
#181520000000
0!
0%
#181525000000
1!
1%
#181530000000
0!
0%
#181535000000
1!
1%
#181540000000
0!
0%
#181545000000
1!
1%
#181550000000
0!
0%
#181555000000
1!
1%
#181560000000
0!
0%
#181565000000
1!
1%
#181570000000
0!
0%
#181575000000
1!
1%
#181580000000
0!
0%
#181585000000
1!
1%
#181590000000
0!
0%
#181595000000
1!
1%
#181600000000
0!
0%
#181605000000
1!
1%
#181610000000
0!
0%
#181615000000
1!
1%
#181620000000
0!
0%
#181625000000
1!
1%
#181630000000
0!
0%
#181635000000
1!
1%
#181640000000
0!
0%
#181645000000
1!
1%
#181650000000
0!
0%
#181655000000
1!
1%
#181660000000
0!
0%
#181665000000
1!
1%
#181670000000
0!
0%
#181675000000
1!
1%
#181680000000
0!
0%
#181685000000
1!
1%
#181690000000
0!
0%
#181695000000
1!
1%
#181700000000
0!
0%
#181705000000
1!
1%
#181710000000
0!
0%
#181715000000
1!
1%
#181720000000
0!
0%
#181725000000
1!
1%
#181730000000
0!
0%
#181735000000
1!
1%
#181740000000
0!
0%
#181745000000
1!
1%
#181750000000
0!
0%
#181755000000
1!
1%
#181760000000
0!
0%
#181765000000
1!
1%
#181770000000
0!
0%
#181775000000
1!
1%
#181780000000
0!
0%
#181785000000
1!
1%
#181790000000
0!
0%
#181795000000
1!
1%
#181800000000
0!
0%
#181805000000
1!
1%
#181810000000
0!
0%
#181815000000
1!
1%
#181820000000
0!
0%
#181825000000
1!
1%
#181830000000
0!
0%
#181835000000
1!
1%
#181840000000
0!
0%
#181845000000
1!
1%
#181850000000
0!
0%
#181855000000
1!
1%
#181860000000
0!
0%
#181865000000
1!
1%
#181870000000
0!
0%
#181875000000
1!
1%
#181880000000
0!
0%
#181885000000
1!
1%
#181890000000
0!
0%
#181895000000
1!
1%
#181900000000
0!
0%
#181905000000
1!
1%
#181910000000
0!
0%
#181915000000
1!
1%
#181920000000
0!
0%
#181925000000
1!
1%
#181930000000
0!
0%
#181935000000
1!
1%
#181940000000
0!
0%
#181945000000
1!
1%
#181950000000
0!
0%
#181955000000
1!
1%
#181960000000
0!
0%
#181965000000
1!
1%
#181970000000
0!
0%
#181975000000
1!
1%
#181980000000
0!
0%
#181985000000
1!
1%
#181990000000
0!
0%
#181995000000
1!
1%
#182000000000
0!
0%
#182005000000
1!
1%
#182010000000
0!
0%
#182015000000
1!
1%
#182020000000
0!
0%
#182025000000
1!
1%
#182030000000
0!
0%
#182035000000
1!
1%
#182040000000
0!
0%
#182045000000
1!
1%
#182050000000
0!
0%
#182055000000
1!
1%
#182060000000
0!
0%
#182065000000
1!
1%
#182070000000
0!
0%
#182075000000
1!
1%
#182080000000
0!
0%
#182085000000
1!
1%
#182090000000
0!
0%
#182095000000
1!
1%
#182100000000
0!
0%
#182105000000
1!
1%
#182110000000
0!
0%
#182115000000
1!
1%
#182120000000
0!
0%
#182125000000
1!
1%
#182130000000
0!
0%
#182135000000
1!
1%
#182140000000
0!
0%
#182145000000
1!
1%
#182150000000
0!
0%
#182155000000
1!
1%
#182160000000
0!
0%
#182165000000
1!
1%
#182170000000
0!
0%
#182175000000
1!
1%
#182180000000
0!
0%
#182185000000
1!
1%
#182190000000
0!
0%
#182195000000
1!
1%
#182200000000
0!
0%
#182205000000
1!
1%
#182210000000
0!
0%
#182215000000
1!
1%
#182220000000
0!
0%
#182225000000
1!
1%
#182230000000
0!
0%
#182235000000
1!
1%
#182240000000
0!
0%
#182245000000
1!
1%
#182250000000
0!
0%
#182255000000
1!
1%
#182260000000
0!
0%
#182265000000
1!
1%
#182270000000
0!
0%
#182275000000
1!
1%
#182280000000
0!
0%
#182285000000
1!
1%
#182290000000
0!
0%
#182295000000
1!
1%
#182300000000
0!
0%
#182305000000
1!
1%
#182310000000
0!
0%
#182315000000
1!
1%
#182320000000
0!
0%
#182325000000
1!
1%
#182330000000
0!
0%
#182335000000
1!
1%
#182340000000
0!
0%
#182345000000
1!
1%
#182350000000
0!
0%
#182355000000
1!
1%
#182360000000
0!
0%
#182365000000
1!
1%
#182370000000
0!
0%
#182375000000
1!
1%
#182380000000
0!
0%
#182385000000
1!
1%
#182390000000
0!
0%
#182395000000
1!
1%
#182400000000
0!
0%
#182405000000
1!
1%
#182410000000
0!
0%
#182415000000
1!
1%
#182420000000
0!
0%
#182425000000
1!
1%
#182430000000
0!
0%
#182435000000
1!
1%
#182440000000
0!
0%
#182445000000
1!
1%
#182450000000
0!
0%
#182455000000
1!
1%
#182460000000
0!
0%
#182465000000
1!
1%
#182470000000
0!
0%
#182475000000
1!
1%
#182480000000
0!
0%
#182485000000
1!
1%
#182490000000
0!
0%
#182495000000
1!
1%
#182500000000
0!
0%
#182505000000
1!
1%
#182510000000
0!
0%
#182515000000
1!
1%
#182520000000
0!
0%
#182525000000
1!
1%
#182530000000
0!
0%
#182535000000
1!
1%
#182540000000
0!
0%
#182545000000
1!
1%
#182550000000
0!
0%
#182555000000
1!
1%
#182560000000
0!
0%
#182565000000
1!
1%
#182570000000
0!
0%
#182575000000
1!
1%
#182580000000
0!
0%
#182585000000
1!
1%
#182590000000
0!
0%
#182595000000
1!
1%
#182600000000
0!
0%
#182605000000
1!
1%
#182610000000
0!
0%
#182615000000
1!
1%
#182620000000
0!
0%
#182625000000
1!
1%
#182630000000
0!
0%
#182635000000
1!
1%
#182640000000
0!
0%
#182645000000
1!
1%
#182650000000
0!
0%
#182655000000
1!
1%
#182660000000
0!
0%
#182665000000
1!
1%
#182670000000
0!
0%
#182675000000
1!
1%
#182680000000
0!
0%
#182685000000
1!
1%
#182690000000
0!
0%
#182695000000
1!
1%
#182700000000
0!
0%
#182705000000
1!
1%
#182710000000
0!
0%
#182715000000
1!
1%
#182720000000
0!
0%
#182725000000
1!
1%
#182730000000
0!
0%
#182735000000
1!
1%
#182740000000
0!
0%
#182745000000
1!
1%
#182750000000
0!
0%
#182755000000
1!
1%
#182760000000
0!
0%
#182765000000
1!
1%
#182770000000
0!
0%
#182775000000
1!
1%
#182780000000
0!
0%
#182785000000
1!
1%
#182790000000
0!
0%
#182795000000
1!
1%
#182800000000
0!
0%
#182805000000
1!
1%
#182810000000
0!
0%
#182815000000
1!
1%
#182820000000
0!
0%
#182825000000
1!
1%
#182830000000
0!
0%
#182835000000
1!
1%
#182840000000
0!
0%
#182845000000
1!
1%
#182850000000
0!
0%
#182855000000
1!
1%
#182860000000
0!
0%
#182865000000
1!
1%
#182870000000
0!
0%
#182875000000
1!
1%
#182880000000
0!
0%
#182885000000
1!
1%
#182890000000
0!
0%
#182895000000
1!
1%
#182900000000
0!
0%
#182905000000
1!
1%
#182910000000
0!
0%
#182915000000
1!
1%
#182920000000
0!
0%
#182925000000
1!
1%
#182930000000
0!
0%
#182935000000
1!
1%
#182940000000
0!
0%
#182945000000
1!
1%
#182950000000
0!
0%
#182955000000
1!
1%
#182960000000
0!
0%
#182965000000
1!
1%
#182970000000
0!
0%
#182975000000
1!
1%
#182980000000
0!
0%
#182985000000
1!
1%
#182990000000
0!
0%
#182995000000
1!
1%
#183000000000
0!
0%
#183005000000
1!
1%
#183010000000
0!
0%
#183015000000
1!
1%
#183020000000
0!
0%
#183025000000
1!
1%
#183030000000
0!
0%
#183035000000
1!
1%
#183040000000
0!
0%
#183045000000
1!
1%
#183050000000
0!
0%
#183055000000
1!
1%
#183060000000
0!
0%
#183065000000
1!
1%
#183070000000
0!
0%
#183075000000
1!
1%
#183080000000
0!
0%
#183085000000
1!
1%
#183090000000
0!
0%
#183095000000
1!
1%
#183100000000
0!
0%
#183105000000
1!
1%
#183110000000
0!
0%
#183115000000
1!
1%
#183120000000
0!
0%
#183125000000
1!
1%
#183130000000
0!
0%
#183135000000
1!
1%
#183140000000
0!
0%
#183145000000
1!
1%
#183150000000
0!
0%
#183155000000
1!
1%
#183160000000
0!
0%
#183165000000
1!
1%
#183170000000
0!
0%
#183175000000
1!
1%
#183180000000
0!
0%
#183185000000
1!
1%
#183190000000
0!
0%
#183195000000
1!
1%
#183200000000
0!
0%
#183205000000
1!
1%
#183210000000
0!
0%
#183215000000
1!
1%
#183220000000
0!
0%
#183225000000
1!
1%
#183230000000
0!
0%
#183235000000
1!
1%
#183240000000
0!
0%
#183245000000
1!
1%
#183250000000
0!
0%
#183255000000
1!
1%
#183260000000
0!
0%
#183265000000
1!
1%
#183270000000
0!
0%
#183275000000
1!
1%
#183280000000
0!
0%
#183285000000
1!
1%
#183290000000
0!
0%
#183295000000
1!
1%
#183300000000
0!
0%
#183305000000
1!
1%
#183310000000
0!
0%
#183315000000
1!
1%
#183320000000
0!
0%
#183325000000
1!
1%
#183330000000
0!
0%
#183335000000
1!
1%
#183340000000
0!
0%
#183345000000
1!
1%
#183350000000
0!
0%
#183355000000
1!
1%
#183360000000
0!
0%
#183365000000
1!
1%
#183370000000
0!
0%
#183375000000
1!
1%
#183380000000
0!
0%
#183385000000
1!
1%
#183390000000
0!
0%
#183395000000
1!
1%
#183400000000
0!
0%
#183405000000
1!
1%
#183410000000
0!
0%
#183415000000
1!
1%
#183420000000
0!
0%
#183425000000
1!
1%
#183430000000
0!
0%
#183435000000
1!
1%
#183440000000
0!
0%
#183445000000
1!
1%
#183450000000
0!
0%
#183455000000
1!
1%
#183460000000
0!
0%
#183465000000
1!
1%
#183470000000
0!
0%
#183475000000
1!
1%
#183480000000
0!
0%
#183485000000
1!
1%
#183490000000
0!
0%
#183495000000
1!
1%
#183500000000
0!
0%
#183505000000
1!
1%
#183510000000
0!
0%
#183515000000
1!
1%
#183520000000
0!
0%
#183525000000
1!
1%
#183530000000
0!
0%
#183535000000
1!
1%
#183540000000
0!
0%
#183545000000
1!
1%
#183550000000
0!
0%
#183555000000
1!
1%
#183560000000
0!
0%
#183565000000
1!
1%
#183570000000
0!
0%
#183575000000
1!
1%
#183580000000
0!
0%
#183585000000
1!
1%
#183590000000
0!
0%
#183595000000
1!
1%
#183600000000
0!
0%
#183605000000
1!
1%
#183610000000
0!
0%
#183615000000
1!
1%
#183620000000
0!
0%
#183625000000
1!
1%
#183630000000
0!
0%
#183635000000
1!
1%
#183640000000
0!
0%
#183645000000
1!
1%
#183650000000
0!
0%
#183655000000
1!
1%
#183660000000
0!
0%
#183665000000
1!
1%
#183670000000
0!
0%
#183675000000
1!
1%
#183680000000
0!
0%
#183685000000
1!
1%
#183690000000
0!
0%
#183695000000
1!
1%
#183700000000
0!
0%
#183705000000
1!
1%
#183710000000
0!
0%
#183715000000
1!
1%
#183720000000
0!
0%
#183725000000
1!
1%
#183730000000
0!
0%
#183735000000
1!
1%
#183740000000
0!
0%
#183745000000
1!
1%
#183750000000
0!
0%
#183755000000
1!
1%
#183760000000
0!
0%
#183765000000
1!
1%
#183770000000
0!
0%
#183775000000
1!
1%
#183780000000
0!
0%
#183785000000
1!
1%
#183790000000
0!
0%
#183795000000
1!
1%
#183800000000
0!
0%
#183805000000
1!
1%
#183810000000
0!
0%
#183815000000
1!
1%
#183820000000
0!
0%
#183825000000
1!
1%
#183830000000
0!
0%
#183835000000
1!
1%
#183840000000
0!
0%
#183845000000
1!
1%
#183850000000
0!
0%
#183855000000
1!
1%
#183860000000
0!
0%
#183865000000
1!
1%
#183870000000
0!
0%
#183875000000
1!
1%
#183880000000
0!
0%
#183885000000
1!
1%
#183890000000
0!
0%
#183895000000
1!
1%
#183900000000
0!
0%
#183905000000
1!
1%
#183910000000
0!
0%
#183915000000
1!
1%
#183920000000
0!
0%
#183925000000
1!
1%
#183930000000
0!
0%
#183935000000
1!
1%
#183940000000
0!
0%
#183945000000
1!
1%
#183950000000
0!
0%
#183955000000
1!
1%
#183960000000
0!
0%
#183965000000
1!
1%
#183970000000
0!
0%
#183975000000
1!
1%
#183980000000
0!
0%
#183985000000
1!
1%
#183990000000
0!
0%
#183995000000
1!
1%
#184000000000
0!
0%
#184005000000
1!
1%
#184010000000
0!
0%
#184015000000
1!
1%
#184020000000
0!
0%
#184025000000
1!
1%
#184030000000
0!
0%
#184035000000
1!
1%
#184040000000
0!
0%
#184045000000
1!
1%
#184050000000
0!
0%
#184055000000
1!
1%
#184060000000
0!
0%
#184065000000
1!
1%
#184070000000
0!
0%
#184075000000
1!
1%
#184080000000
0!
0%
#184085000000
1!
1%
#184090000000
0!
0%
#184095000000
1!
1%
#184100000000
0!
0%
#184105000000
1!
1%
#184110000000
0!
0%
#184115000000
1!
1%
#184120000000
0!
0%
#184125000000
1!
1%
#184130000000
0!
0%
#184135000000
1!
1%
#184140000000
0!
0%
#184145000000
1!
1%
#184150000000
0!
0%
#184155000000
1!
1%
#184160000000
0!
0%
#184165000000
1!
1%
#184170000000
0!
0%
#184175000000
1!
1%
#184180000000
0!
0%
#184185000000
1!
1%
#184190000000
0!
0%
#184195000000
1!
1%
#184200000000
0!
0%
#184205000000
1!
1%
#184210000000
0!
0%
#184215000000
1!
1%
#184220000000
0!
0%
#184225000000
1!
1%
#184230000000
0!
0%
#184235000000
1!
1%
#184240000000
0!
0%
#184245000000
1!
1%
#184250000000
0!
0%
#184255000000
1!
1%
#184260000000
0!
0%
#184265000000
1!
1%
#184270000000
0!
0%
#184275000000
1!
1%
#184280000000
0!
0%
#184285000000
1!
1%
#184290000000
0!
0%
#184295000000
1!
1%
#184300000000
0!
0%
#184305000000
1!
1%
#184310000000
0!
0%
#184315000000
1!
1%
#184320000000
0!
0%
#184325000000
1!
1%
#184330000000
0!
0%
#184335000000
1!
1%
#184340000000
0!
0%
#184345000000
1!
1%
#184350000000
0!
0%
#184355000000
1!
1%
#184360000000
0!
0%
#184365000000
1!
1%
#184370000000
0!
0%
#184375000000
1!
1%
#184380000000
0!
0%
#184385000000
1!
1%
#184390000000
0!
0%
#184395000000
1!
1%
#184400000000
0!
0%
#184405000000
1!
1%
#184410000000
0!
0%
#184415000000
1!
1%
#184420000000
0!
0%
#184425000000
1!
1%
#184430000000
0!
0%
#184435000000
1!
1%
#184440000000
0!
0%
#184445000000
1!
1%
#184450000000
0!
0%
#184455000000
1!
1%
#184460000000
0!
0%
#184465000000
1!
1%
#184470000000
0!
0%
#184475000000
1!
1%
#184480000000
0!
0%
#184485000000
1!
1%
#184490000000
0!
0%
#184495000000
1!
1%
#184500000000
0!
0%
#184505000000
1!
1%
#184510000000
0!
0%
#184515000000
1!
1%
#184520000000
0!
0%
#184525000000
1!
1%
#184530000000
0!
0%
#184535000000
1!
1%
#184540000000
0!
0%
#184545000000
1!
1%
#184550000000
0!
0%
#184555000000
1!
1%
#184560000000
0!
0%
#184565000000
1!
1%
#184570000000
0!
0%
#184575000000
1!
1%
#184580000000
0!
0%
#184585000000
1!
1%
#184590000000
0!
0%
#184595000000
1!
1%
#184600000000
0!
0%
#184605000000
1!
1%
#184610000000
0!
0%
#184615000000
1!
1%
#184620000000
0!
0%
#184625000000
1!
1%
#184630000000
0!
0%
#184635000000
1!
1%
#184640000000
0!
0%
#184645000000
1!
1%
#184650000000
0!
0%
#184655000000
1!
1%
#184660000000
0!
0%
#184665000000
1!
1%
#184670000000
0!
0%
#184675000000
1!
1%
#184680000000
0!
0%
#184685000000
1!
1%
#184690000000
0!
0%
#184695000000
1!
1%
#184700000000
0!
0%
#184705000000
1!
1%
#184710000000
0!
0%
#184715000000
1!
1%
#184720000000
0!
0%
#184725000000
1!
1%
#184730000000
0!
0%
#184735000000
1!
1%
#184740000000
0!
0%
#184745000000
1!
1%
#184750000000
0!
0%
#184755000000
1!
1%
#184760000000
0!
0%
#184765000000
1!
1%
#184770000000
0!
0%
#184775000000
1!
1%
#184780000000
0!
0%
#184785000000
1!
1%
#184790000000
0!
0%
#184795000000
1!
1%
#184800000000
0!
0%
#184805000000
1!
1%
#184810000000
0!
0%
#184815000000
1!
1%
#184820000000
0!
0%
#184825000000
1!
1%
#184830000000
0!
0%
#184835000000
1!
1%
#184840000000
0!
0%
#184845000000
1!
1%
#184850000000
0!
0%
#184855000000
1!
1%
#184860000000
0!
0%
#184865000000
1!
1%
#184870000000
0!
0%
#184875000000
1!
1%
#184880000000
0!
0%
#184885000000
1!
1%
#184890000000
0!
0%
#184895000000
1!
1%
#184900000000
0!
0%
#184905000000
1!
1%
#184910000000
0!
0%
#184915000000
1!
1%
#184920000000
0!
0%
#184925000000
1!
1%
#184930000000
0!
0%
#184935000000
1!
1%
#184940000000
0!
0%
#184945000000
1!
1%
#184950000000
0!
0%
#184955000000
1!
1%
#184960000000
0!
0%
#184965000000
1!
1%
#184970000000
0!
0%
#184975000000
1!
1%
#184980000000
0!
0%
#184985000000
1!
1%
#184990000000
0!
0%
#184995000000
1!
1%
#185000000000
0!
0%
#185005000000
1!
1%
#185010000000
0!
0%
#185015000000
1!
1%
#185020000000
0!
0%
#185025000000
1!
1%
#185030000000
0!
0%
#185035000000
1!
1%
#185040000000
0!
0%
#185045000000
1!
1%
#185050000000
0!
0%
#185055000000
1!
1%
#185060000000
0!
0%
#185065000000
1!
1%
#185070000000
0!
0%
#185075000000
1!
1%
#185080000000
0!
0%
#185085000000
1!
1%
#185090000000
0!
0%
#185095000000
1!
1%
#185100000000
0!
0%
#185105000000
1!
1%
#185110000000
0!
0%
#185115000000
1!
1%
#185120000000
0!
0%
#185125000000
1!
1%
#185130000000
0!
0%
#185135000000
1!
1%
#185140000000
0!
0%
#185145000000
1!
1%
#185150000000
0!
0%
#185155000000
1!
1%
#185160000000
0!
0%
#185165000000
1!
1%
#185170000000
0!
0%
#185175000000
1!
1%
#185180000000
0!
0%
#185185000000
1!
1%
#185190000000
0!
0%
#185195000000
1!
1%
#185200000000
0!
0%
#185205000000
1!
1%
#185210000000
0!
0%
#185215000000
1!
1%
#185220000000
0!
0%
#185225000000
1!
1%
#185230000000
0!
0%
#185235000000
1!
1%
#185240000000
0!
0%
#185245000000
1!
1%
#185250000000
0!
0%
#185255000000
1!
1%
#185260000000
0!
0%
#185265000000
1!
1%
#185270000000
0!
0%
#185275000000
1!
1%
#185280000000
0!
0%
#185285000000
1!
1%
#185290000000
0!
0%
#185295000000
1!
1%
#185300000000
0!
0%
#185305000000
1!
1%
#185310000000
0!
0%
#185315000000
1!
1%
#185320000000
0!
0%
#185325000000
1!
1%
#185330000000
0!
0%
#185335000000
1!
1%
#185340000000
0!
0%
#185345000000
1!
1%
#185350000000
0!
0%
#185355000000
1!
1%
#185360000000
0!
0%
#185365000000
1!
1%
#185370000000
0!
0%
#185375000000
1!
1%
#185380000000
0!
0%
#185385000000
1!
1%
#185390000000
0!
0%
#185395000000
1!
1%
#185400000000
0!
0%
#185405000000
1!
1%
#185410000000
0!
0%
#185415000000
1!
1%
#185420000000
0!
0%
#185425000000
1!
1%
#185430000000
0!
0%
#185435000000
1!
1%
#185440000000
0!
0%
#185445000000
1!
1%
#185450000000
0!
0%
#185455000000
1!
1%
#185460000000
0!
0%
#185465000000
1!
1%
#185470000000
0!
0%
#185475000000
1!
1%
#185480000000
0!
0%
#185485000000
1!
1%
#185490000000
0!
0%
#185495000000
1!
1%
#185500000000
0!
0%
#185505000000
1!
1%
#185510000000
0!
0%
#185515000000
1!
1%
#185520000000
0!
0%
#185525000000
1!
1%
#185530000000
0!
0%
#185535000000
1!
1%
#185540000000
0!
0%
#185545000000
1!
1%
#185550000000
0!
0%
#185555000000
1!
1%
#185560000000
0!
0%
#185565000000
1!
1%
#185570000000
0!
0%
#185575000000
1!
1%
#185580000000
0!
0%
#185585000000
1!
1%
#185590000000
0!
0%
#185595000000
1!
1%
#185600000000
0!
0%
#185605000000
1!
1%
#185610000000
0!
0%
#185615000000
1!
1%
#185620000000
0!
0%
#185625000000
1!
1%
#185630000000
0!
0%
#185635000000
1!
1%
#185640000000
0!
0%
#185645000000
1!
1%
#185650000000
0!
0%
#185655000000
1!
1%
#185660000000
0!
0%
#185665000000
1!
1%
#185670000000
0!
0%
#185675000000
1!
1%
#185680000000
0!
0%
#185685000000
1!
1%
#185690000000
0!
0%
#185695000000
1!
1%
#185700000000
0!
0%
#185705000000
1!
1%
#185710000000
0!
0%
#185715000000
1!
1%
#185720000000
0!
0%
#185725000000
1!
1%
#185730000000
0!
0%
#185735000000
1!
1%
#185740000000
0!
0%
#185745000000
1!
1%
#185750000000
0!
0%
#185755000000
1!
1%
#185760000000
0!
0%
#185765000000
1!
1%
#185770000000
0!
0%
#185775000000
1!
1%
#185780000000
0!
0%
#185785000000
1!
1%
#185790000000
0!
0%
#185795000000
1!
1%
#185800000000
0!
0%
#185805000000
1!
1%
#185810000000
0!
0%
#185815000000
1!
1%
#185820000000
0!
0%
#185825000000
1!
1%
#185830000000
0!
0%
#185835000000
1!
1%
#185840000000
0!
0%
#185845000000
1!
1%
#185850000000
0!
0%
#185855000000
1!
1%
#185860000000
0!
0%
#185865000000
1!
1%
#185870000000
0!
0%
#185875000000
1!
1%
#185880000000
0!
0%
#185885000000
1!
1%
#185890000000
0!
0%
#185895000000
1!
1%
#185900000000
0!
0%
#185905000000
1!
1%
#185910000000
0!
0%
#185915000000
1!
1%
#185920000000
0!
0%
#185925000000
1!
1%
#185930000000
0!
0%
#185935000000
1!
1%
#185940000000
0!
0%
#185945000000
1!
1%
#185950000000
0!
0%
#185955000000
1!
1%
#185960000000
0!
0%
#185965000000
1!
1%
#185970000000
0!
0%
#185975000000
1!
1%
#185980000000
0!
0%
#185985000000
1!
1%
#185990000000
0!
0%
#185995000000
1!
1%
#186000000000
0!
0%
#186005000000
1!
1%
#186010000000
0!
0%
#186015000000
1!
1%
#186020000000
0!
0%
#186025000000
1!
1%
#186030000000
0!
0%
#186035000000
1!
1%
#186040000000
0!
0%
#186045000000
1!
1%
#186050000000
0!
0%
#186055000000
1!
1%
#186060000000
0!
0%
#186065000000
1!
1%
#186070000000
0!
0%
#186075000000
1!
1%
#186080000000
0!
0%
#186085000000
1!
1%
#186090000000
0!
0%
#186095000000
1!
1%
#186100000000
0!
0%
#186105000000
1!
1%
#186110000000
0!
0%
#186115000000
1!
1%
#186120000000
0!
0%
#186125000000
1!
1%
#186130000000
0!
0%
#186135000000
1!
1%
#186140000000
0!
0%
#186145000000
1!
1%
#186150000000
0!
0%
#186155000000
1!
1%
#186160000000
0!
0%
#186165000000
1!
1%
#186170000000
0!
0%
#186175000000
1!
1%
#186180000000
0!
0%
#186185000000
1!
1%
#186190000000
0!
0%
#186195000000
1!
1%
#186200000000
0!
0%
#186205000000
1!
1%
#186210000000
0!
0%
#186215000000
1!
1%
#186220000000
0!
0%
#186225000000
1!
1%
#186230000000
0!
0%
#186235000000
1!
1%
#186240000000
0!
0%
#186245000000
1!
1%
#186250000000
0!
0%
#186255000000
1!
1%
#186260000000
0!
0%
#186265000000
1!
1%
#186270000000
0!
0%
#186275000000
1!
1%
#186280000000
0!
0%
#186285000000
1!
1%
#186290000000
0!
0%
#186295000000
1!
1%
#186300000000
0!
0%
#186305000000
1!
1%
#186310000000
0!
0%
#186315000000
1!
1%
#186320000000
0!
0%
#186325000000
1!
1%
#186330000000
0!
0%
#186335000000
1!
1%
#186340000000
0!
0%
#186345000000
1!
1%
#186350000000
0!
0%
#186355000000
1!
1%
#186360000000
0!
0%
#186365000000
1!
1%
#186370000000
0!
0%
#186375000000
1!
1%
#186380000000
0!
0%
#186385000000
1!
1%
#186390000000
0!
0%
#186395000000
1!
1%
#186400000000
0!
0%
#186405000000
1!
1%
#186410000000
0!
0%
#186415000000
1!
1%
#186420000000
0!
0%
#186425000000
1!
1%
#186430000000
0!
0%
#186435000000
1!
1%
#186440000000
0!
0%
#186445000000
1!
1%
#186450000000
0!
0%
#186455000000
1!
1%
#186460000000
0!
0%
#186465000000
1!
1%
#186470000000
0!
0%
#186475000000
1!
1%
#186480000000
0!
0%
#186485000000
1!
1%
#186490000000
0!
0%
#186495000000
1!
1%
#186500000000
0!
0%
#186505000000
1!
1%
#186510000000
0!
0%
#186515000000
1!
1%
#186520000000
0!
0%
#186525000000
1!
1%
#186530000000
0!
0%
#186535000000
1!
1%
#186540000000
0!
0%
#186545000000
1!
1%
#186550000000
0!
0%
#186555000000
1!
1%
#186560000000
0!
0%
#186565000000
1!
1%
#186570000000
0!
0%
#186575000000
1!
1%
#186580000000
0!
0%
#186585000000
1!
1%
#186590000000
0!
0%
#186595000000
1!
1%
#186600000000
0!
0%
#186605000000
1!
1%
#186610000000
0!
0%
#186615000000
1!
1%
#186620000000
0!
0%
#186625000000
1!
1%
#186630000000
0!
0%
#186635000000
1!
1%
#186640000000
0!
0%
#186645000000
1!
1%
#186650000000
0!
0%
#186655000000
1!
1%
#186660000000
0!
0%
#186665000000
1!
1%
#186670000000
0!
0%
#186675000000
1!
1%
#186680000000
0!
0%
#186685000000
1!
1%
#186690000000
0!
0%
#186695000000
1!
1%
#186700000000
0!
0%
#186705000000
1!
1%
#186710000000
0!
0%
#186715000000
1!
1%
#186720000000
0!
0%
#186725000000
1!
1%
#186730000000
0!
0%
#186735000000
1!
1%
#186740000000
0!
0%
#186745000000
1!
1%
#186750000000
0!
0%
#186755000000
1!
1%
#186760000000
0!
0%
#186765000000
1!
1%
#186770000000
0!
0%
#186775000000
1!
1%
#186780000000
0!
0%
#186785000000
1!
1%
#186790000000
0!
0%
#186795000000
1!
1%
#186800000000
0!
0%
#186805000000
1!
1%
#186810000000
0!
0%
#186815000000
1!
1%
#186820000000
0!
0%
#186825000000
1!
1%
#186830000000
0!
0%
#186835000000
1!
1%
#186840000000
0!
0%
#186845000000
1!
1%
#186850000000
0!
0%
#186855000000
1!
1%
#186860000000
0!
0%
#186865000000
1!
1%
#186870000000
0!
0%
#186875000000
1!
1%
#186880000000
0!
0%
#186885000000
1!
1%
#186890000000
0!
0%
#186895000000
1!
1%
#186900000000
0!
0%
#186905000000
1!
1%
#186910000000
0!
0%
#186915000000
1!
1%
#186920000000
0!
0%
#186925000000
1!
1%
#186930000000
0!
0%
#186935000000
1!
1%
#186940000000
0!
0%
#186945000000
1!
1%
#186950000000
0!
0%
#186955000000
1!
1%
#186960000000
0!
0%
#186965000000
1!
1%
#186970000000
0!
0%
#186975000000
1!
1%
#186980000000
0!
0%
#186985000000
1!
1%
#186990000000
0!
0%
#186995000000
1!
1%
#187000000000
0!
0%
#187005000000
1!
1%
#187010000000
0!
0%
#187015000000
1!
1%
#187020000000
0!
0%
#187025000000
1!
1%
#187030000000
0!
0%
#187035000000
1!
1%
#187040000000
0!
0%
#187045000000
1!
1%
#187050000000
0!
0%
#187055000000
1!
1%
#187060000000
0!
0%
#187065000000
1!
1%
#187070000000
0!
0%
#187075000000
1!
1%
#187080000000
0!
0%
#187085000000
1!
1%
#187090000000
0!
0%
#187095000000
1!
1%
#187100000000
0!
0%
#187105000000
1!
1%
#187110000000
0!
0%
#187115000000
1!
1%
#187120000000
0!
0%
#187125000000
1!
1%
#187130000000
0!
0%
#187135000000
1!
1%
#187140000000
0!
0%
#187145000000
1!
1%
#187150000000
0!
0%
#187155000000
1!
1%
#187160000000
0!
0%
#187165000000
1!
1%
#187170000000
0!
0%
#187175000000
1!
1%
#187180000000
0!
0%
#187185000000
1!
1%
#187190000000
0!
0%
#187195000000
1!
1%
#187200000000
0!
0%
#187205000000
1!
1%
#187210000000
0!
0%
#187215000000
1!
1%
#187220000000
0!
0%
#187225000000
1!
1%
#187230000000
0!
0%
#187235000000
1!
1%
#187240000000
0!
0%
#187245000000
1!
1%
#187250000000
0!
0%
#187255000000
1!
1%
#187260000000
0!
0%
#187265000000
1!
1%
#187270000000
0!
0%
#187275000000
1!
1%
#187280000000
0!
0%
#187285000000
1!
1%
#187290000000
0!
0%
#187295000000
1!
1%
#187300000000
0!
0%
#187305000000
1!
1%
#187310000000
0!
0%
#187315000000
1!
1%
#187320000000
0!
0%
#187325000000
1!
1%
#187330000000
0!
0%
#187335000000
1!
1%
#187340000000
0!
0%
#187345000000
1!
1%
#187350000000
0!
0%
#187355000000
1!
1%
#187360000000
0!
0%
#187365000000
1!
1%
#187370000000
0!
0%
#187375000000
1!
1%
#187380000000
0!
0%
#187385000000
1!
1%
#187390000000
0!
0%
#187395000000
1!
1%
#187400000000
0!
0%
#187405000000
1!
1%
#187410000000
0!
0%
#187415000000
1!
1%
#187420000000
0!
0%
#187425000000
1!
1%
#187430000000
0!
0%
#187435000000
1!
1%
#187440000000
0!
0%
#187445000000
1!
1%
#187450000000
0!
0%
#187455000000
1!
1%
#187460000000
0!
0%
#187465000000
1!
1%
#187470000000
0!
0%
#187475000000
1!
1%
#187480000000
0!
0%
#187485000000
1!
1%
#187490000000
0!
0%
#187495000000
1!
1%
#187500000000
0!
0%
#187505000000
1!
1%
#187510000000
0!
0%
#187515000000
1!
1%
#187520000000
0!
0%
#187525000000
1!
1%
#187530000000
0!
0%
#187535000000
1!
1%
#187540000000
0!
0%
#187545000000
1!
1%
#187550000000
0!
0%
#187555000000
1!
1%
#187560000000
0!
0%
#187565000000
1!
1%
#187570000000
0!
0%
#187575000000
1!
1%
#187580000000
0!
0%
#187585000000
1!
1%
#187590000000
0!
0%
#187595000000
1!
1%
#187600000000
0!
0%
#187605000000
1!
1%
#187610000000
0!
0%
#187615000000
1!
1%
#187620000000
0!
0%
#187625000000
1!
1%
#187630000000
0!
0%
#187635000000
1!
1%
#187640000000
0!
0%
#187645000000
1!
1%
#187650000000
0!
0%
#187655000000
1!
1%
#187660000000
0!
0%
#187665000000
1!
1%
#187670000000
0!
0%
#187675000000
1!
1%
#187680000000
0!
0%
#187685000000
1!
1%
#187690000000
0!
0%
#187695000000
1!
1%
#187700000000
0!
0%
#187705000000
1!
1%
#187710000000
0!
0%
#187715000000
1!
1%
#187720000000
0!
0%
#187725000000
1!
1%
#187730000000
0!
0%
#187735000000
1!
1%
#187740000000
0!
0%
#187745000000
1!
1%
#187750000000
0!
0%
#187755000000
1!
1%
#187760000000
0!
0%
#187765000000
1!
1%
#187770000000
0!
0%
#187775000000
1!
1%
#187780000000
0!
0%
#187785000000
1!
1%
#187790000000
0!
0%
#187795000000
1!
1%
#187800000000
0!
0%
#187805000000
1!
1%
#187810000000
0!
0%
#187815000000
1!
1%
#187820000000
0!
0%
#187825000000
1!
1%
#187830000000
0!
0%
#187835000000
1!
1%
#187840000000
0!
0%
#187845000000
1!
1%
#187850000000
0!
0%
#187855000000
1!
1%
#187860000000
0!
0%
#187865000000
1!
1%
#187870000000
0!
0%
#187875000000
1!
1%
#187880000000
0!
0%
#187885000000
1!
1%
#187890000000
0!
0%
#187895000000
1!
1%
#187900000000
0!
0%
#187905000000
1!
1%
#187910000000
0!
0%
#187915000000
1!
1%
#187920000000
0!
0%
#187925000000
1!
1%
#187930000000
0!
0%
#187935000000
1!
1%
#187940000000
0!
0%
#187945000000
1!
1%
#187950000000
0!
0%
#187955000000
1!
1%
#187960000000
0!
0%
#187965000000
1!
1%
#187970000000
0!
0%
#187975000000
1!
1%
#187980000000
0!
0%
#187985000000
1!
1%
#187990000000
0!
0%
#187995000000
1!
1%
#188000000000
0!
0%
#188005000000
1!
1%
#188010000000
0!
0%
#188015000000
1!
1%
#188020000000
0!
0%
#188025000000
1!
1%
#188030000000
0!
0%
#188035000000
1!
1%
#188040000000
0!
0%
#188045000000
1!
1%
#188050000000
0!
0%
#188055000000
1!
1%
#188060000000
0!
0%
#188065000000
1!
1%
#188070000000
0!
0%
#188075000000
1!
1%
#188080000000
0!
0%
#188085000000
1!
1%
#188090000000
0!
0%
#188095000000
1!
1%
#188100000000
0!
0%
#188105000000
1!
1%
#188110000000
0!
0%
#188115000000
1!
1%
#188120000000
0!
0%
#188125000000
1!
1%
#188130000000
0!
0%
#188135000000
1!
1%
#188140000000
0!
0%
#188145000000
1!
1%
#188150000000
0!
0%
#188155000000
1!
1%
#188160000000
0!
0%
#188165000000
1!
1%
#188170000000
0!
0%
#188175000000
1!
1%
#188180000000
0!
0%
#188185000000
1!
1%
#188190000000
0!
0%
#188195000000
1!
1%
#188200000000
0!
0%
#188205000000
1!
1%
#188210000000
0!
0%
#188215000000
1!
1%
#188220000000
0!
0%
#188225000000
1!
1%
#188230000000
0!
0%
#188235000000
1!
1%
#188240000000
0!
0%
#188245000000
1!
1%
#188250000000
0!
0%
#188255000000
1!
1%
#188260000000
0!
0%
#188265000000
1!
1%
#188270000000
0!
0%
#188275000000
1!
1%
#188280000000
0!
0%
#188285000000
1!
1%
#188290000000
0!
0%
#188295000000
1!
1%
#188300000000
0!
0%
#188305000000
1!
1%
#188310000000
0!
0%
#188315000000
1!
1%
#188320000000
0!
0%
#188325000000
1!
1%
#188330000000
0!
0%
#188335000000
1!
1%
#188340000000
0!
0%
#188345000000
1!
1%
#188350000000
0!
0%
#188355000000
1!
1%
#188360000000
0!
0%
#188365000000
1!
1%
#188370000000
0!
0%
#188375000000
1!
1%
#188380000000
0!
0%
#188385000000
1!
1%
#188390000000
0!
0%
#188395000000
1!
1%
#188400000000
0!
0%
#188405000000
1!
1%
#188410000000
0!
0%
#188415000000
1!
1%
#188420000000
0!
0%
#188425000000
1!
1%
#188430000000
0!
0%
#188435000000
1!
1%
#188440000000
0!
0%
#188445000000
1!
1%
#188450000000
0!
0%
#188455000000
1!
1%
#188460000000
0!
0%
#188465000000
1!
1%
#188470000000
0!
0%
#188475000000
1!
1%
#188480000000
0!
0%
#188485000000
1!
1%
#188490000000
0!
0%
#188495000000
1!
1%
#188500000000
0!
0%
#188505000000
1!
1%
#188510000000
0!
0%
#188515000000
1!
1%
#188520000000
0!
0%
#188525000000
1!
1%
#188530000000
0!
0%
#188535000000
1!
1%
#188540000000
0!
0%
#188545000000
1!
1%
#188550000000
0!
0%
#188555000000
1!
1%
#188560000000
0!
0%
#188565000000
1!
1%
#188570000000
0!
0%
#188575000000
1!
1%
#188580000000
0!
0%
#188585000000
1!
1%
#188590000000
0!
0%
#188595000000
1!
1%
#188600000000
0!
0%
#188605000000
1!
1%
#188610000000
0!
0%
#188615000000
1!
1%
#188620000000
0!
0%
#188625000000
1!
1%
#188630000000
0!
0%
#188635000000
1!
1%
#188640000000
0!
0%
#188645000000
1!
1%
#188650000000
0!
0%
#188655000000
1!
1%
#188660000000
0!
0%
#188665000000
1!
1%
#188670000000
0!
0%
#188675000000
1!
1%
#188680000000
0!
0%
#188685000000
1!
1%
#188690000000
0!
0%
#188695000000
1!
1%
#188700000000
0!
0%
#188705000000
1!
1%
#188710000000
0!
0%
#188715000000
1!
1%
#188720000000
0!
0%
#188725000000
1!
1%
#188730000000
0!
0%
#188735000000
1!
1%
#188740000000
0!
0%
#188745000000
1!
1%
#188750000000
0!
0%
#188755000000
1!
1%
#188760000000
0!
0%
#188765000000
1!
1%
#188770000000
0!
0%
#188775000000
1!
1%
#188780000000
0!
0%
#188785000000
1!
1%
#188790000000
0!
0%
#188795000000
1!
1%
#188800000000
0!
0%
#188805000000
1!
1%
#188810000000
0!
0%
#188815000000
1!
1%
#188820000000
0!
0%
#188825000000
1!
1%
#188830000000
0!
0%
#188835000000
1!
1%
#188840000000
0!
0%
#188845000000
1!
1%
#188850000000
0!
0%
#188855000000
1!
1%
#188860000000
0!
0%
#188865000000
1!
1%
#188870000000
0!
0%
#188875000000
1!
1%
#188880000000
0!
0%
#188885000000
1!
1%
#188890000000
0!
0%
#188895000000
1!
1%
#188900000000
0!
0%
#188905000000
1!
1%
#188910000000
0!
0%
#188915000000
1!
1%
#188920000000
0!
0%
#188925000000
1!
1%
#188930000000
0!
0%
#188935000000
1!
1%
#188940000000
0!
0%
#188945000000
1!
1%
#188950000000
0!
0%
#188955000000
1!
1%
#188960000000
0!
0%
#188965000000
1!
1%
#188970000000
0!
0%
#188975000000
1!
1%
#188980000000
0!
0%
#188985000000
1!
1%
#188990000000
0!
0%
#188995000000
1!
1%
#189000000000
0!
0%
#189005000000
1!
1%
#189010000000
0!
0%
#189015000000
1!
1%
#189020000000
0!
0%
#189025000000
1!
1%
#189030000000
0!
0%
#189035000000
1!
1%
#189040000000
0!
0%
#189045000000
1!
1%
#189050000000
0!
0%
#189055000000
1!
1%
#189060000000
0!
0%
#189065000000
1!
1%
#189070000000
0!
0%
#189075000000
1!
1%
#189080000000
0!
0%
#189085000000
1!
1%
#189090000000
0!
0%
#189095000000
1!
1%
#189100000000
0!
0%
#189105000000
1!
1%
#189110000000
0!
0%
#189115000000
1!
1%
#189120000000
0!
0%
#189125000000
1!
1%
#189130000000
0!
0%
#189135000000
1!
1%
#189140000000
0!
0%
#189145000000
1!
1%
#189150000000
0!
0%
#189155000000
1!
1%
#189160000000
0!
0%
#189165000000
1!
1%
#189170000000
0!
0%
#189175000000
1!
1%
#189180000000
0!
0%
#189185000000
1!
1%
#189190000000
0!
0%
#189195000000
1!
1%
#189200000000
0!
0%
#189205000000
1!
1%
#189210000000
0!
0%
#189215000000
1!
1%
#189220000000
0!
0%
#189225000000
1!
1%
#189230000000
0!
0%
#189235000000
1!
1%
#189240000000
0!
0%
#189245000000
1!
1%
#189250000000
0!
0%
#189255000000
1!
1%
#189260000000
0!
0%
#189265000000
1!
1%
#189270000000
0!
0%
#189275000000
1!
1%
#189280000000
0!
0%
#189285000000
1!
1%
#189290000000
0!
0%
#189295000000
1!
1%
#189300000000
0!
0%
#189305000000
1!
1%
#189310000000
0!
0%
#189315000000
1!
1%
#189320000000
0!
0%
#189325000000
1!
1%
#189330000000
0!
0%
#189335000000
1!
1%
#189340000000
0!
0%
#189345000000
1!
1%
#189350000000
0!
0%
#189355000000
1!
1%
#189360000000
0!
0%
#189365000000
1!
1%
#189370000000
0!
0%
#189375000000
1!
1%
#189380000000
0!
0%
#189385000000
1!
1%
#189390000000
0!
0%
#189395000000
1!
1%
#189400000000
0!
0%
#189405000000
1!
1%
#189410000000
0!
0%
#189415000000
1!
1%
#189420000000
0!
0%
#189425000000
1!
1%
#189430000000
0!
0%
#189435000000
1!
1%
#189440000000
0!
0%
#189445000000
1!
1%
#189450000000
0!
0%
#189455000000
1!
1%
#189460000000
0!
0%
#189465000000
1!
1%
#189470000000
0!
0%
#189475000000
1!
1%
#189480000000
0!
0%
#189485000000
1!
1%
#189490000000
0!
0%
#189495000000
1!
1%
#189500000000
0!
0%
#189505000000
1!
1%
#189510000000
0!
0%
#189515000000
1!
1%
#189520000000
0!
0%
#189525000000
1!
1%
#189530000000
0!
0%
#189535000000
1!
1%
#189540000000
0!
0%
#189545000000
1!
1%
#189550000000
0!
0%
#189555000000
1!
1%
#189560000000
0!
0%
#189565000000
1!
1%
#189570000000
0!
0%
#189575000000
1!
1%
#189580000000
0!
0%
#189585000000
1!
1%
#189590000000
0!
0%
#189595000000
1!
1%
#189600000000
0!
0%
#189605000000
1!
1%
#189610000000
0!
0%
#189615000000
1!
1%
#189620000000
0!
0%
#189625000000
1!
1%
#189630000000
0!
0%
#189635000000
1!
1%
#189640000000
0!
0%
#189645000000
1!
1%
#189650000000
0!
0%
#189655000000
1!
1%
#189660000000
0!
0%
#189665000000
1!
1%
#189670000000
0!
0%
#189675000000
1!
1%
#189680000000
0!
0%
#189685000000
1!
1%
#189690000000
0!
0%
#189695000000
1!
1%
#189700000000
0!
0%
#189705000000
1!
1%
#189710000000
0!
0%
#189715000000
1!
1%
#189720000000
0!
0%
#189725000000
1!
1%
#189730000000
0!
0%
#189735000000
1!
1%
#189740000000
0!
0%
#189745000000
1!
1%
#189750000000
0!
0%
#189755000000
1!
1%
#189760000000
0!
0%
#189765000000
1!
1%
#189770000000
0!
0%
#189775000000
1!
1%
#189780000000
0!
0%
#189785000000
1!
1%
#189790000000
0!
0%
#189795000000
1!
1%
#189800000000
0!
0%
#189805000000
1!
1%
#189810000000
0!
0%
#189815000000
1!
1%
#189820000000
0!
0%
#189825000000
1!
1%
#189830000000
0!
0%
#189835000000
1!
1%
#189840000000
0!
0%
#189845000000
1!
1%
#189850000000
0!
0%
#189855000000
1!
1%
#189860000000
0!
0%
#189865000000
1!
1%
#189870000000
0!
0%
#189875000000
1!
1%
#189880000000
0!
0%
#189885000000
1!
1%
#189890000000
0!
0%
#189895000000
1!
1%
#189900000000
0!
0%
#189905000000
1!
1%
#189910000000
0!
0%
#189915000000
1!
1%
#189920000000
0!
0%
#189925000000
1!
1%
#189930000000
0!
0%
#189935000000
1!
1%
#189940000000
0!
0%
#189945000000
1!
1%
#189950000000
0!
0%
#189955000000
1!
1%
#189960000000
0!
0%
#189965000000
1!
1%
#189970000000
0!
0%
#189975000000
1!
1%
#189980000000
0!
0%
#189985000000
1!
1%
#189990000000
0!
0%
#189995000000
1!
1%
#190000000000
0!
0%
#190005000000
1!
1%
#190010000000
0!
0%
#190015000000
1!
1%
#190020000000
0!
0%
#190025000000
1!
1%
#190030000000
0!
0%
#190035000000
1!
1%
#190040000000
0!
0%
#190045000000
1!
1%
#190050000000
0!
0%
#190055000000
1!
1%
#190060000000
0!
0%
#190065000000
1!
1%
#190070000000
0!
0%
#190075000000
1!
1%
#190080000000
0!
0%
#190085000000
1!
1%
#190090000000
0!
0%
#190095000000
1!
1%
#190100000000
0!
0%
#190105000000
1!
1%
#190110000000
0!
0%
#190115000000
1!
1%
#190120000000
0!
0%
#190125000000
1!
1%
#190130000000
0!
0%
#190135000000
1!
1%
#190140000000
0!
0%
#190145000000
1!
1%
#190150000000
0!
0%
#190155000000
1!
1%
#190160000000
0!
0%
#190165000000
1!
1%
#190170000000
0!
0%
#190175000000
1!
1%
#190180000000
0!
0%
#190185000000
1!
1%
#190190000000
0!
0%
#190195000000
1!
1%
#190200000000
0!
0%
#190205000000
1!
1%
#190210000000
0!
0%
#190215000000
1!
1%
#190220000000
0!
0%
#190225000000
1!
1%
#190230000000
0!
0%
#190235000000
1!
1%
#190240000000
0!
0%
#190245000000
1!
1%
#190250000000
0!
0%
#190255000000
1!
1%
#190260000000
0!
0%
#190265000000
1!
1%
#190270000000
0!
0%
#190275000000
1!
1%
#190280000000
0!
0%
#190285000000
1!
1%
#190290000000
0!
0%
#190295000000
1!
1%
#190300000000
0!
0%
#190305000000
1!
1%
#190310000000
0!
0%
#190315000000
1!
1%
#190320000000
0!
0%
#190325000000
1!
1%
#190330000000
0!
0%
#190335000000
1!
1%
#190340000000
0!
0%
#190345000000
1!
1%
#190350000000
0!
0%
#190355000000
1!
1%
#190360000000
0!
0%
#190365000000
1!
1%
#190370000000
0!
0%
#190375000000
1!
1%
#190380000000
0!
0%
#190385000000
1!
1%
#190390000000
0!
0%
#190395000000
1!
1%
#190400000000
0!
0%
#190405000000
1!
1%
#190410000000
0!
0%
#190415000000
1!
1%
#190420000000
0!
0%
#190425000000
1!
1%
#190430000000
0!
0%
#190435000000
1!
1%
#190440000000
0!
0%
#190445000000
1!
1%
#190450000000
0!
0%
#190455000000
1!
1%
#190460000000
0!
0%
#190465000000
1!
1%
#190470000000
0!
0%
#190475000000
1!
1%
#190480000000
0!
0%
#190485000000
1!
1%
#190490000000
0!
0%
#190495000000
1!
1%
#190500000000
0!
0%
#190505000000
1!
1%
#190510000000
0!
0%
#190515000000
1!
1%
#190520000000
0!
0%
#190525000000
1!
1%
#190530000000
0!
0%
#190535000000
1!
1%
#190540000000
0!
0%
#190545000000
1!
1%
#190550000000
0!
0%
#190555000000
1!
1%
#190560000000
0!
0%
#190565000000
1!
1%
#190570000000
0!
0%
#190575000000
1!
1%
#190580000000
0!
0%
#190585000000
1!
1%
#190590000000
0!
0%
#190595000000
1!
1%
#190600000000
0!
0%
#190605000000
1!
1%
#190610000000
0!
0%
#190615000000
1!
1%
#190620000000
0!
0%
#190625000000
1!
1%
#190630000000
0!
0%
#190635000000
1!
1%
#190640000000
0!
0%
#190645000000
1!
1%
#190650000000
0!
0%
#190655000000
1!
1%
#190660000000
0!
0%
#190665000000
1!
1%
#190670000000
0!
0%
#190675000000
1!
1%
#190680000000
0!
0%
#190685000000
1!
1%
#190690000000
0!
0%
#190695000000
1!
1%
#190700000000
0!
0%
#190705000000
1!
1%
#190710000000
0!
0%
#190715000000
1!
1%
#190720000000
0!
0%
#190725000000
1!
1%
#190730000000
0!
0%
#190735000000
1!
1%
#190740000000
0!
0%
#190745000000
1!
1%
#190750000000
0!
0%
#190755000000
1!
1%
#190760000000
0!
0%
#190765000000
1!
1%
#190770000000
0!
0%
#190775000000
1!
1%
#190780000000
0!
0%
#190785000000
1!
1%
#190790000000
0!
0%
#190795000000
1!
1%
#190800000000
0!
0%
#190805000000
1!
1%
#190810000000
0!
0%
#190815000000
1!
1%
#190820000000
0!
0%
#190825000000
1!
1%
#190830000000
0!
0%
#190835000000
1!
1%
#190840000000
0!
0%
#190845000000
1!
1%
#190850000000
0!
0%
#190855000000
1!
1%
#190860000000
0!
0%
#190865000000
1!
1%
#190870000000
0!
0%
#190875000000
1!
1%
#190880000000
0!
0%
#190885000000
1!
1%
#190890000000
0!
0%
#190895000000
1!
1%
#190900000000
0!
0%
#190905000000
1!
1%
#190910000000
0!
0%
#190915000000
1!
1%
#190920000000
0!
0%
#190925000000
1!
1%
#190930000000
0!
0%
#190935000000
1!
1%
#190940000000
0!
0%
#190945000000
1!
1%
#190950000000
0!
0%
#190955000000
1!
1%
#190960000000
0!
0%
#190965000000
1!
1%
#190970000000
0!
0%
#190975000000
1!
1%
#190980000000
0!
0%
#190985000000
1!
1%
#190990000000
0!
0%
#190995000000
1!
1%
#191000000000
0!
0%
#191005000000
1!
1%
#191010000000
0!
0%
#191015000000
1!
1%
#191020000000
0!
0%
#191025000000
1!
1%
#191030000000
0!
0%
#191035000000
1!
1%
#191040000000
0!
0%
#191045000000
1!
1%
#191050000000
0!
0%
#191055000000
1!
1%
#191060000000
0!
0%
#191065000000
1!
1%
#191070000000
0!
0%
#191075000000
1!
1%
#191080000000
0!
0%
#191085000000
1!
1%
#191090000000
0!
0%
#191095000000
1!
1%
#191100000000
0!
0%
#191105000000
1!
1%
#191110000000
0!
0%
#191115000000
1!
1%
#191120000000
0!
0%
#191125000000
1!
1%
#191130000000
0!
0%
#191135000000
1!
1%
#191140000000
0!
0%
#191145000000
1!
1%
#191150000000
0!
0%
#191155000000
1!
1%
#191160000000
0!
0%
#191165000000
1!
1%
#191170000000
0!
0%
#191175000000
1!
1%
#191180000000
0!
0%
#191185000000
1!
1%
#191190000000
0!
0%
#191195000000
1!
1%
#191200000000
0!
0%
#191205000000
1!
1%
#191210000000
0!
0%
#191215000000
1!
1%
#191220000000
0!
0%
#191225000000
1!
1%
#191230000000
0!
0%
#191235000000
1!
1%
#191240000000
0!
0%
#191245000000
1!
1%
#191250000000
0!
0%
#191255000000
1!
1%
#191260000000
0!
0%
#191265000000
1!
1%
#191270000000
0!
0%
#191275000000
1!
1%
#191280000000
0!
0%
#191285000000
1!
1%
#191290000000
0!
0%
#191295000000
1!
1%
#191300000000
0!
0%
#191305000000
1!
1%
#191310000000
0!
0%
#191315000000
1!
1%
#191320000000
0!
0%
#191325000000
1!
1%
#191330000000
0!
0%
#191335000000
1!
1%
#191340000000
0!
0%
#191345000000
1!
1%
#191350000000
0!
0%
#191355000000
1!
1%
#191360000000
0!
0%
#191365000000
1!
1%
#191370000000
0!
0%
#191375000000
1!
1%
#191380000000
0!
0%
#191385000000
1!
1%
#191390000000
0!
0%
#191395000000
1!
1%
#191400000000
0!
0%
#191405000000
1!
1%
#191410000000
0!
0%
#191415000000
1!
1%
#191420000000
0!
0%
#191425000000
1!
1%
#191430000000
0!
0%
#191435000000
1!
1%
#191440000000
0!
0%
#191445000000
1!
1%
#191450000000
0!
0%
#191455000000
1!
1%
#191460000000
0!
0%
#191465000000
1!
1%
#191470000000
0!
0%
#191475000000
1!
1%
#191480000000
0!
0%
#191485000000
1!
1%
#191490000000
0!
0%
#191495000000
1!
1%
#191500000000
0!
0%
#191505000000
1!
1%
#191510000000
0!
0%
#191515000000
1!
1%
#191520000000
0!
0%
#191525000000
1!
1%
#191530000000
0!
0%
#191535000000
1!
1%
#191540000000
0!
0%
#191545000000
1!
1%
#191550000000
0!
0%
#191555000000
1!
1%
#191560000000
0!
0%
#191565000000
1!
1%
#191570000000
0!
0%
#191575000000
1!
1%
#191580000000
0!
0%
#191585000000
1!
1%
#191590000000
0!
0%
#191595000000
1!
1%
#191600000000
0!
0%
#191605000000
1!
1%
#191610000000
0!
0%
#191615000000
1!
1%
#191620000000
0!
0%
#191625000000
1!
1%
#191630000000
0!
0%
#191635000000
1!
1%
#191640000000
0!
0%
#191645000000
1!
1%
#191650000000
0!
0%
#191655000000
1!
1%
#191660000000
0!
0%
#191665000000
1!
1%
#191670000000
0!
0%
#191675000000
1!
1%
#191680000000
0!
0%
#191685000000
1!
1%
#191690000000
0!
0%
#191695000000
1!
1%
#191700000000
0!
0%
#191705000000
1!
1%
#191710000000
0!
0%
#191715000000
1!
1%
#191720000000
0!
0%
#191725000000
1!
1%
#191730000000
0!
0%
#191735000000
1!
1%
#191740000000
0!
0%
#191745000000
1!
1%
#191750000000
0!
0%
#191755000000
1!
1%
#191760000000
0!
0%
#191765000000
1!
1%
#191770000000
0!
0%
#191775000000
1!
1%
#191780000000
0!
0%
#191785000000
1!
1%
#191790000000
0!
0%
#191795000000
1!
1%
#191800000000
0!
0%
#191805000000
1!
1%
#191810000000
0!
0%
#191815000000
1!
1%
#191820000000
0!
0%
#191825000000
1!
1%
#191830000000
0!
0%
#191835000000
1!
1%
#191840000000
0!
0%
#191845000000
1!
1%
#191850000000
0!
0%
#191855000000
1!
1%
#191860000000
0!
0%
#191865000000
1!
1%
#191870000000
0!
0%
#191875000000
1!
1%
#191880000000
0!
0%
#191885000000
1!
1%
#191890000000
0!
0%
#191895000000
1!
1%
#191900000000
0!
0%
#191905000000
1!
1%
#191910000000
0!
0%
#191915000000
1!
1%
#191920000000
0!
0%
#191925000000
1!
1%
#191930000000
0!
0%
#191935000000
1!
1%
#191940000000
0!
0%
#191945000000
1!
1%
#191950000000
0!
0%
#191955000000
1!
1%
#191960000000
0!
0%
#191965000000
1!
1%
#191970000000
0!
0%
#191975000000
1!
1%
#191980000000
0!
0%
#191985000000
1!
1%
#191990000000
0!
0%
#191995000000
1!
1%
#192000000000
0!
0%
#192005000000
1!
1%
#192010000000
0!
0%
#192015000000
1!
1%
#192020000000
0!
0%
#192025000000
1!
1%
#192030000000
0!
0%
#192035000000
1!
1%
#192040000000
0!
0%
#192045000000
1!
1%
#192050000000
0!
0%
#192055000000
1!
1%
#192060000000
0!
0%
#192065000000
1!
1%
#192070000000
0!
0%
#192075000000
1!
1%
#192080000000
0!
0%
#192085000000
1!
1%
#192090000000
0!
0%
#192095000000
1!
1%
#192100000000
0!
0%
#192105000000
1!
1%
#192110000000
0!
0%
#192115000000
1!
1%
#192120000000
0!
0%
#192125000000
1!
1%
#192130000000
0!
0%
#192135000000
1!
1%
#192140000000
0!
0%
#192145000000
1!
1%
#192150000000
0!
0%
#192155000000
1!
1%
#192160000000
0!
0%
#192165000000
1!
1%
#192170000000
0!
0%
#192175000000
1!
1%
#192180000000
0!
0%
#192185000000
1!
1%
#192190000000
0!
0%
#192195000000
1!
1%
#192200000000
0!
0%
#192205000000
1!
1%
#192210000000
0!
0%
#192215000000
1!
1%
#192220000000
0!
0%
#192225000000
1!
1%
#192230000000
0!
0%
#192235000000
1!
1%
#192240000000
0!
0%
#192245000000
1!
1%
#192250000000
0!
0%
#192255000000
1!
1%
#192260000000
0!
0%
#192265000000
1!
1%
#192270000000
0!
0%
#192275000000
1!
1%
#192280000000
0!
0%
#192285000000
1!
1%
#192290000000
0!
0%
#192295000000
1!
1%
#192300000000
0!
0%
#192305000000
1!
1%
#192310000000
0!
0%
#192315000000
1!
1%
#192320000000
0!
0%
#192325000000
1!
1%
#192330000000
0!
0%
#192335000000
1!
1%
#192340000000
0!
0%
#192345000000
1!
1%
#192350000000
0!
0%
#192355000000
1!
1%
#192360000000
0!
0%
#192365000000
1!
1%
#192370000000
0!
0%
#192375000000
1!
1%
#192380000000
0!
0%
#192385000000
1!
1%
#192390000000
0!
0%
#192395000000
1!
1%
#192400000000
0!
0%
#192405000000
1!
1%
#192410000000
0!
0%
#192415000000
1!
1%
#192420000000
0!
0%
#192425000000
1!
1%
#192430000000
0!
0%
#192435000000
1!
1%
#192440000000
0!
0%
#192445000000
1!
1%
#192450000000
0!
0%
#192455000000
1!
1%
#192460000000
0!
0%
#192465000000
1!
1%
#192470000000
0!
0%
#192475000000
1!
1%
#192480000000
0!
0%
#192485000000
1!
1%
#192490000000
0!
0%
#192495000000
1!
1%
#192500000000
0!
0%
#192505000000
1!
1%
#192510000000
0!
0%
#192515000000
1!
1%
#192520000000
0!
0%
#192525000000
1!
1%
#192530000000
0!
0%
#192535000000
1!
1%
#192540000000
0!
0%
#192545000000
1!
1%
#192550000000
0!
0%
#192555000000
1!
1%
#192560000000
0!
0%
#192565000000
1!
1%
#192570000000
0!
0%
#192575000000
1!
1%
#192580000000
0!
0%
#192585000000
1!
1%
#192590000000
0!
0%
#192595000000
1!
1%
#192600000000
0!
0%
#192605000000
1!
1%
#192610000000
0!
0%
#192615000000
1!
1%
#192620000000
0!
0%
#192625000000
1!
1%
#192630000000
0!
0%
#192635000000
1!
1%
#192640000000
0!
0%
#192645000000
1!
1%
#192650000000
0!
0%
#192655000000
1!
1%
#192660000000
0!
0%
#192665000000
1!
1%
#192670000000
0!
0%
#192675000000
1!
1%
#192680000000
0!
0%
#192685000000
1!
1%
#192690000000
0!
0%
#192695000000
1!
1%
#192700000000
0!
0%
#192705000000
1!
1%
#192710000000
0!
0%
#192715000000
1!
1%
#192720000000
0!
0%
#192725000000
1!
1%
#192730000000
0!
0%
#192735000000
1!
1%
#192740000000
0!
0%
#192745000000
1!
1%
#192750000000
0!
0%
#192755000000
1!
1%
#192760000000
0!
0%
#192765000000
1!
1%
#192770000000
0!
0%
#192775000000
1!
1%
#192780000000
0!
0%
#192785000000
1!
1%
#192790000000
0!
0%
#192795000000
1!
1%
#192800000000
0!
0%
#192805000000
1!
1%
#192810000000
0!
0%
#192815000000
1!
1%
#192820000000
0!
0%
#192825000000
1!
1%
#192830000000
0!
0%
#192835000000
1!
1%
#192840000000
0!
0%
#192845000000
1!
1%
#192850000000
0!
0%
#192855000000
1!
1%
#192860000000
0!
0%
#192865000000
1!
1%
#192870000000
0!
0%
#192875000000
1!
1%
#192880000000
0!
0%
#192885000000
1!
1%
#192890000000
0!
0%
#192895000000
1!
1%
#192900000000
0!
0%
#192905000000
1!
1%
#192910000000
0!
0%
#192915000000
1!
1%
#192920000000
0!
0%
#192925000000
1!
1%
#192930000000
0!
0%
#192935000000
1!
1%
#192940000000
0!
0%
#192945000000
1!
1%
#192950000000
0!
0%
#192955000000
1!
1%
#192960000000
0!
0%
#192965000000
1!
1%
#192970000000
0!
0%
#192975000000
1!
1%
#192980000000
0!
0%
#192985000000
1!
1%
#192990000000
0!
0%
#192995000000
1!
1%
#193000000000
0!
0%
#193005000000
1!
1%
#193010000000
0!
0%
#193015000000
1!
1%
#193020000000
0!
0%
#193025000000
1!
1%
#193030000000
0!
0%
#193035000000
1!
1%
#193040000000
0!
0%
#193045000000
1!
1%
#193050000000
0!
0%
#193055000000
1!
1%
#193060000000
0!
0%
#193065000000
1!
1%
#193070000000
0!
0%
#193075000000
1!
1%
#193080000000
0!
0%
#193085000000
1!
1%
#193090000000
0!
0%
#193095000000
1!
1%
#193100000000
0!
0%
#193105000000
1!
1%
#193110000000
0!
0%
#193115000000
1!
1%
#193120000000
0!
0%
#193125000000
1!
1%
#193130000000
0!
0%
#193135000000
1!
1%
#193140000000
0!
0%
#193145000000
1!
1%
#193150000000
0!
0%
#193155000000
1!
1%
#193160000000
0!
0%
#193165000000
1!
1%
#193170000000
0!
0%
#193175000000
1!
1%
#193180000000
0!
0%
#193185000000
1!
1%
#193190000000
0!
0%
#193195000000
1!
1%
#193200000000
0!
0%
#193205000000
1!
1%
#193210000000
0!
0%
#193215000000
1!
1%
#193220000000
0!
0%
#193225000000
1!
1%
#193230000000
0!
0%
#193235000000
1!
1%
#193240000000
0!
0%
#193245000000
1!
1%
#193250000000
0!
0%
#193255000000
1!
1%
#193260000000
0!
0%
#193265000000
1!
1%
#193270000000
0!
0%
#193275000000
1!
1%
#193280000000
0!
0%
#193285000000
1!
1%
#193290000000
0!
0%
#193295000000
1!
1%
#193300000000
0!
0%
#193305000000
1!
1%
#193310000000
0!
0%
#193315000000
1!
1%
#193320000000
0!
0%
#193325000000
1!
1%
#193330000000
0!
0%
#193335000000
1!
1%
#193340000000
0!
0%
#193345000000
1!
1%
#193350000000
0!
0%
#193355000000
1!
1%
#193360000000
0!
0%
#193365000000
1!
1%
#193370000000
0!
0%
#193375000000
1!
1%
#193380000000
0!
0%
#193385000000
1!
1%
#193390000000
0!
0%
#193395000000
1!
1%
#193400000000
0!
0%
#193405000000
1!
1%
#193410000000
0!
0%
#193415000000
1!
1%
#193420000000
0!
0%
#193425000000
1!
1%
#193430000000
0!
0%
#193435000000
1!
1%
#193440000000
0!
0%
#193445000000
1!
1%
#193450000000
0!
0%
#193455000000
1!
1%
#193460000000
0!
0%
#193465000000
1!
1%
#193470000000
0!
0%
#193475000000
1!
1%
#193480000000
0!
0%
#193485000000
1!
1%
#193490000000
0!
0%
#193495000000
1!
1%
#193500000000
0!
0%
#193505000000
1!
1%
#193510000000
0!
0%
#193515000000
1!
1%
#193520000000
0!
0%
#193525000000
1!
1%
#193530000000
0!
0%
#193535000000
1!
1%
#193540000000
0!
0%
#193545000000
1!
1%
#193550000000
0!
0%
#193555000000
1!
1%
#193560000000
0!
0%
#193565000000
1!
1%
#193570000000
0!
0%
#193575000000
1!
1%
#193580000000
0!
0%
#193585000000
1!
1%
#193590000000
0!
0%
#193595000000
1!
1%
#193600000000
0!
0%
#193605000000
1!
1%
#193610000000
0!
0%
#193615000000
1!
1%
#193620000000
0!
0%
#193625000000
1!
1%
#193630000000
0!
0%
#193635000000
1!
1%
#193640000000
0!
0%
#193645000000
1!
1%
#193650000000
0!
0%
#193655000000
1!
1%
#193660000000
0!
0%
#193665000000
1!
1%
#193670000000
0!
0%
#193675000000
1!
1%
#193680000000
0!
0%
#193685000000
1!
1%
#193690000000
0!
0%
#193695000000
1!
1%
#193700000000
0!
0%
#193705000000
1!
1%
#193710000000
0!
0%
#193715000000
1!
1%
#193720000000
0!
0%
#193725000000
1!
1%
#193730000000
0!
0%
#193735000000
1!
1%
#193740000000
0!
0%
#193745000000
1!
1%
#193750000000
0!
0%
#193755000000
1!
1%
#193760000000
0!
0%
#193765000000
1!
1%
#193770000000
0!
0%
#193775000000
1!
1%
#193780000000
0!
0%
#193785000000
1!
1%
#193790000000
0!
0%
#193795000000
1!
1%
#193800000000
0!
0%
#193805000000
1!
1%
#193810000000
0!
0%
#193815000000
1!
1%
#193820000000
0!
0%
#193825000000
1!
1%
#193830000000
0!
0%
#193835000000
1!
1%
#193840000000
0!
0%
#193845000000
1!
1%
#193850000000
0!
0%
#193855000000
1!
1%
#193860000000
0!
0%
#193865000000
1!
1%
#193870000000
0!
0%
#193875000000
1!
1%
#193880000000
0!
0%
#193885000000
1!
1%
#193890000000
0!
0%
#193895000000
1!
1%
#193900000000
0!
0%
#193905000000
1!
1%
#193910000000
0!
0%
#193915000000
1!
1%
#193920000000
0!
0%
#193925000000
1!
1%
#193930000000
0!
0%
#193935000000
1!
1%
#193940000000
0!
0%
#193945000000
1!
1%
#193950000000
0!
0%
#193955000000
1!
1%
#193960000000
0!
0%
#193965000000
1!
1%
#193970000000
0!
0%
#193975000000
1!
1%
#193980000000
0!
0%
#193985000000
1!
1%
#193990000000
0!
0%
#193995000000
1!
1%
#194000000000
0!
0%
#194005000000
1!
1%
#194010000000
0!
0%
#194015000000
1!
1%
#194020000000
0!
0%
#194025000000
1!
1%
#194030000000
0!
0%
#194035000000
1!
1%
#194040000000
0!
0%
#194045000000
1!
1%
#194050000000
0!
0%
#194055000000
1!
1%
#194060000000
0!
0%
#194065000000
1!
1%
#194070000000
0!
0%
#194075000000
1!
1%
#194080000000
0!
0%
#194085000000
1!
1%
#194090000000
0!
0%
#194095000000
1!
1%
#194100000000
0!
0%
#194105000000
1!
1%
#194110000000
0!
0%
#194115000000
1!
1%
#194120000000
0!
0%
#194125000000
1!
1%
#194130000000
0!
0%
#194135000000
1!
1%
#194140000000
0!
0%
#194145000000
1!
1%
#194150000000
0!
0%
#194155000000
1!
1%
#194160000000
0!
0%
#194165000000
1!
1%
#194170000000
0!
0%
#194175000000
1!
1%
#194180000000
0!
0%
#194185000000
1!
1%
#194190000000
0!
0%
#194195000000
1!
1%
#194200000000
0!
0%
#194205000000
1!
1%
#194210000000
0!
0%
#194215000000
1!
1%
#194220000000
0!
0%
#194225000000
1!
1%
#194230000000
0!
0%
#194235000000
1!
1%
#194240000000
0!
0%
#194245000000
1!
1%
#194250000000
0!
0%
#194255000000
1!
1%
#194260000000
0!
0%
#194265000000
1!
1%
#194270000000
0!
0%
#194275000000
1!
1%
#194280000000
0!
0%
#194285000000
1!
1%
#194290000000
0!
0%
#194295000000
1!
1%
#194300000000
0!
0%
#194305000000
1!
1%
#194310000000
0!
0%
#194315000000
1!
1%
#194320000000
0!
0%
#194325000000
1!
1%
#194330000000
0!
0%
#194335000000
1!
1%
#194340000000
0!
0%
#194345000000
1!
1%
#194350000000
0!
0%
#194355000000
1!
1%
#194360000000
0!
0%
#194365000000
1!
1%
#194370000000
0!
0%
#194375000000
1!
1%
#194380000000
0!
0%
#194385000000
1!
1%
#194390000000
0!
0%
#194395000000
1!
1%
#194400000000
0!
0%
#194405000000
1!
1%
#194410000000
0!
0%
#194415000000
1!
1%
#194420000000
0!
0%
#194425000000
1!
1%
#194430000000
0!
0%
#194435000000
1!
1%
#194440000000
0!
0%
#194445000000
1!
1%
#194450000000
0!
0%
#194455000000
1!
1%
#194460000000
0!
0%
#194465000000
1!
1%
#194470000000
0!
0%
#194475000000
1!
1%
#194480000000
0!
0%
#194485000000
1!
1%
#194490000000
0!
0%
#194495000000
1!
1%
#194500000000
0!
0%
#194505000000
1!
1%
#194510000000
0!
0%
#194515000000
1!
1%
#194520000000
0!
0%
#194525000000
1!
1%
#194530000000
0!
0%
#194535000000
1!
1%
#194540000000
0!
0%
#194545000000
1!
1%
#194550000000
0!
0%
#194555000000
1!
1%
#194560000000
0!
0%
#194565000000
1!
1%
#194570000000
0!
0%
#194575000000
1!
1%
#194580000000
0!
0%
#194585000000
1!
1%
#194590000000
0!
0%
#194595000000
1!
1%
#194600000000
0!
0%
#194605000000
1!
1%
#194610000000
0!
0%
#194615000000
1!
1%
#194620000000
0!
0%
#194625000000
1!
1%
#194630000000
0!
0%
#194635000000
1!
1%
#194640000000
0!
0%
#194645000000
1!
1%
#194650000000
0!
0%
#194655000000
1!
1%
#194660000000
0!
0%
#194665000000
1!
1%
#194670000000
0!
0%
#194675000000
1!
1%
#194680000000
0!
0%
#194685000000
1!
1%
#194690000000
0!
0%
#194695000000
1!
1%
#194700000000
0!
0%
#194705000000
1!
1%
#194710000000
0!
0%
#194715000000
1!
1%
#194720000000
0!
0%
#194725000000
1!
1%
#194730000000
0!
0%
#194735000000
1!
1%
#194740000000
0!
0%
#194745000000
1!
1%
#194750000000
0!
0%
#194755000000
1!
1%
#194760000000
0!
0%
#194765000000
1!
1%
#194770000000
0!
0%
#194775000000
1!
1%
#194780000000
0!
0%
#194785000000
1!
1%
#194790000000
0!
0%
#194795000000
1!
1%
#194800000000
0!
0%
#194805000000
1!
1%
#194810000000
0!
0%
#194815000000
1!
1%
#194820000000
0!
0%
#194825000000
1!
1%
#194830000000
0!
0%
#194835000000
1!
1%
#194840000000
0!
0%
#194845000000
1!
1%
#194850000000
0!
0%
#194855000000
1!
1%
#194860000000
0!
0%
#194865000000
1!
1%
#194870000000
0!
0%
#194875000000
1!
1%
#194880000000
0!
0%
#194885000000
1!
1%
#194890000000
0!
0%
#194895000000
1!
1%
#194900000000
0!
0%
#194905000000
1!
1%
#194910000000
0!
0%
#194915000000
1!
1%
#194920000000
0!
0%
#194925000000
1!
1%
#194930000000
0!
0%
#194935000000
1!
1%
#194940000000
0!
0%
#194945000000
1!
1%
#194950000000
0!
0%
#194955000000
1!
1%
#194960000000
0!
0%
#194965000000
1!
1%
#194970000000
0!
0%
#194975000000
1!
1%
#194980000000
0!
0%
#194985000000
1!
1%
#194990000000
0!
0%
#194995000000
1!
1%
#195000000000
0!
0%
#195005000000
1!
1%
#195010000000
0!
0%
#195015000000
1!
1%
#195020000000
0!
0%
#195025000000
1!
1%
#195030000000
0!
0%
#195035000000
1!
1%
#195040000000
0!
0%
#195045000000
1!
1%
#195050000000
0!
0%
#195055000000
1!
1%
#195060000000
0!
0%
#195065000000
1!
1%
#195070000000
0!
0%
#195075000000
1!
1%
#195080000000
0!
0%
#195085000000
1!
1%
#195090000000
0!
0%
#195095000000
1!
1%
#195100000000
0!
0%
#195105000000
1!
1%
#195110000000
0!
0%
#195115000000
1!
1%
#195120000000
0!
0%
#195125000000
1!
1%
#195130000000
0!
0%
#195135000000
1!
1%
#195140000000
0!
0%
#195145000000
1!
1%
#195150000000
0!
0%
#195155000000
1!
1%
#195160000000
0!
0%
#195165000000
1!
1%
#195170000000
0!
0%
#195175000000
1!
1%
#195180000000
0!
0%
#195185000000
1!
1%
#195190000000
0!
0%
#195195000000
1!
1%
#195200000000
0!
0%
#195205000000
1!
1%
#195210000000
0!
0%
#195215000000
1!
1%
#195220000000
0!
0%
#195225000000
1!
1%
#195230000000
0!
0%
#195235000000
1!
1%
#195240000000
0!
0%
#195245000000
1!
1%
#195250000000
0!
0%
#195255000000
1!
1%
#195260000000
0!
0%
#195265000000
1!
1%
#195270000000
0!
0%
#195275000000
1!
1%
#195280000000
0!
0%
#195285000000
1!
1%
#195290000000
0!
0%
#195295000000
1!
1%
#195300000000
0!
0%
#195305000000
1!
1%
#195310000000
0!
0%
#195315000000
1!
1%
#195320000000
0!
0%
#195325000000
1!
1%
#195330000000
0!
0%
#195335000000
1!
1%
#195340000000
0!
0%
#195345000000
1!
1%
#195350000000
0!
0%
#195355000000
1!
1%
#195360000000
0!
0%
#195365000000
1!
1%
#195370000000
0!
0%
#195375000000
1!
1%
#195380000000
0!
0%
#195385000000
1!
1%
#195390000000
0!
0%
#195395000000
1!
1%
#195400000000
0!
0%
#195405000000
1!
1%
#195410000000
0!
0%
#195415000000
1!
1%
#195420000000
0!
0%
#195425000000
1!
1%
#195430000000
0!
0%
#195435000000
1!
1%
#195440000000
0!
0%
#195445000000
1!
1%
#195450000000
0!
0%
#195455000000
1!
1%
#195460000000
0!
0%
#195465000000
1!
1%
#195470000000
0!
0%
#195475000000
1!
1%
#195480000000
0!
0%
#195485000000
1!
1%
#195490000000
0!
0%
#195495000000
1!
1%
#195500000000
0!
0%
#195505000000
1!
1%
#195510000000
0!
0%
#195515000000
1!
1%
#195520000000
0!
0%
#195525000000
1!
1%
#195530000000
0!
0%
#195535000000
1!
1%
#195540000000
0!
0%
#195545000000
1!
1%
#195550000000
0!
0%
#195555000000
1!
1%
#195560000000
0!
0%
#195565000000
1!
1%
#195570000000
0!
0%
#195575000000
1!
1%
#195580000000
0!
0%
#195585000000
1!
1%
#195590000000
0!
0%
#195595000000
1!
1%
#195600000000
0!
0%
#195605000000
1!
1%
#195610000000
0!
0%
#195615000000
1!
1%
#195620000000
0!
0%
#195625000000
1!
1%
#195630000000
0!
0%
#195635000000
1!
1%
#195640000000
0!
0%
#195645000000
1!
1%
#195650000000
0!
0%
#195655000000
1!
1%
#195660000000
0!
0%
#195665000000
1!
1%
#195670000000
0!
0%
#195675000000
1!
1%
#195680000000
0!
0%
#195685000000
1!
1%
#195690000000
0!
0%
#195695000000
1!
1%
#195700000000
0!
0%
#195705000000
1!
1%
#195710000000
0!
0%
#195715000000
1!
1%
#195720000000
0!
0%
#195725000000
1!
1%
#195730000000
0!
0%
#195735000000
1!
1%
#195740000000
0!
0%
#195745000000
1!
1%
#195750000000
0!
0%
#195755000000
1!
1%
#195760000000
0!
0%
#195765000000
1!
1%
#195770000000
0!
0%
#195775000000
1!
1%
#195780000000
0!
0%
#195785000000
1!
1%
#195790000000
0!
0%
#195795000000
1!
1%
#195800000000
0!
0%
#195805000000
1!
1%
#195810000000
0!
0%
#195815000000
1!
1%
#195820000000
0!
0%
#195825000000
1!
1%
#195830000000
0!
0%
#195835000000
1!
1%
#195840000000
0!
0%
#195845000000
1!
1%
#195850000000
0!
0%
#195855000000
1!
1%
#195860000000
0!
0%
#195865000000
1!
1%
#195870000000
0!
0%
#195875000000
1!
1%
#195880000000
0!
0%
#195885000000
1!
1%
#195890000000
0!
0%
#195895000000
1!
1%
#195900000000
0!
0%
#195905000000
1!
1%
#195910000000
0!
0%
#195915000000
1!
1%
#195920000000
0!
0%
#195925000000
1!
1%
#195930000000
0!
0%
#195935000000
1!
1%
#195940000000
0!
0%
#195945000000
1!
1%
#195950000000
0!
0%
#195955000000
1!
1%
#195960000000
0!
0%
#195965000000
1!
1%
#195970000000
0!
0%
#195975000000
1!
1%
#195980000000
0!
0%
#195985000000
1!
1%
#195990000000
0!
0%
#195995000000
1!
1%
#196000000000
0!
0%
#196005000000
1!
1%
#196010000000
0!
0%
#196015000000
1!
1%
#196020000000
0!
0%
#196025000000
1!
1%
#196030000000
0!
0%
#196035000000
1!
1%
#196040000000
0!
0%
#196045000000
1!
1%
#196050000000
0!
0%
#196055000000
1!
1%
#196060000000
0!
0%
#196065000000
1!
1%
#196070000000
0!
0%
#196075000000
1!
1%
#196080000000
0!
0%
#196085000000
1!
1%
#196090000000
0!
0%
#196095000000
1!
1%
#196100000000
0!
0%
#196105000000
1!
1%
#196110000000
0!
0%
#196115000000
1!
1%
#196120000000
0!
0%
#196125000000
1!
1%
#196130000000
0!
0%
#196135000000
1!
1%
#196140000000
0!
0%
#196145000000
1!
1%
#196150000000
0!
0%
#196155000000
1!
1%
#196160000000
0!
0%
#196165000000
1!
1%
#196170000000
0!
0%
#196175000000
1!
1%
#196180000000
0!
0%
#196185000000
1!
1%
#196190000000
0!
0%
#196195000000
1!
1%
#196200000000
0!
0%
#196205000000
1!
1%
#196210000000
0!
0%
#196215000000
1!
1%
#196220000000
0!
0%
#196225000000
1!
1%
#196230000000
0!
0%
#196235000000
1!
1%
#196240000000
0!
0%
#196245000000
1!
1%
#196250000000
0!
0%
#196255000000
1!
1%
#196260000000
0!
0%
#196265000000
1!
1%
#196270000000
0!
0%
#196275000000
1!
1%
#196280000000
0!
0%
#196285000000
1!
1%
#196290000000
0!
0%
#196295000000
1!
1%
#196300000000
0!
0%
#196305000000
1!
1%
#196310000000
0!
0%
#196315000000
1!
1%
#196320000000
0!
0%
#196325000000
1!
1%
#196330000000
0!
0%
#196335000000
1!
1%
#196340000000
0!
0%
#196345000000
1!
1%
#196350000000
0!
0%
#196355000000
1!
1%
#196360000000
0!
0%
#196365000000
1!
1%
#196370000000
0!
0%
#196375000000
1!
1%
#196380000000
0!
0%
#196385000000
1!
1%
#196390000000
0!
0%
#196395000000
1!
1%
#196400000000
0!
0%
#196405000000
1!
1%
#196410000000
0!
0%
#196415000000
1!
1%
#196420000000
0!
0%
#196425000000
1!
1%
#196430000000
0!
0%
#196435000000
1!
1%
#196440000000
0!
0%
#196445000000
1!
1%
#196450000000
0!
0%
#196455000000
1!
1%
#196460000000
0!
0%
#196465000000
1!
1%
#196470000000
0!
0%
#196475000000
1!
1%
#196480000000
0!
0%
#196485000000
1!
1%
#196490000000
0!
0%
#196495000000
1!
1%
#196500000000
0!
0%
#196505000000
1!
1%
#196510000000
0!
0%
#196515000000
1!
1%
#196520000000
0!
0%
#196525000000
1!
1%
#196530000000
0!
0%
#196535000000
1!
1%
#196540000000
0!
0%
#196545000000
1!
1%
#196550000000
0!
0%
#196555000000
1!
1%
#196560000000
0!
0%
#196565000000
1!
1%
#196570000000
0!
0%
#196575000000
1!
1%
#196580000000
0!
0%
#196585000000
1!
1%
#196590000000
0!
0%
#196595000000
1!
1%
#196600000000
0!
0%
#196605000000
1!
1%
#196610000000
0!
0%
#196615000000
1!
1%
#196620000000
0!
0%
#196625000000
1!
1%
#196630000000
0!
0%
#196635000000
1!
1%
#196640000000
0!
0%
#196645000000
1!
1%
#196650000000
0!
0%
#196655000000
1!
1%
#196660000000
0!
0%
#196665000000
1!
1%
#196670000000
0!
0%
#196675000000
1!
1%
#196680000000
0!
0%
#196685000000
1!
1%
#196690000000
0!
0%
#196695000000
1!
1%
#196700000000
0!
0%
#196705000000
1!
1%
#196710000000
0!
0%
#196715000000
1!
1%
#196720000000
0!
0%
#196725000000
1!
1%
#196730000000
0!
0%
#196735000000
1!
1%
#196740000000
0!
0%
#196745000000
1!
1%
#196750000000
0!
0%
#196755000000
1!
1%
#196760000000
0!
0%
#196765000000
1!
1%
#196770000000
0!
0%
#196775000000
1!
1%
#196780000000
0!
0%
#196785000000
1!
1%
#196790000000
0!
0%
#196795000000
1!
1%
#196800000000
0!
0%
#196805000000
1!
1%
#196810000000
0!
0%
#196815000000
1!
1%
#196820000000
0!
0%
#196825000000
1!
1%
#196830000000
0!
0%
#196835000000
1!
1%
#196840000000
0!
0%
#196845000000
1!
1%
#196850000000
0!
0%
#196855000000
1!
1%
#196860000000
0!
0%
#196865000000
1!
1%
#196870000000
0!
0%
#196875000000
1!
1%
#196880000000
0!
0%
#196885000000
1!
1%
#196890000000
0!
0%
#196895000000
1!
1%
#196900000000
0!
0%
#196905000000
1!
1%
#196910000000
0!
0%
#196915000000
1!
1%
#196920000000
0!
0%
#196925000000
1!
1%
#196930000000
0!
0%
#196935000000
1!
1%
#196940000000
0!
0%
#196945000000
1!
1%
#196950000000
0!
0%
#196955000000
1!
1%
#196960000000
0!
0%
#196965000000
1!
1%
#196970000000
0!
0%
#196975000000
1!
1%
#196980000000
0!
0%
#196985000000
1!
1%
#196990000000
0!
0%
#196995000000
1!
1%
#197000000000
0!
0%
#197005000000
1!
1%
#197010000000
0!
0%
#197015000000
1!
1%
#197020000000
0!
0%
#197025000000
1!
1%
#197030000000
0!
0%
#197035000000
1!
1%
#197040000000
0!
0%
#197045000000
1!
1%
#197050000000
0!
0%
#197055000000
1!
1%
#197060000000
0!
0%
#197065000000
1!
1%
#197070000000
0!
0%
#197075000000
1!
1%
#197080000000
0!
0%
#197085000000
1!
1%
#197090000000
0!
0%
#197095000000
1!
1%
#197100000000
0!
0%
#197105000000
1!
1%
#197110000000
0!
0%
#197115000000
1!
1%
#197120000000
0!
0%
#197125000000
1!
1%
#197130000000
0!
0%
#197135000000
1!
1%
#197140000000
0!
0%
#197145000000
1!
1%
#197150000000
0!
0%
#197155000000
1!
1%
#197160000000
0!
0%
#197165000000
1!
1%
#197170000000
0!
0%
#197175000000
1!
1%
#197180000000
0!
0%
#197185000000
1!
1%
#197190000000
0!
0%
#197195000000
1!
1%
#197200000000
0!
0%
#197205000000
1!
1%
#197210000000
0!
0%
#197215000000
1!
1%
#197220000000
0!
0%
#197225000000
1!
1%
#197230000000
0!
0%
#197235000000
1!
1%
#197240000000
0!
0%
#197245000000
1!
1%
#197250000000
0!
0%
#197255000000
1!
1%
#197260000000
0!
0%
#197265000000
1!
1%
#197270000000
0!
0%
#197275000000
1!
1%
#197280000000
0!
0%
#197285000000
1!
1%
#197290000000
0!
0%
#197295000000
1!
1%
#197300000000
0!
0%
#197305000000
1!
1%
#197310000000
0!
0%
#197315000000
1!
1%
#197320000000
0!
0%
#197325000000
1!
1%
#197330000000
0!
0%
#197335000000
1!
1%
#197340000000
0!
0%
#197345000000
1!
1%
#197350000000
0!
0%
#197355000000
1!
1%
#197360000000
0!
0%
#197365000000
1!
1%
#197370000000
0!
0%
#197375000000
1!
1%
#197380000000
0!
0%
#197385000000
1!
1%
#197390000000
0!
0%
#197395000000
1!
1%
#197400000000
0!
0%
#197405000000
1!
1%
#197410000000
0!
0%
#197415000000
1!
1%
#197420000000
0!
0%
#197425000000
1!
1%
#197430000000
0!
0%
#197435000000
1!
1%
#197440000000
0!
0%
#197445000000
1!
1%
#197450000000
0!
0%
#197455000000
1!
1%
#197460000000
0!
0%
#197465000000
1!
1%
#197470000000
0!
0%
#197475000000
1!
1%
#197480000000
0!
0%
#197485000000
1!
1%
#197490000000
0!
0%
#197495000000
1!
1%
#197500000000
0!
0%
#197505000000
1!
1%
#197510000000
0!
0%
#197515000000
1!
1%
#197520000000
0!
0%
#197525000000
1!
1%
#197530000000
0!
0%
#197535000000
1!
1%
#197540000000
0!
0%
#197545000000
1!
1%
#197550000000
0!
0%
#197555000000
1!
1%
#197560000000
0!
0%
#197565000000
1!
1%
#197570000000
0!
0%
#197575000000
1!
1%
#197580000000
0!
0%
#197585000000
1!
1%
#197590000000
0!
0%
#197595000000
1!
1%
#197600000000
0!
0%
#197605000000
1!
1%
#197610000000
0!
0%
#197615000000
1!
1%
#197620000000
0!
0%
#197625000000
1!
1%
#197630000000
0!
0%
#197635000000
1!
1%
#197640000000
0!
0%
#197645000000
1!
1%
#197650000000
0!
0%
#197655000000
1!
1%
#197660000000
0!
0%
#197665000000
1!
1%
#197670000000
0!
0%
#197675000000
1!
1%
#197680000000
0!
0%
#197685000000
1!
1%
#197690000000
0!
0%
#197695000000
1!
1%
#197700000000
0!
0%
#197705000000
1!
1%
#197710000000
0!
0%
#197715000000
1!
1%
#197720000000
0!
0%
#197725000000
1!
1%
#197730000000
0!
0%
#197735000000
1!
1%
#197740000000
0!
0%
#197745000000
1!
1%
#197750000000
0!
0%
#197755000000
1!
1%
#197760000000
0!
0%
#197765000000
1!
1%
#197770000000
0!
0%
#197775000000
1!
1%
#197780000000
0!
0%
#197785000000
1!
1%
#197790000000
0!
0%
#197795000000
1!
1%
#197800000000
0!
0%
#197805000000
1!
1%
#197810000000
0!
0%
#197815000000
1!
1%
#197820000000
0!
0%
#197825000000
1!
1%
#197830000000
0!
0%
#197835000000
1!
1%
#197840000000
0!
0%
#197845000000
1!
1%
#197850000000
0!
0%
#197855000000
1!
1%
#197860000000
0!
0%
#197865000000
1!
1%
#197870000000
0!
0%
#197875000000
1!
1%
#197880000000
0!
0%
#197885000000
1!
1%
#197890000000
0!
0%
#197895000000
1!
1%
#197900000000
0!
0%
#197905000000
1!
1%
#197910000000
0!
0%
#197915000000
1!
1%
#197920000000
0!
0%
#197925000000
1!
1%
#197930000000
0!
0%
#197935000000
1!
1%
#197940000000
0!
0%
#197945000000
1!
1%
#197950000000
0!
0%
#197955000000
1!
1%
#197960000000
0!
0%
#197965000000
1!
1%
#197970000000
0!
0%
#197975000000
1!
1%
#197980000000
0!
0%
#197985000000
1!
1%
#197990000000
0!
0%
#197995000000
1!
1%
#198000000000
0!
0%
#198005000000
1!
1%
#198010000000
0!
0%
#198015000000
1!
1%
#198020000000
0!
0%
#198025000000
1!
1%
#198030000000
0!
0%
#198035000000
1!
1%
#198040000000
0!
0%
#198045000000
1!
1%
#198050000000
0!
0%
#198055000000
1!
1%
#198060000000
0!
0%
#198065000000
1!
1%
#198070000000
0!
0%
#198075000000
1!
1%
#198080000000
0!
0%
#198085000000
1!
1%
#198090000000
0!
0%
#198095000000
1!
1%
#198100000000
0!
0%
#198105000000
1!
1%
#198110000000
0!
0%
#198115000000
1!
1%
#198120000000
0!
0%
#198125000000
1!
1%
#198130000000
0!
0%
#198135000000
1!
1%
#198140000000
0!
0%
#198145000000
1!
1%
#198150000000
0!
0%
#198155000000
1!
1%
#198160000000
0!
0%
#198165000000
1!
1%
#198170000000
0!
0%
#198175000000
1!
1%
#198180000000
0!
0%
#198185000000
1!
1%
#198190000000
0!
0%
#198195000000
1!
1%
#198200000000
0!
0%
#198205000000
1!
1%
#198210000000
0!
0%
#198215000000
1!
1%
#198220000000
0!
0%
#198225000000
1!
1%
#198230000000
0!
0%
#198235000000
1!
1%
#198240000000
0!
0%
#198245000000
1!
1%
#198250000000
0!
0%
#198255000000
1!
1%
#198260000000
0!
0%
#198265000000
1!
1%
#198270000000
0!
0%
#198275000000
1!
1%
#198280000000
0!
0%
#198285000000
1!
1%
#198290000000
0!
0%
#198295000000
1!
1%
#198300000000
0!
0%
#198305000000
1!
1%
#198310000000
0!
0%
#198315000000
1!
1%
#198320000000
0!
0%
#198325000000
1!
1%
#198330000000
0!
0%
#198335000000
1!
1%
#198340000000
0!
0%
#198345000000
1!
1%
#198350000000
0!
0%
#198355000000
1!
1%
#198360000000
0!
0%
#198365000000
1!
1%
#198370000000
0!
0%
#198375000000
1!
1%
#198380000000
0!
0%
#198385000000
1!
1%
#198390000000
0!
0%
#198395000000
1!
1%
#198400000000
0!
0%
#198405000000
1!
1%
#198410000000
0!
0%
#198415000000
1!
1%
#198420000000
0!
0%
#198425000000
1!
1%
#198430000000
0!
0%
#198435000000
1!
1%
#198440000000
0!
0%
#198445000000
1!
1%
#198450000000
0!
0%
#198455000000
1!
1%
#198460000000
0!
0%
#198465000000
1!
1%
#198470000000
0!
0%
#198475000000
1!
1%
#198480000000
0!
0%
#198485000000
1!
1%
#198490000000
0!
0%
#198495000000
1!
1%
#198500000000
0!
0%
#198505000000
1!
1%
#198510000000
0!
0%
#198515000000
1!
1%
#198520000000
0!
0%
#198525000000
1!
1%
#198530000000
0!
0%
#198535000000
1!
1%
#198540000000
0!
0%
#198545000000
1!
1%
#198550000000
0!
0%
#198555000000
1!
1%
#198560000000
0!
0%
#198565000000
1!
1%
#198570000000
0!
0%
#198575000000
1!
1%
#198580000000
0!
0%
#198585000000
1!
1%
#198590000000
0!
0%
#198595000000
1!
1%
#198600000000
0!
0%
#198605000000
1!
1%
#198610000000
0!
0%
#198615000000
1!
1%
#198620000000
0!
0%
#198625000000
1!
1%
#198630000000
0!
0%
#198635000000
1!
1%
#198640000000
0!
0%
#198645000000
1!
1%
#198650000000
0!
0%
#198655000000
1!
1%
#198660000000
0!
0%
#198665000000
1!
1%
#198670000000
0!
0%
#198675000000
1!
1%
#198680000000
0!
0%
#198685000000
1!
1%
#198690000000
0!
0%
#198695000000
1!
1%
#198700000000
0!
0%
#198705000000
1!
1%
#198710000000
0!
0%
#198715000000
1!
1%
#198720000000
0!
0%
#198725000000
1!
1%
#198730000000
0!
0%
#198735000000
1!
1%
#198740000000
0!
0%
#198745000000
1!
1%
#198750000000
0!
0%
#198755000000
1!
1%
#198760000000
0!
0%
#198765000000
1!
1%
#198770000000
0!
0%
#198775000000
1!
1%
#198780000000
0!
0%
#198785000000
1!
1%
#198790000000
0!
0%
#198795000000
1!
1%
#198800000000
0!
0%
#198805000000
1!
1%
#198810000000
0!
0%
#198815000000
1!
1%
#198820000000
0!
0%
#198825000000
1!
1%
#198830000000
0!
0%
#198835000000
1!
1%
#198840000000
0!
0%
#198845000000
1!
1%
#198850000000
0!
0%
#198855000000
1!
1%
#198860000000
0!
0%
#198865000000
1!
1%
#198870000000
0!
0%
#198875000000
1!
1%
#198880000000
0!
0%
#198885000000
1!
1%
#198890000000
0!
0%
#198895000000
1!
1%
#198900000000
0!
0%
#198905000000
1!
1%
#198910000000
0!
0%
#198915000000
1!
1%
#198920000000
0!
0%
#198925000000
1!
1%
#198930000000
0!
0%
#198935000000
1!
1%
#198940000000
0!
0%
#198945000000
1!
1%
#198950000000
0!
0%
#198955000000
1!
1%
#198960000000
0!
0%
#198965000000
1!
1%
#198970000000
0!
0%
#198975000000
1!
1%
#198980000000
0!
0%
#198985000000
1!
1%
#198990000000
0!
0%
#198995000000
1!
1%
#199000000000
0!
0%
#199005000000
1!
1%
#199010000000
0!
0%
#199015000000
1!
1%
#199020000000
0!
0%
#199025000000
1!
1%
#199030000000
0!
0%
#199035000000
1!
1%
#199040000000
0!
0%
#199045000000
1!
1%
#199050000000
0!
0%
#199055000000
1!
1%
#199060000000
0!
0%
#199065000000
1!
1%
#199070000000
0!
0%
#199075000000
1!
1%
#199080000000
0!
0%
#199085000000
1!
1%
#199090000000
0!
0%
#199095000000
1!
1%
#199100000000
0!
0%
#199105000000
1!
1%
#199110000000
0!
0%
#199115000000
1!
1%
#199120000000
0!
0%
#199125000000
1!
1%
#199130000000
0!
0%
#199135000000
1!
1%
#199140000000
0!
0%
#199145000000
1!
1%
#199150000000
0!
0%
#199155000000
1!
1%
#199160000000
0!
0%
#199165000000
1!
1%
#199170000000
0!
0%
#199175000000
1!
1%
#199180000000
0!
0%
#199185000000
1!
1%
#199190000000
0!
0%
#199195000000
1!
1%
#199200000000
0!
0%
#199205000000
1!
1%
#199210000000
0!
0%
#199215000000
1!
1%
#199220000000
0!
0%
#199225000000
1!
1%
#199230000000
0!
0%
#199235000000
1!
1%
#199240000000
0!
0%
#199245000000
1!
1%
#199250000000
0!
0%
#199255000000
1!
1%
#199260000000
0!
0%
#199265000000
1!
1%
#199270000000
0!
0%
#199275000000
1!
1%
#199280000000
0!
0%
#199285000000
1!
1%
#199290000000
0!
0%
#199295000000
1!
1%
#199300000000
0!
0%
#199305000000
1!
1%
#199310000000
0!
0%
#199315000000
1!
1%
#199320000000
0!
0%
#199325000000
1!
1%
#199330000000
0!
0%
#199335000000
1!
1%
#199340000000
0!
0%
#199345000000
1!
1%
#199350000000
0!
0%
#199355000000
1!
1%
#199360000000
0!
0%
#199365000000
1!
1%
#199370000000
0!
0%
#199375000000
1!
1%
#199380000000
0!
0%
#199385000000
1!
1%
#199390000000
0!
0%
#199395000000
1!
1%
#199400000000
0!
0%
#199405000000
1!
1%
#199410000000
0!
0%
#199415000000
1!
1%
#199420000000
0!
0%
#199425000000
1!
1%
#199430000000
0!
0%
#199435000000
1!
1%
#199440000000
0!
0%
#199445000000
1!
1%
#199450000000
0!
0%
#199455000000
1!
1%
#199460000000
0!
0%
#199465000000
1!
1%
#199470000000
0!
0%
#199475000000
1!
1%
#199480000000
0!
0%
#199485000000
1!
1%
#199490000000
0!
0%
#199495000000
1!
1%
#199500000000
0!
0%
#199505000000
1!
1%
#199510000000
0!
0%
#199515000000
1!
1%
#199520000000
0!
0%
#199525000000
1!
1%
#199530000000
0!
0%
#199535000000
1!
1%
#199540000000
0!
0%
#199545000000
1!
1%
#199550000000
0!
0%
#199555000000
1!
1%
#199560000000
0!
0%
#199565000000
1!
1%
#199570000000
0!
0%
#199575000000
1!
1%
#199580000000
0!
0%
#199585000000
1!
1%
#199590000000
0!
0%
#199595000000
1!
1%
#199600000000
0!
0%
#199605000000
1!
1%
#199610000000
0!
0%
#199615000000
1!
1%
#199620000000
0!
0%
#199625000000
1!
1%
#199630000000
0!
0%
#199635000000
1!
1%
#199640000000
0!
0%
#199645000000
1!
1%
#199650000000
0!
0%
#199655000000
1!
1%
#199660000000
0!
0%
#199665000000
1!
1%
#199670000000
0!
0%
#199675000000
1!
1%
#199680000000
0!
0%
#199685000000
1!
1%
#199690000000
0!
0%
#199695000000
1!
1%
#199700000000
0!
0%
#199705000000
1!
1%
#199710000000
0!
0%
#199715000000
1!
1%
#199720000000
0!
0%
#199725000000
1!
1%
#199730000000
0!
0%
#199735000000
1!
1%
#199740000000
0!
0%
#199745000000
1!
1%
#199750000000
0!
0%
#199755000000
1!
1%
#199760000000
0!
0%
#199765000000
1!
1%
#199770000000
0!
0%
#199775000000
1!
1%
#199780000000
0!
0%
#199785000000
1!
1%
#199790000000
0!
0%
#199795000000
1!
1%
#199800000000
0!
0%
#199805000000
1!
1%
#199810000000
0!
0%
#199815000000
1!
1%
#199820000000
0!
0%
#199825000000
1!
1%
#199830000000
0!
0%
#199835000000
1!
1%
#199840000000
0!
0%
#199845000000
1!
1%
#199850000000
0!
0%
#199855000000
1!
1%
#199860000000
0!
0%
#199865000000
1!
1%
#199870000000
0!
0%
#199875000000
1!
1%
#199880000000
0!
0%
#199885000000
1!
1%
#199890000000
0!
0%
#199895000000
1!
1%
#199900000000
0!
0%
#199905000000
1!
1%
#199910000000
0!
0%
#199915000000
1!
1%
#199920000000
0!
0%
#199925000000
1!
1%
#199930000000
0!
0%
#199935000000
1!
1%
#199940000000
0!
0%
#199945000000
1!
1%
#199950000000
0!
0%
#199955000000
1!
1%
#199960000000
0!
0%
#199965000000
1!
1%
#199970000000
0!
0%
#199975000000
1!
1%
#199980000000
0!
0%
#199985000000
1!
1%
#199990000000
0!
0%
#199995000000
1!
1%
#200000000000
0!
0%
#200005000000
1!
1%
#200010000000
0!
0%
#200015000000
1!
1%
#200020000000
0!
0%
#200025000000
1!
1%
#200030000000
0!
0%
#200035000000
1!
1%
#200040000000
0!
0%
#200045000000
1!
1%
#200050000000
0!
0%
#200055000000
1!
1%
#200060000000
0!
0%
#200065000000
1!
1%
#200070000000
0!
0%
#200075000000
1!
1%
#200080000000
0!
0%
#200085000000
1!
1%
#200090000000
0!
0%
#200095000000
1!
1%
#200100000000
0!
0%
#200105000000
1!
1%
#200110000000
0!
0%
#200115000000
1!
1%
#200120000000
0!
0%
#200125000000
1!
1%
#200130000000
0!
0%
#200135000000
1!
1%
#200140000000
0!
0%
#200145000000
1!
1%
#200150000000
0!
0%
#200155000000
1!
1%
#200160000000
0!
0%
#200165000000
1!
1%
#200170000000
0!
0%
#200175000000
1!
1%
#200180000000
0!
0%
#200185000000
1!
1%
#200190000000
0!
0%
#200195000000
1!
1%
#200200000000
0!
0%
#200205000000
1!
1%
#200210000000
0!
0%
#200215000000
1!
1%
#200220000000
0!
0%
#200225000000
1!
1%
#200230000000
0!
0%
#200235000000
1!
1%
#200240000000
0!
0%
#200245000000
1!
1%
#200250000000
0!
0%
#200255000000
1!
1%
#200260000000
0!
0%
#200265000000
1!
1%
#200270000000
0!
0%
#200275000000
1!
1%
#200280000000
0!
0%
#200285000000
1!
1%
#200290000000
0!
0%
#200295000000
1!
1%
#200300000000
0!
0%
#200305000000
1!
1%
#200310000000
0!
0%
#200315000000
1!
1%
#200320000000
0!
0%
#200325000000
1!
1%
#200330000000
0!
0%
#200335000000
1!
1%
#200340000000
0!
0%
#200345000000
1!
1%
#200350000000
0!
0%
#200355000000
1!
1%
#200360000000
0!
0%
#200365000000
1!
1%
#200370000000
0!
0%
#200375000000
1!
1%
#200380000000
0!
0%
#200385000000
1!
1%
#200390000000
0!
0%
#200395000000
1!
1%
#200400000000
0!
0%
#200405000000
1!
1%
#200410000000
0!
0%
#200415000000
1!
1%
#200420000000
0!
0%
#200425000000
1!
1%
#200430000000
0!
0%
#200435000000
1!
1%
#200440000000
0!
0%
#200445000000
1!
1%
#200450000000
0!
0%
#200455000000
1!
1%
#200460000000
0!
0%
#200465000000
1!
1%
#200470000000
0!
0%
#200475000000
1!
1%
#200480000000
0!
0%
#200485000000
1!
1%
#200490000000
0!
0%
#200495000000
1!
1%
#200500000000
0!
0%
#200505000000
1!
1%
#200510000000
0!
0%
#200515000000
1!
1%
#200520000000
0!
0%
#200525000000
1!
1%
#200530000000
0!
0%
#200535000000
1!
1%
#200540000000
0!
0%
#200545000000
1!
1%
#200550000000
0!
0%
#200555000000
1!
1%
#200560000000
0!
0%
#200565000000
1!
1%
#200570000000
0!
0%
#200575000000
1!
1%
#200580000000
0!
0%
#200585000000
1!
1%
#200590000000
0!
0%
#200595000000
1!
1%
#200600000000
0!
0%
#200605000000
1!
1%
#200610000000
0!
0%
#200615000000
1!
1%
#200620000000
0!
0%
#200625000000
1!
1%
#200630000000
0!
0%
#200635000000
1!
1%
#200640000000
0!
0%
#200645000000
1!
1%
#200650000000
0!
0%
#200655000000
1!
1%
#200660000000
0!
0%
#200665000000
1!
1%
#200670000000
0!
0%
#200675000000
1!
1%
#200680000000
0!
0%
#200685000000
1!
1%
#200690000000
0!
0%
#200695000000
1!
1%
#200700000000
0!
0%
#200705000000
1!
1%
#200710000000
0!
0%
#200715000000
1!
1%
#200720000000
0!
0%
#200725000000
1!
1%
#200730000000
0!
0%
#200735000000
1!
1%
#200740000000
0!
0%
#200745000000
1!
1%
#200750000000
0!
0%
#200755000000
1!
1%
#200760000000
0!
0%
#200765000000
1!
1%
#200770000000
0!
0%
#200775000000
1!
1%
#200780000000
0!
0%
#200785000000
1!
1%
#200790000000
0!
0%
#200795000000
1!
1%
#200800000000
0!
0%
#200805000000
1!
1%
#200810000000
0!
0%
#200815000000
1!
1%
#200820000000
0!
0%
#200825000000
1!
1%
#200830000000
0!
0%
#200835000000
1!
1%
#200840000000
0!
0%
#200845000000
1!
1%
#200850000000
0!
0%
#200855000000
1!
1%
#200860000000
0!
0%
#200865000000
1!
1%
#200870000000
0!
0%
#200875000000
1!
1%
#200880000000
0!
0%
#200885000000
1!
1%
#200890000000
0!
0%
#200895000000
1!
1%
#200900000000
0!
0%
#200905000000
1!
1%
#200910000000
0!
0%
#200915000000
1!
1%
#200920000000
0!
0%
#200925000000
1!
1%
#200930000000
0!
0%
#200935000000
1!
1%
#200940000000
0!
0%
#200945000000
1!
1%
#200950000000
0!
0%
#200955000000
1!
1%
#200960000000
0!
0%
#200965000000
1!
1%
#200970000000
0!
0%
#200975000000
1!
1%
#200980000000
0!
0%
#200985000000
1!
1%
#200990000000
0!
0%
#200995000000
1!
1%
#201000000000
0!
0%
#201005000000
1!
1%
#201010000000
0!
0%
#201015000000
1!
1%
#201020000000
0!
0%
#201025000000
1!
1%
#201030000000
0!
0%
#201035000000
1!
1%
#201040000000
0!
0%
#201045000000
1!
1%
#201050000000
0!
0%
#201055000000
1!
1%
#201060000000
0!
0%
#201065000000
1!
1%
#201070000000
0!
0%
#201075000000
1!
1%
#201080000000
0!
0%
#201085000000
1!
1%
#201090000000
0!
0%
#201095000000
1!
1%
#201100000000
0!
0%
#201105000000
1!
1%
#201110000000
0!
0%
#201115000000
1!
1%
#201120000000
0!
0%
#201125000000
1!
1%
#201130000000
0!
0%
#201135000000
1!
1%
#201140000000
0!
0%
#201145000000
1!
1%
#201150000000
0!
0%
#201155000000
1!
1%
#201160000000
0!
0%
#201165000000
1!
1%
#201170000000
0!
0%
#201175000000
1!
1%
#201180000000
0!
0%
#201185000000
1!
1%
#201190000000
0!
0%
#201195000000
1!
1%
#201200000000
0!
0%
#201205000000
1!
1%
#201210000000
0!
0%
#201215000000
1!
1%
#201220000000
0!
0%
#201225000000
1!
1%
#201230000000
0!
0%
#201235000000
1!
1%
#201240000000
0!
0%
#201245000000
1!
1%
#201250000000
0!
0%
#201255000000
1!
1%
#201260000000
0!
0%
#201265000000
1!
1%
#201270000000
0!
0%
#201275000000
1!
1%
#201280000000
0!
0%
#201285000000
1!
1%
#201290000000
0!
0%
#201295000000
1!
1%
#201300000000
0!
0%
#201305000000
1!
1%
#201310000000
0!
0%
#201315000000
1!
1%
#201320000000
0!
0%
#201325000000
1!
1%
#201330000000
0!
0%
#201335000000
1!
1%
#201340000000
0!
0%
#201345000000
1!
1%
#201350000000
0!
0%
#201355000000
1!
1%
#201360000000
0!
0%
#201365000000
1!
1%
#201370000000
0!
0%
#201375000000
1!
1%
#201380000000
0!
0%
#201385000000
1!
1%
#201390000000
0!
0%
#201395000000
1!
1%
#201400000000
0!
0%
#201405000000
1!
1%
#201410000000
0!
0%
#201415000000
1!
1%
#201420000000
0!
0%
#201425000000
1!
1%
#201430000000
0!
0%
#201435000000
1!
1%
#201440000000
0!
0%
#201445000000
1!
1%
#201450000000
0!
0%
#201455000000
1!
1%
#201460000000
0!
0%
#201465000000
1!
1%
#201470000000
0!
0%
#201475000000
1!
1%
#201480000000
0!
0%
#201485000000
1!
1%
#201490000000
0!
0%
#201495000000
1!
1%
#201500000000
0!
0%
#201505000000
1!
1%
#201510000000
0!
0%
#201515000000
1!
1%
#201520000000
0!
0%
#201525000000
1!
1%
#201530000000
0!
0%
#201535000000
1!
1%
#201540000000
0!
0%
#201545000000
1!
1%
#201550000000
0!
0%
#201555000000
1!
1%
#201560000000
0!
0%
#201565000000
1!
1%
#201570000000
0!
0%
#201575000000
1!
1%
#201580000000
0!
0%
#201585000000
1!
1%
#201590000000
0!
0%
#201595000000
1!
1%
#201600000000
0!
0%
#201605000000
1!
1%
#201610000000
0!
0%
#201615000000
1!
1%
#201620000000
0!
0%
#201625000000
1!
1%
#201630000000
0!
0%
#201635000000
1!
1%
#201640000000
0!
0%
#201645000000
1!
1%
#201650000000
0!
0%
#201655000000
1!
1%
#201660000000
0!
0%
#201665000000
1!
1%
#201670000000
0!
0%
#201675000000
1!
1%
#201680000000
0!
0%
#201685000000
1!
1%
#201690000000
0!
0%
#201695000000
1!
1%
#201700000000
0!
0%
#201705000000
1!
1%
#201710000000
0!
0%
#201715000000
1!
1%
#201720000000
0!
0%
#201725000000
1!
1%
#201730000000
0!
0%
#201735000000
1!
1%
#201740000000
0!
0%
#201745000000
1!
1%
#201750000000
0!
0%
#201755000000
1!
1%
#201760000000
0!
0%
#201765000000
1!
1%
#201770000000
0!
0%
#201775000000
1!
1%
#201780000000
0!
0%
#201785000000
1!
1%
#201790000000
0!
0%
#201795000000
1!
1%
#201800000000
0!
0%
#201805000000
1!
1%
#201810000000
0!
0%
#201815000000
1!
1%
#201820000000
0!
0%
#201825000000
1!
1%
#201830000000
0!
0%
#201835000000
1!
1%
#201840000000
0!
0%
#201845000000
1!
1%
#201850000000
0!
0%
#201855000000
1!
1%
#201860000000
0!
0%
#201865000000
1!
1%
#201870000000
0!
0%
#201875000000
1!
1%
#201880000000
0!
0%
#201885000000
1!
1%
#201890000000
0!
0%
#201895000000
1!
1%
#201900000000
0!
0%
#201905000000
1!
1%
#201910000000
0!
0%
#201915000000
1!
1%
#201920000000
0!
0%
#201925000000
1!
1%
#201930000000
0!
0%
#201935000000
1!
1%
#201940000000
0!
0%
#201945000000
1!
1%
#201950000000
0!
0%
#201955000000
1!
1%
#201960000000
0!
0%
#201965000000
1!
1%
#201970000000
0!
0%
#201975000000
1!
1%
#201980000000
0!
0%
#201985000000
1!
1%
#201990000000
0!
0%
#201995000000
1!
1%
#202000000000
0!
0%
#202005000000
1!
1%
#202010000000
0!
0%
#202015000000
1!
1%
#202020000000
0!
0%
#202025000000
1!
1%
#202030000000
0!
0%
#202035000000
1!
1%
#202040000000
0!
0%
#202045000000
1!
1%
#202050000000
0!
0%
#202055000000
1!
1%
#202060000000
0!
0%
#202065000000
1!
1%
#202070000000
0!
0%
#202075000000
1!
1%
#202080000000
0!
0%
#202085000000
1!
1%
#202090000000
0!
0%
#202095000000
1!
1%
#202100000000
0!
0%
#202105000000
1!
1%
#202110000000
0!
0%
#202115000000
1!
1%
#202120000000
0!
0%
#202125000000
1!
1%
#202130000000
0!
0%
#202135000000
1!
1%
#202140000000
0!
0%
#202145000000
1!
1%
#202150000000
0!
0%
#202155000000
1!
1%
#202160000000
0!
0%
#202165000000
1!
1%
#202170000000
0!
0%
#202175000000
1!
1%
#202180000000
0!
0%
#202185000000
1!
1%
#202190000000
0!
0%
#202195000000
1!
1%
#202200000000
0!
0%
#202205000000
1!
1%
#202210000000
0!
0%
#202215000000
1!
1%
#202220000000
0!
0%
#202225000000
1!
1%
#202230000000
0!
0%
#202235000000
1!
1%
#202240000000
0!
0%
#202245000000
1!
1%
#202250000000
0!
0%
#202255000000
1!
1%
#202260000000
0!
0%
#202265000000
1!
1%
#202270000000
0!
0%
#202275000000
1!
1%
#202280000000
0!
0%
#202285000000
1!
1%
#202290000000
0!
0%
#202295000000
1!
1%
#202300000000
0!
0%
#202305000000
1!
1%
#202310000000
0!
0%
#202315000000
1!
1%
#202320000000
0!
0%
#202325000000
1!
1%
#202330000000
0!
0%
#202335000000
1!
1%
#202340000000
0!
0%
#202345000000
1!
1%
#202350000000
0!
0%
#202355000000
1!
1%
#202360000000
0!
0%
#202365000000
1!
1%
#202370000000
0!
0%
#202375000000
1!
1%
#202380000000
0!
0%
#202385000000
1!
1%
#202390000000
0!
0%
#202395000000
1!
1%
#202400000000
0!
0%
#202405000000
1!
1%
#202410000000
0!
0%
#202415000000
1!
1%
#202420000000
0!
0%
#202425000000
1!
1%
#202430000000
0!
0%
#202435000000
1!
1%
#202440000000
0!
0%
#202445000000
1!
1%
#202450000000
0!
0%
#202455000000
1!
1%
#202460000000
0!
0%
#202465000000
1!
1%
#202470000000
0!
0%
#202475000000
1!
1%
#202480000000
0!
0%
#202485000000
1!
1%
#202490000000
0!
0%
#202495000000
1!
1%
#202500000000
0!
0%
#202505000000
1!
1%
#202510000000
0!
0%
#202515000000
1!
1%
#202520000000
0!
0%
#202525000000
1!
1%
#202530000000
0!
0%
#202535000000
1!
1%
#202540000000
0!
0%
#202545000000
1!
1%
#202550000000
0!
0%
#202555000000
1!
1%
#202560000000
0!
0%
#202565000000
1!
1%
#202570000000
0!
0%
#202575000000
1!
1%
#202580000000
0!
0%
#202585000000
1!
1%
#202590000000
0!
0%
#202595000000
1!
1%
#202600000000
0!
0%
#202605000000
1!
1%
#202610000000
0!
0%
#202615000000
1!
1%
#202620000000
0!
0%
#202625000000
1!
1%
#202630000000
0!
0%
#202635000000
1!
1%
#202640000000
0!
0%
#202645000000
1!
1%
#202650000000
0!
0%
#202655000000
1!
1%
#202660000000
0!
0%
#202665000000
1!
1%
#202670000000
0!
0%
#202675000000
1!
1%
#202680000000
0!
0%
#202685000000
1!
1%
#202690000000
0!
0%
#202695000000
1!
1%
#202700000000
0!
0%
#202705000000
1!
1%
#202710000000
0!
0%
#202715000000
1!
1%
#202720000000
0!
0%
#202725000000
1!
1%
#202730000000
0!
0%
#202735000000
1!
1%
#202740000000
0!
0%
#202745000000
1!
1%
#202750000000
0!
0%
#202755000000
1!
1%
#202760000000
0!
0%
#202765000000
1!
1%
#202770000000
0!
0%
#202775000000
1!
1%
#202780000000
0!
0%
#202785000000
1!
1%
#202790000000
0!
0%
#202795000000
1!
1%
#202800000000
0!
0%
#202805000000
1!
1%
#202810000000
0!
0%
#202815000000
1!
1%
#202820000000
0!
0%
#202825000000
1!
1%
#202830000000
0!
0%
#202835000000
1!
1%
#202840000000
0!
0%
#202845000000
1!
1%
#202850000000
0!
0%
#202855000000
1!
1%
#202860000000
0!
0%
#202865000000
1!
1%
#202870000000
0!
0%
#202875000000
1!
1%
#202880000000
0!
0%
#202885000000
1!
1%
#202890000000
0!
0%
#202895000000
1!
1%
#202900000000
0!
0%
#202905000000
1!
1%
#202910000000
0!
0%
#202915000000
1!
1%
#202920000000
0!
0%
#202925000000
1!
1%
#202930000000
0!
0%
#202935000000
1!
1%
#202940000000
0!
0%
#202945000000
1!
1%
#202950000000
0!
0%
#202955000000
1!
1%
#202960000000
0!
0%
#202965000000
1!
1%
#202970000000
0!
0%
#202975000000
1!
1%
#202980000000
0!
0%
#202985000000
1!
1%
#202990000000
0!
0%
#202995000000
1!
1%
#203000000000
0!
0%
#203005000000
1!
1%
#203010000000
0!
0%
#203015000000
1!
1%
#203020000000
0!
0%
#203025000000
1!
1%
#203030000000
0!
0%
#203035000000
1!
1%
#203040000000
0!
0%
#203045000000
1!
1%
#203050000000
0!
0%
#203055000000
1!
1%
#203060000000
0!
0%
#203065000000
1!
1%
#203070000000
0!
0%
#203075000000
1!
1%
#203080000000
0!
0%
#203085000000
1!
1%
#203090000000
0!
0%
#203095000000
1!
1%
#203100000000
0!
0%
#203105000000
1!
1%
#203110000000
0!
0%
#203115000000
1!
1%
#203120000000
0!
0%
#203125000000
1!
1%
#203130000000
0!
0%
#203135000000
1!
1%
#203140000000
0!
0%
#203145000000
1!
1%
#203150000000
0!
0%
#203155000000
1!
1%
#203160000000
0!
0%
#203165000000
1!
1%
#203170000000
0!
0%
#203175000000
1!
1%
#203180000000
0!
0%
#203185000000
1!
1%
#203190000000
0!
0%
#203195000000
1!
1%
#203200000000
0!
0%
#203205000000
1!
1%
#203210000000
0!
0%
#203215000000
1!
1%
#203220000000
0!
0%
#203225000000
1!
1%
#203230000000
0!
0%
#203235000000
1!
1%
#203240000000
0!
0%
#203245000000
1!
1%
#203250000000
0!
0%
#203255000000
1!
1%
#203260000000
0!
0%
#203265000000
1!
1%
#203270000000
0!
0%
#203275000000
1!
1%
#203280000000
0!
0%
#203285000000
1!
1%
#203290000000
0!
0%
#203295000000
1!
1%
#203300000000
0!
0%
#203305000000
1!
1%
#203310000000
0!
0%
#203315000000
1!
1%
#203320000000
0!
0%
#203325000000
1!
1%
#203330000000
0!
0%
#203335000000
1!
1%
#203340000000
0!
0%
#203345000000
1!
1%
#203350000000
0!
0%
#203355000000
1!
1%
#203360000000
0!
0%
#203365000000
1!
1%
#203370000000
0!
0%
#203375000000
1!
1%
#203380000000
0!
0%
#203385000000
1!
1%
#203390000000
0!
0%
#203395000000
1!
1%
#203400000000
0!
0%
#203405000000
1!
1%
#203410000000
0!
0%
#203415000000
1!
1%
#203420000000
0!
0%
#203425000000
1!
1%
#203430000000
0!
0%
#203435000000
1!
1%
#203440000000
0!
0%
#203445000000
1!
1%
#203450000000
0!
0%
#203455000000
1!
1%
#203460000000
0!
0%
#203465000000
1!
1%
#203470000000
0!
0%
#203475000000
1!
1%
#203480000000
0!
0%
#203485000000
1!
1%
#203490000000
0!
0%
#203495000000
1!
1%
#203500000000
0!
0%
#203505000000
1!
1%
#203510000000
0!
0%
#203515000000
1!
1%
#203520000000
0!
0%
#203525000000
1!
1%
#203530000000
0!
0%
#203535000000
1!
1%
#203540000000
0!
0%
#203545000000
1!
1%
#203550000000
0!
0%
#203555000000
1!
1%
#203560000000
0!
0%
#203565000000
1!
1%
#203570000000
0!
0%
#203575000000
1!
1%
#203580000000
0!
0%
#203585000000
1!
1%
#203590000000
0!
0%
#203595000000
1!
1%
#203600000000
0!
0%
#203605000000
1!
1%
#203610000000
0!
0%
#203615000000
1!
1%
#203620000000
0!
0%
#203625000000
1!
1%
#203630000000
0!
0%
#203635000000
1!
1%
#203640000000
0!
0%
#203645000000
1!
1%
#203650000000
0!
0%
#203655000000
1!
1%
#203660000000
0!
0%
#203665000000
1!
1%
#203670000000
0!
0%
#203675000000
1!
1%
#203680000000
0!
0%
#203685000000
1!
1%
#203690000000
0!
0%
#203695000000
1!
1%
#203700000000
0!
0%
#203705000000
1!
1%
#203710000000
0!
0%
#203715000000
1!
1%
#203720000000
0!
0%
#203725000000
1!
1%
#203730000000
0!
0%
#203735000000
1!
1%
#203740000000
0!
0%
#203745000000
1!
1%
#203750000000
0!
0%
#203755000000
1!
1%
#203760000000
0!
0%
#203765000000
1!
1%
#203770000000
0!
0%
#203775000000
1!
1%
#203780000000
0!
0%
#203785000000
1!
1%
#203790000000
0!
0%
#203795000000
1!
1%
#203800000000
0!
0%
#203805000000
1!
1%
#203810000000
0!
0%
#203815000000
1!
1%
#203820000000
0!
0%
#203825000000
1!
1%
#203830000000
0!
0%
#203835000000
1!
1%
#203840000000
0!
0%
#203845000000
1!
1%
#203850000000
0!
0%
#203855000000
1!
1%
#203860000000
0!
0%
#203865000000
1!
1%
#203870000000
0!
0%
#203875000000
1!
1%
#203880000000
0!
0%
#203885000000
1!
1%
#203890000000
0!
0%
#203895000000
1!
1%
#203900000000
0!
0%
#203905000000
1!
1%
#203910000000
0!
0%
#203915000000
1!
1%
#203920000000
0!
0%
#203925000000
1!
1%
#203930000000
0!
0%
#203935000000
1!
1%
#203940000000
0!
0%
#203945000000
1!
1%
#203950000000
0!
0%
#203955000000
1!
1%
#203960000000
0!
0%
#203965000000
1!
1%
#203970000000
0!
0%
#203975000000
1!
1%
#203980000000
0!
0%
#203985000000
1!
1%
#203990000000
0!
0%
#203995000000
1!
1%
#204000000000
0!
0%
#204005000000
1!
1%
#204010000000
0!
0%
#204015000000
1!
1%
#204020000000
0!
0%
#204025000000
1!
1%
#204030000000
0!
0%
#204035000000
1!
1%
#204040000000
0!
0%
#204045000000
1!
1%
#204050000000
0!
0%
#204055000000
1!
1%
#204060000000
0!
0%
#204065000000
1!
1%
#204070000000
0!
0%
#204075000000
1!
1%
#204080000000
0!
0%
#204085000000
1!
1%
#204090000000
0!
0%
#204095000000
1!
1%
#204100000000
0!
0%
#204105000000
1!
1%
#204110000000
0!
0%
#204115000000
1!
1%
#204120000000
0!
0%
#204125000000
1!
1%
#204130000000
0!
0%
#204135000000
1!
1%
#204140000000
0!
0%
#204145000000
1!
1%
#204150000000
0!
0%
#204155000000
1!
1%
#204160000000
0!
0%
#204165000000
1!
1%
#204170000000
0!
0%
#204175000000
1!
1%
#204180000000
0!
0%
#204185000000
1!
1%
#204190000000
0!
0%
#204195000000
1!
1%
#204200000000
0!
0%
#204205000000
1!
1%
#204210000000
0!
0%
#204215000000
1!
1%
#204220000000
0!
0%
#204225000000
1!
1%
#204230000000
0!
0%
#204235000000
1!
1%
#204240000000
0!
0%
#204245000000
1!
1%
#204250000000
0!
0%
#204255000000
1!
1%
#204260000000
0!
0%
#204265000000
1!
1%
#204270000000
0!
0%
#204275000000
1!
1%
#204280000000
0!
0%
#204285000000
1!
1%
#204290000000
0!
0%
#204295000000
1!
1%
#204300000000
0!
0%
#204305000000
1!
1%
#204310000000
0!
0%
#204315000000
1!
1%
#204320000000
0!
0%
#204325000000
1!
1%
#204330000000
0!
0%
#204335000000
1!
1%
#204340000000
0!
0%
#204345000000
1!
1%
#204350000000
0!
0%
#204355000000
1!
1%
#204360000000
0!
0%
#204365000000
1!
1%
#204370000000
0!
0%
#204375000000
1!
1%
#204380000000
0!
0%
#204385000000
1!
1%
#204390000000
0!
0%
#204395000000
1!
1%
#204400000000
0!
0%
#204405000000
1!
1%
#204410000000
0!
0%
#204415000000
1!
1%
#204420000000
0!
0%
#204425000000
1!
1%
#204430000000
0!
0%
#204435000000
1!
1%
#204440000000
0!
0%
#204445000000
1!
1%
#204450000000
0!
0%
#204455000000
1!
1%
#204460000000
0!
0%
#204465000000
1!
1%
#204470000000
0!
0%
#204475000000
1!
1%
#204480000000
0!
0%
#204485000000
1!
1%
#204490000000
0!
0%
#204495000000
1!
1%
#204500000000
0!
0%
#204505000000
1!
1%
#204510000000
0!
0%
#204515000000
1!
1%
#204520000000
0!
0%
#204525000000
1!
1%
#204530000000
0!
0%
#204535000000
1!
1%
#204540000000
0!
0%
#204545000000
1!
1%
#204550000000
0!
0%
#204555000000
1!
1%
#204560000000
0!
0%
#204565000000
1!
1%
#204570000000
0!
0%
#204575000000
1!
1%
#204580000000
0!
0%
#204585000000
1!
1%
#204590000000
0!
0%
#204595000000
1!
1%
#204600000000
0!
0%
#204605000000
1!
1%
#204610000000
0!
0%
#204615000000
1!
1%
#204620000000
0!
0%
#204625000000
1!
1%
#204630000000
0!
0%
#204635000000
1!
1%
#204640000000
0!
0%
#204645000000
1!
1%
#204650000000
0!
0%
#204655000000
1!
1%
#204660000000
0!
0%
#204665000000
1!
1%
#204670000000
0!
0%
#204675000000
1!
1%
#204680000000
0!
0%
#204685000000
1!
1%
#204690000000
0!
0%
#204695000000
1!
1%
#204700000000
0!
0%
#204705000000
1!
1%
#204710000000
0!
0%
#204715000000
1!
1%
#204720000000
0!
0%
#204725000000
1!
1%
#204730000000
0!
0%
#204735000000
1!
1%
#204740000000
0!
0%
#204745000000
1!
1%
#204750000000
0!
0%
#204755000000
1!
1%
#204760000000
0!
0%
#204765000000
1!
1%
#204770000000
0!
0%
#204775000000
1!
1%
#204780000000
0!
0%
#204785000000
1!
1%
#204790000000
0!
0%
#204795000000
1!
1%
#204800000000
0!
0%
#204805000000
1!
1%
#204810000000
0!
0%
#204815000000
1!
1%
#204820000000
0!
0%
#204825000000
1!
1%
#204830000000
0!
0%
#204835000000
1!
1%
#204840000000
0!
0%
#204845000000
1!
1%
#204850000000
0!
0%
#204855000000
1!
1%
#204860000000
0!
0%
#204865000000
1!
1%
#204870000000
0!
0%
#204875000000
1!
1%
#204880000000
0!
0%
#204885000000
1!
1%
#204890000000
0!
0%
#204895000000
1!
1%
#204900000000
0!
0%
#204905000000
1!
1%
#204910000000
0!
0%
#204915000000
1!
1%
#204920000000
0!
0%
#204925000000
1!
1%
#204930000000
0!
0%
#204935000000
1!
1%
#204940000000
0!
0%
#204945000000
1!
1%
#204950000000
0!
0%
#204955000000
1!
1%
#204960000000
0!
0%
#204965000000
1!
1%
#204970000000
0!
0%
#204975000000
1!
1%
#204980000000
0!
0%
#204985000000
1!
1%
#204990000000
0!
0%
#204995000000
1!
1%
#205000000000
0!
0%
#205005000000
1!
1%
#205010000000
0!
0%
#205015000000
1!
1%
#205020000000
0!
0%
#205025000000
1!
1%
#205030000000
0!
0%
#205035000000
1!
1%
#205040000000
0!
0%
#205045000000
1!
1%
#205050000000
0!
0%
#205055000000
1!
1%
#205060000000
0!
0%
#205065000000
1!
1%
#205070000000
0!
0%
#205075000000
1!
1%
#205080000000
0!
0%
#205085000000
1!
1%
#205090000000
0!
0%
#205095000000
1!
1%
#205100000000
0!
0%
#205105000000
1!
1%
#205110000000
0!
0%
#205115000000
1!
1%
#205120000000
0!
0%
#205125000000
1!
1%
#205130000000
0!
0%
#205135000000
1!
1%
#205140000000
0!
0%
#205145000000
1!
1%
#205150000000
0!
0%
#205155000000
1!
1%
#205160000000
0!
0%
#205165000000
1!
1%
#205170000000
0!
0%
#205175000000
1!
1%
#205180000000
0!
0%
#205185000000
1!
1%
#205190000000
0!
0%
#205195000000
1!
1%
#205200000000
0!
0%
#205205000000
1!
1%
#205210000000
0!
0%
#205215000000
1!
1%
#205220000000
0!
0%
#205225000000
1!
1%
#205230000000
0!
0%
#205235000000
1!
1%
#205240000000
0!
0%
#205245000000
1!
1%
#205250000000
0!
0%
#205255000000
1!
1%
#205260000000
0!
0%
#205265000000
1!
1%
#205270000000
0!
0%
#205275000000
1!
1%
#205280000000
0!
0%
#205285000000
1!
1%
#205290000000
0!
0%
#205295000000
1!
1%
#205300000000
0!
0%
#205305000000
1!
1%
#205310000000
0!
0%
#205315000000
1!
1%
#205320000000
0!
0%
#205325000000
1!
1%
#205330000000
0!
0%
#205335000000
1!
1%
#205340000000
0!
0%
#205345000000
1!
1%
#205350000000
0!
0%
#205355000000
1!
1%
#205360000000
0!
0%
#205365000000
1!
1%
#205370000000
0!
0%
#205375000000
1!
1%
#205380000000
0!
0%
#205385000000
1!
1%
#205390000000
0!
0%
#205395000000
1!
1%
#205400000000
0!
0%
#205405000000
1!
1%
#205410000000
0!
0%
#205415000000
1!
1%
#205420000000
0!
0%
#205425000000
1!
1%
#205430000000
0!
0%
#205435000000
1!
1%
#205440000000
0!
0%
#205445000000
1!
1%
#205450000000
0!
0%
#205455000000
1!
1%
#205460000000
0!
0%
#205465000000
1!
1%
#205470000000
0!
0%
#205475000000
1!
1%
#205480000000
0!
0%
#205485000000
1!
1%
#205490000000
0!
0%
#205495000000
1!
1%
#205500000000
0!
0%
#205505000000
1!
1%
#205510000000
0!
0%
#205515000000
1!
1%
#205520000000
0!
0%
#205525000000
1!
1%
#205530000000
0!
0%
#205535000000
1!
1%
#205540000000
0!
0%
#205545000000
1!
1%
#205550000000
0!
0%
#205555000000
1!
1%
#205560000000
0!
0%
#205565000000
1!
1%
#205570000000
0!
0%
#205575000000
1!
1%
#205580000000
0!
0%
#205585000000
1!
1%
#205590000000
0!
0%
#205595000000
1!
1%
#205600000000
0!
0%
#205605000000
1!
1%
#205610000000
0!
0%
#205615000000
1!
1%
#205620000000
0!
0%
#205625000000
1!
1%
#205630000000
0!
0%
#205635000000
1!
1%
#205640000000
0!
0%
#205645000000
1!
1%
#205650000000
0!
0%
#205655000000
1!
1%
#205660000000
0!
0%
#205665000000
1!
1%
#205670000000
0!
0%
#205675000000
1!
1%
#205680000000
0!
0%
#205685000000
1!
1%
#205690000000
0!
0%
#205695000000
1!
1%
#205700000000
0!
0%
#205705000000
1!
1%
#205710000000
0!
0%
#205715000000
1!
1%
#205720000000
0!
0%
#205725000000
1!
1%
#205730000000
0!
0%
#205735000000
1!
1%
#205740000000
0!
0%
#205745000000
1!
1%
#205750000000
0!
0%
#205755000000
1!
1%
#205760000000
0!
0%
#205765000000
1!
1%
#205770000000
0!
0%
#205775000000
1!
1%
#205780000000
0!
0%
#205785000000
1!
1%
#205790000000
0!
0%
#205795000000
1!
1%
#205800000000
0!
0%
#205805000000
1!
1%
#205810000000
0!
0%
#205815000000
1!
1%
#205820000000
0!
0%
#205825000000
1!
1%
#205830000000
0!
0%
#205835000000
1!
1%
#205840000000
0!
0%
#205845000000
1!
1%
#205850000000
0!
0%
#205855000000
1!
1%
#205860000000
0!
0%
#205865000000
1!
1%
#205870000000
0!
0%
#205875000000
1!
1%
#205880000000
0!
0%
#205885000000
1!
1%
#205890000000
0!
0%
#205895000000
1!
1%
#205900000000
0!
0%
#205905000000
1!
1%
#205910000000
0!
0%
#205915000000
1!
1%
#205920000000
0!
0%
#205925000000
1!
1%
#205930000000
0!
0%
#205935000000
1!
1%
#205940000000
0!
0%
#205945000000
1!
1%
#205950000000
0!
0%
#205955000000
1!
1%
#205960000000
0!
0%
#205965000000
1!
1%
#205970000000
0!
0%
#205975000000
1!
1%
#205980000000
0!
0%
#205985000000
1!
1%
#205990000000
0!
0%
#205995000000
1!
1%
#206000000000
0!
0%
#206005000000
1!
1%
#206010000000
0!
0%
#206015000000
1!
1%
#206020000000
0!
0%
#206025000000
1!
1%
#206030000000
0!
0%
#206035000000
1!
1%
#206040000000
0!
0%
#206045000000
1!
1%
#206050000000
0!
0%
#206055000000
1!
1%
#206060000000
0!
0%
#206065000000
1!
1%
#206070000000
0!
0%
#206075000000
1!
1%
#206080000000
0!
0%
#206085000000
1!
1%
#206090000000
0!
0%
#206095000000
1!
1%
#206100000000
0!
0%
#206105000000
1!
1%
#206110000000
0!
0%
#206115000000
1!
1%
#206120000000
0!
0%
#206125000000
1!
1%
#206130000000
0!
0%
#206135000000
1!
1%
#206140000000
0!
0%
#206145000000
1!
1%
#206150000000
0!
0%
#206155000000
1!
1%
#206160000000
0!
0%
#206165000000
1!
1%
#206170000000
0!
0%
#206175000000
1!
1%
#206180000000
0!
0%
#206185000000
1!
1%
#206190000000
0!
0%
#206195000000
1!
1%
#206200000000
0!
0%
#206205000000
1!
1%
#206210000000
0!
0%
#206215000000
1!
1%
#206220000000
0!
0%
#206225000000
1!
1%
#206230000000
0!
0%
#206235000000
1!
1%
#206240000000
0!
0%
#206245000000
1!
1%
#206250000000
0!
0%
#206255000000
1!
1%
#206260000000
0!
0%
#206265000000
1!
1%
#206270000000
0!
0%
#206275000000
1!
1%
#206280000000
0!
0%
#206285000000
1!
1%
#206290000000
0!
0%
#206295000000
1!
1%
#206300000000
0!
0%
#206305000000
1!
1%
#206310000000
0!
0%
#206315000000
1!
1%
#206320000000
0!
0%
#206325000000
1!
1%
#206330000000
0!
0%
#206335000000
1!
1%
#206340000000
0!
0%
#206345000000
1!
1%
#206350000000
0!
0%
#206355000000
1!
1%
#206360000000
0!
0%
#206365000000
1!
1%
#206370000000
0!
0%
#206375000000
1!
1%
#206380000000
0!
0%
#206385000000
1!
1%
#206390000000
0!
0%
#206395000000
1!
1%
#206400000000
0!
0%
#206405000000
1!
1%
#206410000000
0!
0%
#206415000000
1!
1%
#206420000000
0!
0%
#206425000000
1!
1%
#206430000000
0!
0%
#206435000000
1!
1%
#206440000000
0!
0%
#206445000000
1!
1%
#206450000000
0!
0%
#206455000000
1!
1%
#206460000000
0!
0%
#206465000000
1!
1%
#206470000000
0!
0%
#206475000000
1!
1%
#206480000000
0!
0%
#206485000000
1!
1%
#206490000000
0!
0%
#206495000000
1!
1%
#206500000000
0!
0%
#206505000000
1!
1%
#206510000000
0!
0%
#206515000000
1!
1%
#206520000000
0!
0%
#206525000000
1!
1%
#206530000000
0!
0%
#206535000000
1!
1%
#206540000000
0!
0%
#206545000000
1!
1%
#206550000000
0!
0%
#206555000000
1!
1%
#206560000000
0!
0%
#206565000000
1!
1%
#206570000000
0!
0%
#206575000000
1!
1%
#206580000000
0!
0%
#206585000000
1!
1%
#206590000000
0!
0%
#206595000000
1!
1%
#206600000000
0!
0%
#206605000000
1!
1%
#206610000000
0!
0%
#206615000000
1!
1%
#206620000000
0!
0%
#206625000000
1!
1%
#206630000000
0!
0%
#206635000000
1!
1%
#206640000000
0!
0%
#206645000000
1!
1%
#206650000000
0!
0%
#206655000000
1!
1%
#206660000000
0!
0%
#206665000000
1!
1%
#206670000000
0!
0%
#206675000000
1!
1%
#206680000000
0!
0%
#206685000000
1!
1%
#206690000000
0!
0%
#206695000000
1!
1%
#206700000000
0!
0%
#206705000000
1!
1%
#206710000000
0!
0%
#206715000000
1!
1%
#206720000000
0!
0%
#206725000000
1!
1%
#206730000000
0!
0%
#206735000000
1!
1%
#206740000000
0!
0%
#206745000000
1!
1%
#206750000000
0!
0%
#206755000000
1!
1%
#206760000000
0!
0%
#206765000000
1!
1%
#206770000000
0!
0%
#206775000000
1!
1%
#206780000000
0!
0%
#206785000000
1!
1%
#206790000000
0!
0%
#206795000000
1!
1%
#206800000000
0!
0%
#206805000000
1!
1%
#206810000000
0!
0%
#206815000000
1!
1%
#206820000000
0!
0%
#206825000000
1!
1%
#206830000000
0!
0%
#206835000000
1!
1%
#206840000000
0!
0%
#206845000000
1!
1%
#206850000000
0!
0%
#206855000000
1!
1%
#206860000000
0!
0%
#206865000000
1!
1%
#206870000000
0!
0%
#206875000000
1!
1%
#206880000000
0!
0%
#206885000000
1!
1%
#206890000000
0!
0%
#206895000000
1!
1%
#206900000000
0!
0%
#206905000000
1!
1%
#206910000000
0!
0%
#206915000000
1!
1%
#206920000000
0!
0%
#206925000000
1!
1%
#206930000000
0!
0%
#206935000000
1!
1%
#206940000000
0!
0%
#206945000000
1!
1%
#206950000000
0!
0%
#206955000000
1!
1%
#206960000000
0!
0%
#206965000000
1!
1%
#206970000000
0!
0%
#206975000000
1!
1%
#206980000000
0!
0%
#206985000000
1!
1%
#206990000000
0!
0%
#206995000000
1!
1%
#207000000000
0!
0%
#207005000000
1!
1%
#207010000000
0!
0%
#207015000000
1!
1%
#207020000000
0!
0%
#207025000000
1!
1%
#207030000000
0!
0%
#207035000000
1!
1%
#207040000000
0!
0%
#207045000000
1!
1%
#207050000000
0!
0%
#207055000000
1!
1%
#207060000000
0!
0%
#207065000000
1!
1%
#207070000000
0!
0%
#207075000000
1!
1%
#207080000000
0!
0%
#207085000000
1!
1%
#207090000000
0!
0%
#207095000000
1!
1%
#207100000000
0!
0%
#207105000000
1!
1%
#207110000000
0!
0%
#207115000000
1!
1%
#207120000000
0!
0%
#207125000000
1!
1%
#207130000000
0!
0%
#207135000000
1!
1%
#207140000000
0!
0%
#207145000000
1!
1%
#207150000000
0!
0%
#207155000000
1!
1%
#207160000000
0!
0%
#207165000000
1!
1%
#207170000000
0!
0%
#207175000000
1!
1%
#207180000000
0!
0%
#207185000000
1!
1%
#207190000000
0!
0%
#207195000000
1!
1%
#207200000000
0!
0%
#207205000000
1!
1%
#207210000000
0!
0%
#207215000000
1!
1%
#207220000000
0!
0%
#207225000000
1!
1%
#207230000000
0!
0%
#207235000000
1!
1%
#207240000000
0!
0%
#207245000000
1!
1%
#207250000000
0!
0%
#207255000000
1!
1%
#207260000000
0!
0%
#207265000000
1!
1%
#207270000000
0!
0%
#207275000000
1!
1%
#207280000000
0!
0%
#207285000000
1!
1%
#207290000000
0!
0%
#207295000000
1!
1%
#207300000000
0!
0%
#207305000000
1!
1%
#207310000000
0!
0%
#207315000000
1!
1%
#207320000000
0!
0%
#207325000000
1!
1%
#207330000000
0!
0%
#207335000000
1!
1%
#207340000000
0!
0%
#207345000000
1!
1%
#207350000000
0!
0%
#207355000000
1!
1%
#207360000000
0!
0%
#207365000000
1!
1%
#207370000000
0!
0%
#207375000000
1!
1%
#207380000000
0!
0%
#207385000000
1!
1%
#207390000000
0!
0%
#207395000000
1!
1%
#207400000000
0!
0%
#207405000000
1!
1%
#207410000000
0!
0%
#207415000000
1!
1%
#207420000000
0!
0%
#207425000000
1!
1%
#207430000000
0!
0%
#207435000000
1!
1%
#207440000000
0!
0%
#207445000000
1!
1%
#207450000000
0!
0%
#207455000000
1!
1%
#207460000000
0!
0%
#207465000000
1!
1%
#207470000000
0!
0%
#207475000000
1!
1%
#207480000000
0!
0%
#207485000000
1!
1%
#207490000000
0!
0%
#207495000000
1!
1%
#207500000000
0!
0%
#207505000000
1!
1%
#207510000000
0!
0%
#207515000000
1!
1%
#207520000000
0!
0%
#207525000000
1!
1%
#207530000000
0!
0%
#207535000000
1!
1%
#207540000000
0!
0%
#207545000000
1!
1%
#207550000000
0!
0%
#207555000000
1!
1%
#207560000000
0!
0%
#207565000000
1!
1%
#207570000000
0!
0%
#207575000000
1!
1%
#207580000000
0!
0%
#207585000000
1!
1%
#207590000000
0!
0%
#207595000000
1!
1%
#207600000000
0!
0%
#207605000000
1!
1%
#207610000000
0!
0%
#207615000000
1!
1%
#207620000000
0!
0%
#207625000000
1!
1%
#207630000000
0!
0%
#207635000000
1!
1%
#207640000000
0!
0%
#207645000000
1!
1%
#207650000000
0!
0%
#207655000000
1!
1%
#207660000000
0!
0%
#207665000000
1!
1%
#207670000000
0!
0%
#207675000000
1!
1%
#207680000000
0!
0%
#207685000000
1!
1%
#207690000000
0!
0%
#207695000000
1!
1%
#207700000000
0!
0%
#207705000000
1!
1%
#207710000000
0!
0%
#207715000000
1!
1%
#207720000000
0!
0%
#207725000000
1!
1%
#207730000000
0!
0%
#207735000000
1!
1%
#207740000000
0!
0%
#207745000000
1!
1%
#207750000000
0!
0%
#207755000000
1!
1%
#207760000000
0!
0%
#207765000000
1!
1%
#207770000000
0!
0%
#207775000000
1!
1%
#207780000000
0!
0%
#207785000000
1!
1%
#207790000000
0!
0%
#207795000000
1!
1%
#207800000000
0!
0%
#207805000000
1!
1%
#207810000000
0!
0%
#207815000000
1!
1%
#207820000000
0!
0%
#207825000000
1!
1%
#207830000000
0!
0%
#207835000000
1!
1%
#207840000000
0!
0%
#207845000000
1!
1%
#207850000000
0!
0%
#207855000000
1!
1%
#207860000000
0!
0%
#207865000000
1!
1%
#207870000000
0!
0%
#207875000000
1!
1%
#207880000000
0!
0%
#207885000000
1!
1%
#207890000000
0!
0%
#207895000000
1!
1%
#207900000000
0!
0%
#207905000000
1!
1%
#207910000000
0!
0%
#207915000000
1!
1%
#207920000000
0!
0%
#207925000000
1!
1%
#207930000000
0!
0%
#207935000000
1!
1%
#207940000000
0!
0%
#207945000000
1!
1%
#207950000000
0!
0%
#207955000000
1!
1%
#207960000000
0!
0%
#207965000000
1!
1%
#207970000000
0!
0%
#207975000000
1!
1%
#207980000000
0!
0%
#207985000000
1!
1%
#207990000000
0!
0%
#207995000000
1!
1%
#208000000000
0!
0%
#208005000000
1!
1%
#208010000000
0!
0%
#208015000000
1!
1%
#208020000000
0!
0%
#208025000000
1!
1%
#208030000000
0!
0%
#208035000000
1!
1%
#208040000000
0!
0%
#208045000000
1!
1%
#208050000000
0!
0%
#208055000000
1!
1%
#208060000000
0!
0%
#208065000000
1!
1%
#208070000000
0!
0%
#208075000000
1!
1%
#208080000000
0!
0%
#208085000000
1!
1%
#208090000000
0!
0%
#208095000000
1!
1%
#208100000000
0!
0%
#208105000000
1!
1%
#208110000000
0!
0%
#208115000000
1!
1%
#208120000000
0!
0%
#208125000000
1!
1%
#208130000000
0!
0%
#208135000000
1!
1%
#208140000000
0!
0%
#208145000000
1!
1%
#208150000000
0!
0%
#208155000000
1!
1%
#208160000000
0!
0%
#208165000000
1!
1%
#208170000000
0!
0%
#208175000000
1!
1%
#208180000000
0!
0%
#208185000000
1!
1%
#208190000000
0!
0%
#208195000000
1!
1%
#208200000000
0!
0%
#208205000000
1!
1%
#208210000000
0!
0%
#208215000000
1!
1%
#208220000000
0!
0%
#208225000000
1!
1%
#208230000000
0!
0%
#208235000000
1!
1%
#208240000000
0!
0%
#208245000000
1!
1%
#208250000000
0!
0%
#208255000000
1!
1%
#208260000000
0!
0%
#208265000000
1!
1%
#208270000000
0!
0%
#208275000000
1!
1%
#208280000000
0!
0%
#208285000000
1!
1%
#208290000000
0!
0%
#208295000000
1!
1%
#208300000000
0!
0%
#208305000000
1!
1%
#208310000000
0!
0%
#208315000000
1!
1%
#208320000000
0!
0%
#208325000000
1!
1%
#208330000000
0!
0%
#208335000000
1!
1%
#208340000000
0!
0%
#208345000000
1!
1%
#208350000000
0!
0%
#208355000000
1!
1%
#208360000000
0!
0%
#208365000000
1!
1%
#208370000000
0!
0%
#208375000000
1!
1%
#208380000000
0!
0%
#208385000000
1!
1%
#208390000000
0!
0%
#208395000000
1!
1%
#208400000000
0!
0%
#208405000000
1!
1%
#208410000000
0!
0%
#208415000000
1!
1%
#208420000000
0!
0%
#208425000000
1!
1%
#208430000000
0!
0%
#208435000000
1!
1%
#208440000000
0!
0%
#208445000000
1!
1%
#208450000000
0!
0%
#208455000000
1!
1%
#208460000000
0!
0%
#208465000000
1!
1%
#208470000000
0!
0%
#208475000000
1!
1%
#208480000000
0!
0%
#208485000000
1!
1%
#208490000000
0!
0%
#208495000000
1!
1%
#208500000000
0!
0%
#208505000000
1!
1%
#208510000000
0!
0%
#208515000000
1!
1%
#208520000000
0!
0%
#208525000000
1!
1%
#208530000000
0!
0%
#208535000000
1!
1%
#208540000000
0!
0%
#208545000000
1!
1%
#208550000000
0!
0%
#208555000000
1!
1%
#208560000000
0!
0%
#208565000000
1!
1%
#208570000000
0!
0%
#208575000000
1!
1%
#208580000000
0!
0%
#208585000000
1!
1%
#208590000000
0!
0%
#208595000000
1!
1%
#208600000000
0!
0%
#208605000000
1!
1%
#208610000000
0!
0%
#208615000000
1!
1%
#208620000000
0!
0%
#208625000000
1!
1%
#208630000000
0!
0%
#208635000000
1!
1%
#208640000000
0!
0%
#208645000000
1!
1%
#208650000000
0!
0%
#208655000000
1!
1%
#208660000000
0!
0%
#208665000000
1!
1%
#208670000000
0!
0%
#208675000000
1!
1%
#208680000000
0!
0%
#208685000000
1!
1%
#208690000000
0!
0%
#208695000000
1!
1%
#208700000000
0!
0%
#208705000000
1!
1%
#208710000000
0!
0%
#208715000000
1!
1%
#208720000000
0!
0%
#208725000000
1!
1%
#208730000000
0!
0%
#208735000000
1!
1%
#208740000000
0!
0%
#208745000000
1!
1%
#208750000000
0!
0%
#208755000000
1!
1%
#208760000000
0!
0%
#208765000000
1!
1%
#208770000000
0!
0%
#208775000000
1!
1%
#208780000000
0!
0%
#208785000000
1!
1%
#208790000000
0!
0%
#208795000000
1!
1%
#208800000000
0!
0%
#208805000000
1!
1%
#208810000000
0!
0%
#208815000000
1!
1%
#208820000000
0!
0%
#208825000000
1!
1%
#208830000000
0!
0%
#208835000000
1!
1%
#208840000000
0!
0%
#208845000000
1!
1%
#208850000000
0!
0%
#208855000000
1!
1%
#208860000000
0!
0%
#208865000000
1!
1%
#208870000000
0!
0%
#208875000000
1!
1%
#208880000000
0!
0%
#208885000000
1!
1%
#208890000000
0!
0%
#208895000000
1!
1%
#208900000000
0!
0%
#208905000000
1!
1%
#208910000000
0!
0%
#208915000000
1!
1%
#208920000000
0!
0%
#208925000000
1!
1%
#208930000000
0!
0%
#208935000000
1!
1%
#208940000000
0!
0%
#208945000000
1!
1%
#208950000000
0!
0%
#208955000000
1!
1%
#208960000000
0!
0%
#208965000000
1!
1%
#208970000000
0!
0%
#208975000000
1!
1%
#208980000000
0!
0%
#208985000000
1!
1%
#208990000000
0!
0%
#208995000000
1!
1%
#209000000000
0!
0%
#209005000000
1!
1%
#209010000000
0!
0%
#209015000000
1!
1%
#209020000000
0!
0%
#209025000000
1!
1%
#209030000000
0!
0%
#209035000000
1!
1%
#209040000000
0!
0%
#209045000000
1!
1%
#209050000000
0!
0%
#209055000000
1!
1%
#209060000000
0!
0%
#209065000000
1!
1%
#209070000000
0!
0%
#209075000000
1!
1%
#209080000000
0!
0%
#209085000000
1!
1%
#209090000000
0!
0%
#209095000000
1!
1%
#209100000000
0!
0%
#209105000000
1!
1%
#209110000000
0!
0%
#209115000000
1!
1%
#209120000000
0!
0%
#209125000000
1!
1%
#209130000000
0!
0%
#209135000000
1!
1%
#209140000000
0!
0%
#209145000000
1!
1%
#209150000000
0!
0%
#209155000000
1!
1%
#209160000000
0!
0%
#209165000000
1!
1%
#209170000000
0!
0%
#209175000000
1!
1%
#209180000000
0!
0%
#209185000000
1!
1%
#209190000000
0!
0%
#209195000000
1!
1%
#209200000000
0!
0%
#209205000000
1!
1%
#209210000000
0!
0%
#209215000000
1!
1%
#209220000000
0!
0%
#209225000000
1!
1%
#209230000000
0!
0%
#209235000000
1!
1%
#209240000000
0!
0%
#209245000000
1!
1%
#209250000000
0!
0%
#209255000000
1!
1%
#209260000000
0!
0%
#209265000000
1!
1%
#209270000000
0!
0%
#209275000000
1!
1%
#209280000000
0!
0%
#209285000000
1!
1%
#209290000000
0!
0%
#209295000000
1!
1%
#209300000000
0!
0%
#209305000000
1!
1%
#209310000000
0!
0%
#209315000000
1!
1%
#209320000000
0!
0%
#209325000000
1!
1%
#209330000000
0!
0%
#209335000000
1!
1%
#209340000000
0!
0%
#209345000000
1!
1%
#209350000000
0!
0%
#209355000000
1!
1%
#209360000000
0!
0%
#209365000000
1!
1%
#209370000000
0!
0%
#209375000000
1!
1%
#209380000000
0!
0%
#209385000000
1!
1%
#209390000000
0!
0%
#209395000000
1!
1%
#209400000000
0!
0%
#209405000000
1!
1%
#209410000000
0!
0%
#209415000000
1!
1%
#209420000000
0!
0%
#209425000000
1!
1%
#209430000000
0!
0%
#209435000000
1!
1%
#209440000000
0!
0%
#209445000000
1!
1%
#209450000000
0!
0%
#209455000000
1!
1%
#209460000000
0!
0%
#209465000000
1!
1%
#209470000000
0!
0%
#209475000000
1!
1%
#209480000000
0!
0%
#209485000000
1!
1%
#209490000000
0!
0%
#209495000000
1!
1%
#209500000000
0!
0%
#209505000000
1!
1%
#209510000000
0!
0%
#209515000000
1!
1%
#209520000000
0!
0%
#209525000000
1!
1%
#209530000000
0!
0%
#209535000000
1!
1%
#209540000000
0!
0%
#209545000000
1!
1%
#209550000000
0!
0%
#209555000000
1!
1%
#209560000000
0!
0%
#209565000000
1!
1%
#209570000000
0!
0%
#209575000000
1!
1%
#209580000000
0!
0%
#209585000000
1!
1%
#209590000000
0!
0%
#209595000000
1!
1%
#209600000000
0!
0%
#209605000000
1!
1%
#209610000000
0!
0%
#209615000000
1!
1%
#209620000000
0!
0%
#209625000000
1!
1%
#209630000000
0!
0%
#209635000000
1!
1%
#209640000000
0!
0%
#209645000000
1!
1%
#209650000000
0!
0%
#209655000000
1!
1%
#209660000000
0!
0%
#209665000000
1!
1%
#209670000000
0!
0%
#209675000000
1!
1%
#209680000000
0!
0%
#209685000000
1!
1%
#209690000000
0!
0%
#209695000000
1!
1%
#209700000000
0!
0%
#209705000000
1!
1%
#209710000000
0!
0%
#209715000000
1!
1%
#209720000000
0!
0%
#209725000000
1!
1%
#209730000000
0!
0%
#209735000000
1!
1%
#209740000000
0!
0%
#209745000000
1!
1%
#209750000000
0!
0%
#209755000000
1!
1%
#209760000000
0!
0%
#209765000000
1!
1%
#209770000000
0!
0%
#209775000000
1!
1%
#209780000000
0!
0%
#209785000000
1!
1%
#209790000000
0!
0%
#209795000000
1!
1%
#209800000000
0!
0%
#209805000000
1!
1%
#209810000000
0!
0%
#209815000000
1!
1%
#209820000000
0!
0%
#209825000000
1!
1%
#209830000000
0!
0%
#209835000000
1!
1%
#209840000000
0!
0%
#209845000000
1!
1%
#209850000000
0!
0%
#209855000000
1!
1%
#209860000000
0!
0%
#209865000000
1!
1%
#209870000000
0!
0%
#209875000000
1!
1%
#209880000000
0!
0%
#209885000000
1!
1%
#209890000000
0!
0%
#209895000000
1!
1%
#209900000000
0!
0%
#209905000000
1!
1%
#209910000000
0!
0%
#209915000000
1!
1%
#209920000000
0!
0%
#209925000000
1!
1%
#209930000000
0!
0%
#209935000000
1!
1%
#209940000000
0!
0%
#209945000000
1!
1%
#209950000000
0!
0%
#209955000000
1!
1%
#209960000000
0!
0%
#209965000000
1!
1%
#209970000000
0!
0%
#209975000000
1!
1%
#209980000000
0!
0%
#209985000000
1!
1%
#209990000000
0!
0%
#209995000000
1!
1%
#210000000000
0!
0%
#210005000000
1!
1%
#210010000000
0!
0%
#210015000000
1!
1%
#210020000000
0!
0%
#210025000000
1!
1%
#210030000000
0!
0%
#210035000000
1!
1%
#210040000000
0!
0%
#210045000000
1!
1%
#210050000000
0!
0%
#210055000000
1!
1%
#210060000000
0!
0%
#210065000000
1!
1%
#210070000000
0!
0%
#210075000000
1!
1%
#210080000000
0!
0%
#210085000000
1!
1%
#210090000000
0!
0%
#210095000000
1!
1%
#210100000000
0!
0%
#210105000000
1!
1%
#210110000000
0!
0%
#210115000000
1!
1%
#210120000000
0!
0%
#210125000000
1!
1%
#210130000000
0!
0%
#210135000000
1!
1%
#210140000000
0!
0%
#210145000000
1!
1%
#210150000000
0!
0%
#210155000000
1!
1%
#210160000000
0!
0%
#210165000000
1!
1%
#210170000000
0!
0%
#210175000000
1!
1%
#210180000000
0!
0%
#210185000000
1!
1%
#210190000000
0!
0%
#210195000000
1!
1%
#210200000000
0!
0%
#210205000000
1!
1%
#210210000000
0!
0%
#210215000000
1!
1%
#210220000000
0!
0%
#210225000000
1!
1%
#210230000000
0!
0%
#210235000000
1!
1%
#210240000000
0!
0%
#210245000000
1!
1%
#210250000000
0!
0%
#210255000000
1!
1%
#210260000000
0!
0%
#210265000000
1!
1%
#210270000000
0!
0%
#210275000000
1!
1%
#210280000000
0!
0%
#210285000000
1!
1%
#210290000000
0!
0%
#210295000000
1!
1%
#210300000000
0!
0%
#210305000000
1!
1%
#210310000000
0!
0%
#210315000000
1!
1%
#210320000000
0!
0%
#210325000000
1!
1%
#210330000000
0!
0%
#210335000000
1!
1%
#210340000000
0!
0%
#210345000000
1!
1%
#210350000000
0!
0%
#210355000000
1!
1%
#210360000000
0!
0%
#210365000000
1!
1%
#210370000000
0!
0%
#210375000000
1!
1%
#210380000000
0!
0%
#210385000000
1!
1%
#210390000000
0!
0%
#210395000000
1!
1%
#210400000000
0!
0%
#210405000000
1!
1%
#210410000000
0!
0%
#210415000000
1!
1%
#210420000000
0!
0%
#210425000000
1!
1%
#210430000000
0!
0%
#210435000000
1!
1%
#210440000000
0!
0%
#210445000000
1!
1%
#210450000000
0!
0%
#210455000000
1!
1%
#210460000000
0!
0%
#210465000000
1!
1%
#210470000000
0!
0%
#210475000000
1!
1%
#210480000000
0!
0%
#210485000000
1!
1%
#210490000000
0!
0%
#210495000000
1!
1%
#210500000000
0!
0%
#210505000000
1!
1%
#210510000000
0!
0%
#210515000000
1!
1%
#210520000000
0!
0%
#210525000000
1!
1%
#210530000000
0!
0%
#210535000000
1!
1%
#210540000000
0!
0%
#210545000000
1!
1%
#210550000000
0!
0%
#210555000000
1!
1%
#210560000000
0!
0%
#210565000000
1!
1%
#210570000000
0!
0%
#210575000000
1!
1%
#210580000000
0!
0%
#210585000000
1!
1%
#210590000000
0!
0%
#210595000000
1!
1%
#210600000000
0!
0%
#210605000000
1!
1%
#210610000000
0!
0%
#210615000000
1!
1%
#210620000000
0!
0%
#210625000000
1!
1%
#210630000000
0!
0%
#210635000000
1!
1%
#210640000000
0!
0%
#210645000000
1!
1%
#210650000000
0!
0%
#210655000000
1!
1%
#210660000000
0!
0%
#210665000000
1!
1%
#210670000000
0!
0%
#210675000000
1!
1%
#210680000000
0!
0%
#210685000000
1!
1%
#210690000000
0!
0%
#210695000000
1!
1%
#210700000000
0!
0%
#210705000000
1!
1%
#210710000000
0!
0%
#210715000000
1!
1%
#210720000000
0!
0%
#210725000000
1!
1%
#210730000000
0!
0%
#210735000000
1!
1%
#210740000000
0!
0%
#210745000000
1!
1%
#210750000000
0!
0%
#210755000000
1!
1%
#210760000000
0!
0%
#210765000000
1!
1%
#210770000000
0!
0%
#210775000000
1!
1%
#210780000000
0!
0%
#210785000000
1!
1%
#210790000000
0!
0%
#210795000000
1!
1%
#210800000000
0!
0%
#210805000000
1!
1%
#210810000000
0!
0%
#210815000000
1!
1%
#210820000000
0!
0%
#210825000000
1!
1%
#210830000000
0!
0%
#210835000000
1!
1%
#210840000000
0!
0%
#210845000000
1!
1%
#210850000000
0!
0%
#210855000000
1!
1%
#210860000000
0!
0%
#210865000000
1!
1%
#210870000000
0!
0%
#210875000000
1!
1%
#210880000000
0!
0%
#210885000000
1!
1%
#210890000000
0!
0%
#210895000000
1!
1%
#210900000000
0!
0%
#210905000000
1!
1%
#210910000000
0!
0%
#210915000000
1!
1%
#210920000000
0!
0%
#210925000000
1!
1%
#210930000000
0!
0%
#210935000000
1!
1%
#210940000000
0!
0%
#210945000000
1!
1%
#210950000000
0!
0%
#210955000000
1!
1%
#210960000000
0!
0%
#210965000000
1!
1%
#210970000000
0!
0%
#210975000000
1!
1%
#210980000000
0!
0%
#210985000000
1!
1%
#210990000000
0!
0%
#210995000000
1!
1%
#211000000000
0!
0%
#211005000000
1!
1%
#211010000000
0!
0%
#211015000000
1!
1%
#211020000000
0!
0%
#211025000000
1!
1%
#211030000000
0!
0%
#211035000000
1!
1%
#211040000000
0!
0%
#211045000000
1!
1%
#211050000000
0!
0%
#211055000000
1!
1%
#211060000000
0!
0%
#211065000000
1!
1%
#211070000000
0!
0%
#211075000000
1!
1%
#211080000000
0!
0%
#211085000000
1!
1%
#211090000000
0!
0%
#211095000000
1!
1%
#211100000000
0!
0%
#211105000000
1!
1%
#211110000000
0!
0%
#211115000000
1!
1%
#211120000000
0!
0%
#211125000000
1!
1%
#211130000000
0!
0%
#211135000000
1!
1%
#211140000000
0!
0%
#211145000000
1!
1%
#211150000000
0!
0%
#211155000000
1!
1%
#211160000000
0!
0%
#211165000000
1!
1%
#211170000000
0!
0%
#211175000000
1!
1%
#211180000000
0!
0%
#211185000000
1!
1%
#211190000000
0!
0%
#211195000000
1!
1%
#211200000000
0!
0%
#211205000000
1!
1%
#211210000000
0!
0%
#211215000000
1!
1%
#211220000000
0!
0%
#211225000000
1!
1%
#211230000000
0!
0%
#211235000000
1!
1%
#211240000000
0!
0%
#211245000000
1!
1%
#211250000000
0!
0%
#211255000000
1!
1%
#211260000000
0!
0%
#211265000000
1!
1%
#211270000000
0!
0%
#211275000000
1!
1%
#211280000000
0!
0%
#211285000000
1!
1%
#211290000000
0!
0%
#211295000000
1!
1%
#211300000000
0!
0%
#211305000000
1!
1%
#211310000000
0!
0%
#211315000000
1!
1%
#211320000000
0!
0%
#211325000000
1!
1%
#211330000000
0!
0%
#211335000000
1!
1%
#211340000000
0!
0%
#211345000000
1!
1%
#211350000000
0!
0%
#211355000000
1!
1%
#211360000000
0!
0%
#211365000000
1!
1%
#211370000000
0!
0%
#211375000000
1!
1%
#211380000000
0!
0%
#211385000000
1!
1%
#211390000000
0!
0%
#211395000000
1!
1%
#211400000000
0!
0%
#211405000000
1!
1%
#211410000000
0!
0%
#211415000000
1!
1%
#211420000000
0!
0%
#211425000000
1!
1%
#211430000000
0!
0%
#211435000000
1!
1%
#211440000000
0!
0%
#211445000000
1!
1%
#211450000000
0!
0%
#211455000000
1!
1%
#211460000000
0!
0%
#211465000000
1!
1%
#211470000000
0!
0%
#211475000000
1!
1%
#211480000000
0!
0%
#211485000000
1!
1%
#211490000000
0!
0%
#211495000000
1!
1%
#211500000000
0!
0%
#211505000000
1!
1%
#211510000000
0!
0%
#211515000000
1!
1%
#211520000000
0!
0%
#211525000000
1!
1%
#211530000000
0!
0%
#211535000000
1!
1%
#211540000000
0!
0%
#211545000000
1!
1%
#211550000000
0!
0%
#211555000000
1!
1%
#211560000000
0!
0%
#211565000000
1!
1%
#211570000000
0!
0%
#211575000000
1!
1%
#211580000000
0!
0%
#211585000000
1!
1%
#211590000000
0!
0%
#211595000000
1!
1%
#211600000000
0!
0%
#211605000000
1!
1%
#211610000000
0!
0%
#211615000000
1!
1%
#211620000000
0!
0%
#211625000000
1!
1%
#211630000000
0!
0%
#211635000000
1!
1%
#211640000000
0!
0%
#211645000000
1!
1%
#211650000000
0!
0%
#211655000000
1!
1%
#211660000000
0!
0%
#211665000000
1!
1%
#211670000000
0!
0%
#211675000000
1!
1%
#211680000000
0!
0%
#211685000000
1!
1%
#211690000000
0!
0%
#211695000000
1!
1%
#211700000000
0!
0%
#211705000000
1!
1%
#211710000000
0!
0%
#211715000000
1!
1%
#211720000000
0!
0%
#211725000000
1!
1%
#211730000000
0!
0%
#211735000000
1!
1%
#211740000000
0!
0%
#211745000000
1!
1%
#211750000000
0!
0%
#211755000000
1!
1%
#211760000000
0!
0%
#211765000000
1!
1%
#211770000000
0!
0%
#211775000000
1!
1%
#211780000000
0!
0%
#211785000000
1!
1%
#211790000000
0!
0%
#211795000000
1!
1%
#211800000000
0!
0%
#211805000000
1!
1%
#211810000000
0!
0%
#211815000000
1!
1%
#211820000000
0!
0%
#211825000000
1!
1%
#211830000000
0!
0%
#211835000000
1!
1%
#211840000000
0!
0%
#211845000000
1!
1%
#211850000000
0!
0%
#211855000000
1!
1%
#211860000000
0!
0%
#211865000000
1!
1%
#211870000000
0!
0%
#211875000000
1!
1%
#211880000000
0!
0%
#211885000000
1!
1%
#211890000000
0!
0%
#211895000000
1!
1%
#211900000000
0!
0%
#211905000000
1!
1%
#211910000000
0!
0%
#211915000000
1!
1%
#211920000000
0!
0%
#211925000000
1!
1%
#211930000000
0!
0%
#211935000000
1!
1%
#211940000000
0!
0%
#211945000000
1!
1%
#211950000000
0!
0%
#211955000000
1!
1%
#211960000000
0!
0%
#211965000000
1!
1%
#211970000000
0!
0%
#211975000000
1!
1%
#211980000000
0!
0%
#211985000000
1!
1%
#211990000000
0!
0%
#211995000000
1!
1%
#212000000000
0!
0%
#212005000000
1!
1%
#212010000000
0!
0%
#212015000000
1!
1%
#212020000000
0!
0%
#212025000000
1!
1%
#212030000000
0!
0%
#212035000000
1!
1%
#212040000000
0!
0%
#212045000000
1!
1%
#212050000000
0!
0%
#212055000000
1!
1%
#212060000000
0!
0%
#212065000000
1!
1%
#212070000000
0!
0%
#212075000000
1!
1%
#212080000000
0!
0%
#212085000000
1!
1%
#212090000000
0!
0%
#212095000000
1!
1%
#212100000000
0!
0%
#212105000000
1!
1%
#212110000000
0!
0%
#212115000000
1!
1%
#212120000000
0!
0%
#212125000000
1!
1%
#212130000000
0!
0%
#212135000000
1!
1%
#212140000000
0!
0%
#212145000000
1!
1%
#212150000000
0!
0%
#212155000000
1!
1%
#212160000000
0!
0%
#212165000000
1!
1%
#212170000000
0!
0%
#212175000000
1!
1%
#212180000000
0!
0%
#212185000000
1!
1%
#212190000000
0!
0%
#212195000000
1!
1%
#212200000000
0!
0%
#212205000000
1!
1%
#212210000000
0!
0%
#212215000000
1!
1%
#212220000000
0!
0%
#212225000000
1!
1%
#212230000000
0!
0%
#212235000000
1!
1%
#212240000000
0!
0%
#212245000000
1!
1%
#212250000000
0!
0%
#212255000000
1!
1%
#212260000000
0!
0%
#212265000000
1!
1%
#212270000000
0!
0%
#212275000000
1!
1%
#212280000000
0!
0%
#212285000000
1!
1%
#212290000000
0!
0%
#212295000000
1!
1%
#212300000000
0!
0%
#212305000000
1!
1%
#212310000000
0!
0%
#212315000000
1!
1%
#212320000000
0!
0%
#212325000000
1!
1%
#212330000000
0!
0%
#212335000000
1!
1%
#212340000000
0!
0%
#212345000000
1!
1%
#212350000000
0!
0%
#212355000000
1!
1%
#212360000000
0!
0%
#212365000000
1!
1%
#212370000000
0!
0%
#212375000000
1!
1%
#212380000000
0!
0%
#212385000000
1!
1%
#212390000000
0!
0%
#212395000000
1!
1%
#212400000000
0!
0%
#212405000000
1!
1%
#212410000000
0!
0%
#212415000000
1!
1%
#212420000000
0!
0%
#212425000000
1!
1%
#212430000000
0!
0%
#212435000000
1!
1%
#212440000000
0!
0%
#212445000000
1!
1%
#212450000000
0!
0%
#212455000000
1!
1%
#212460000000
0!
0%
#212465000000
1!
1%
#212470000000
0!
0%
#212475000000
1!
1%
#212480000000
0!
0%
#212485000000
1!
1%
#212490000000
0!
0%
#212495000000
1!
1%
#212500000000
0!
0%
#212505000000
1!
1%
#212510000000
0!
0%
#212515000000
1!
1%
#212520000000
0!
0%
#212525000000
1!
1%
#212530000000
0!
0%
#212535000000
1!
1%
#212540000000
0!
0%
#212545000000
1!
1%
#212550000000
0!
0%
#212555000000
1!
1%
#212560000000
0!
0%
#212565000000
1!
1%
#212570000000
0!
0%
#212575000000
1!
1%
#212580000000
0!
0%
#212585000000
1!
1%
#212590000000
0!
0%
#212595000000
1!
1%
#212600000000
0!
0%
#212605000000
1!
1%
#212610000000
0!
0%
#212615000000
1!
1%
#212620000000
0!
0%
#212625000000
1!
1%
#212630000000
0!
0%
#212635000000
1!
1%
#212640000000
0!
0%
#212645000000
1!
1%
#212650000000
0!
0%
#212655000000
1!
1%
#212660000000
0!
0%
#212665000000
1!
1%
#212670000000
0!
0%
#212675000000
1!
1%
#212680000000
0!
0%
#212685000000
1!
1%
#212690000000
0!
0%
#212695000000
1!
1%
#212700000000
0!
0%
#212705000000
1!
1%
#212710000000
0!
0%
#212715000000
1!
1%
#212720000000
0!
0%
#212725000000
1!
1%
#212730000000
0!
0%
#212735000000
1!
1%
#212740000000
0!
0%
#212745000000
1!
1%
#212750000000
0!
0%
#212755000000
1!
1%
#212760000000
0!
0%
#212765000000
1!
1%
#212770000000
0!
0%
#212775000000
1!
1%
#212780000000
0!
0%
#212785000000
1!
1%
#212790000000
0!
0%
#212795000000
1!
1%
#212800000000
0!
0%
#212805000000
1!
1%
#212810000000
0!
0%
#212815000000
1!
1%
#212820000000
0!
0%
#212825000000
1!
1%
#212830000000
0!
0%
#212835000000
1!
1%
#212840000000
0!
0%
#212845000000
1!
1%
#212850000000
0!
0%
#212855000000
1!
1%
#212860000000
0!
0%
#212865000000
1!
1%
#212870000000
0!
0%
#212875000000
1!
1%
#212880000000
0!
0%
#212885000000
1!
1%
#212890000000
0!
0%
#212895000000
1!
1%
#212900000000
0!
0%
#212905000000
1!
1%
#212910000000
0!
0%
#212915000000
1!
1%
#212920000000
0!
0%
#212925000000
1!
1%
#212930000000
0!
0%
#212935000000
1!
1%
#212940000000
0!
0%
#212945000000
1!
1%
#212950000000
0!
0%
#212955000000
1!
1%
#212960000000
0!
0%
#212965000000
1!
1%
#212970000000
0!
0%
#212975000000
1!
1%
#212980000000
0!
0%
#212985000000
1!
1%
#212990000000
0!
0%
#212995000000
1!
1%
#213000000000
0!
0%
#213005000000
1!
1%
#213010000000
0!
0%
#213015000000
1!
1%
#213020000000
0!
0%
#213025000000
1!
1%
#213030000000
0!
0%
#213035000000
1!
1%
#213040000000
0!
0%
#213045000000
1!
1%
#213050000000
0!
0%
#213055000000
1!
1%
#213060000000
0!
0%
#213065000000
1!
1%
#213070000000
0!
0%
#213075000000
1!
1%
#213080000000
0!
0%
#213085000000
1!
1%
#213090000000
0!
0%
#213095000000
1!
1%
#213100000000
0!
0%
#213105000000
1!
1%
#213110000000
0!
0%
#213115000000
1!
1%
#213120000000
0!
0%
#213125000000
1!
1%
#213130000000
0!
0%
#213135000000
1!
1%
#213140000000
0!
0%
#213145000000
1!
1%
#213150000000
0!
0%
#213155000000
1!
1%
#213160000000
0!
0%
#213165000000
1!
1%
#213170000000
0!
0%
#213175000000
1!
1%
#213180000000
0!
0%
#213185000000
1!
1%
#213190000000
0!
0%
#213195000000
1!
1%
#213200000000
0!
0%
#213205000000
1!
1%
#213210000000
0!
0%
#213215000000
1!
1%
#213220000000
0!
0%
#213225000000
1!
1%
#213230000000
0!
0%
#213235000000
1!
1%
#213240000000
0!
0%
#213245000000
1!
1%
#213250000000
0!
0%
#213255000000
1!
1%
#213260000000
0!
0%
#213265000000
1!
1%
#213270000000
0!
0%
#213275000000
1!
1%
#213280000000
0!
0%
#213285000000
1!
1%
#213290000000
0!
0%
#213295000000
1!
1%
#213300000000
0!
0%
#213305000000
1!
1%
#213310000000
0!
0%
#213315000000
1!
1%
#213320000000
0!
0%
#213325000000
1!
1%
#213330000000
0!
0%
#213335000000
1!
1%
#213340000000
0!
0%
#213345000000
1!
1%
#213350000000
0!
0%
#213355000000
1!
1%
#213360000000
0!
0%
#213365000000
1!
1%
#213370000000
0!
0%
#213375000000
1!
1%
#213380000000
0!
0%
#213385000000
1!
1%
#213390000000
0!
0%
#213395000000
1!
1%
#213400000000
0!
0%
#213405000000
1!
1%
#213410000000
0!
0%
#213415000000
1!
1%
#213420000000
0!
0%
#213425000000
1!
1%
#213430000000
0!
0%
#213435000000
1!
1%
#213440000000
0!
0%
#213445000000
1!
1%
#213450000000
0!
0%
#213455000000
1!
1%
#213460000000
0!
0%
#213465000000
1!
1%
#213470000000
0!
0%
#213475000000
1!
1%
#213480000000
0!
0%
#213485000000
1!
1%
#213490000000
0!
0%
#213495000000
1!
1%
#213500000000
0!
0%
#213505000000
1!
1%
#213510000000
0!
0%
#213515000000
1!
1%
#213520000000
0!
0%
#213525000000
1!
1%
#213530000000
0!
0%
#213535000000
1!
1%
#213540000000
0!
0%
#213545000000
1!
1%
#213550000000
0!
0%
#213555000000
1!
1%
#213560000000
0!
0%
#213565000000
1!
1%
#213570000000
0!
0%
#213575000000
1!
1%
#213580000000
0!
0%
#213585000000
1!
1%
#213590000000
0!
0%
#213595000000
1!
1%
#213600000000
0!
0%
#213605000000
1!
1%
#213610000000
0!
0%
#213615000000
1!
1%
#213620000000
0!
0%
#213625000000
1!
1%
#213630000000
0!
0%
#213635000000
1!
1%
#213640000000
0!
0%
#213645000000
1!
1%
#213650000000
0!
0%
#213655000000
1!
1%
#213660000000
0!
0%
#213665000000
1!
1%
#213670000000
0!
0%
#213675000000
1!
1%
#213680000000
0!
0%
#213685000000
1!
1%
#213690000000
0!
0%
#213695000000
1!
1%
#213700000000
0!
0%
#213705000000
1!
1%
#213710000000
0!
0%
#213715000000
1!
1%
#213720000000
0!
0%
#213725000000
1!
1%
#213730000000
0!
0%
#213735000000
1!
1%
#213740000000
0!
0%
#213745000000
1!
1%
#213750000000
0!
0%
#213755000000
1!
1%
#213760000000
0!
0%
#213765000000
1!
1%
#213770000000
0!
0%
#213775000000
1!
1%
#213780000000
0!
0%
#213785000000
1!
1%
#213790000000
0!
0%
#213795000000
1!
1%
#213800000000
0!
0%
#213805000000
1!
1%
#213810000000
0!
0%
#213815000000
1!
1%
#213820000000
0!
0%
#213825000000
1!
1%
#213830000000
0!
0%
#213835000000
1!
1%
#213840000000
0!
0%
#213845000000
1!
1%
#213850000000
0!
0%
#213855000000
1!
1%
#213860000000
0!
0%
#213865000000
1!
1%
#213870000000
0!
0%
#213875000000
1!
1%
#213880000000
0!
0%
#213885000000
1!
1%
#213890000000
0!
0%
#213895000000
1!
1%
#213900000000
0!
0%
#213905000000
1!
1%
#213910000000
0!
0%
#213915000000
1!
1%
#213920000000
0!
0%
#213925000000
1!
1%
#213930000000
0!
0%
#213935000000
1!
1%
#213940000000
0!
0%
#213945000000
1!
1%
#213950000000
0!
0%
#213955000000
1!
1%
#213960000000
0!
0%
#213965000000
1!
1%
#213970000000
0!
0%
#213975000000
1!
1%
#213980000000
0!
0%
#213985000000
1!
1%
#213990000000
0!
0%
#213995000000
1!
1%
#214000000000
0!
0%
#214005000000
1!
1%
#214010000000
0!
0%
#214015000000
1!
1%
#214020000000
0!
0%
#214025000000
1!
1%
#214030000000
0!
0%
#214035000000
1!
1%
#214040000000
0!
0%
#214045000000
1!
1%
#214050000000
0!
0%
#214055000000
1!
1%
#214060000000
0!
0%
#214065000000
1!
1%
#214070000000
0!
0%
#214075000000
1!
1%
#214080000000
0!
0%
#214085000000
1!
1%
#214090000000
0!
0%
#214095000000
1!
1%
#214100000000
0!
0%
#214105000000
1!
1%
#214110000000
0!
0%
#214115000000
1!
1%
#214120000000
0!
0%
#214125000000
1!
1%
#214130000000
0!
0%
#214135000000
1!
1%
#214140000000
0!
0%
#214145000000
1!
1%
#214150000000
0!
0%
#214155000000
1!
1%
#214160000000
0!
0%
#214165000000
1!
1%
#214170000000
0!
0%
#214175000000
1!
1%
#214180000000
0!
0%
#214185000000
1!
1%
#214190000000
0!
0%
#214195000000
1!
1%
#214200000000
0!
0%
#214205000000
1!
1%
#214210000000
0!
0%
#214215000000
1!
1%
#214220000000
0!
0%
#214225000000
1!
1%
#214230000000
0!
0%
#214235000000
1!
1%
#214240000000
0!
0%
#214245000000
1!
1%
#214250000000
0!
0%
#214255000000
1!
1%
#214260000000
0!
0%
#214265000000
1!
1%
#214270000000
0!
0%
#214275000000
1!
1%
#214280000000
0!
0%
#214285000000
1!
1%
#214290000000
0!
0%
#214295000000
1!
1%
#214300000000
0!
0%
#214305000000
1!
1%
#214310000000
0!
0%
#214315000000
1!
1%
#214320000000
0!
0%
#214325000000
1!
1%
#214330000000
0!
0%
#214335000000
1!
1%
#214340000000
0!
0%
#214345000000
1!
1%
#214350000000
0!
0%
#214355000000
1!
1%
#214360000000
0!
0%
#214365000000
1!
1%
#214370000000
0!
0%
#214375000000
1!
1%
#214380000000
0!
0%
#214385000000
1!
1%
#214390000000
0!
0%
#214395000000
1!
1%
#214400000000
0!
0%
#214405000000
1!
1%
#214410000000
0!
0%
#214415000000
1!
1%
#214420000000
0!
0%
#214425000000
1!
1%
#214430000000
0!
0%
#214435000000
1!
1%
#214440000000
0!
0%
#214445000000
1!
1%
#214450000000
0!
0%
#214455000000
1!
1%
#214460000000
0!
0%
#214465000000
1!
1%
#214470000000
0!
0%
#214475000000
1!
1%
#214480000000
0!
0%
#214485000000
1!
1%
#214490000000
0!
0%
#214495000000
1!
1%
#214500000000
0!
0%
#214505000000
1!
1%
#214510000000
0!
0%
#214515000000
1!
1%
#214520000000
0!
0%
#214525000000
1!
1%
#214530000000
0!
0%
#214535000000
1!
1%
#214540000000
0!
0%
#214545000000
1!
1%
#214550000000
0!
0%
#214555000000
1!
1%
#214560000000
0!
0%
#214565000000
1!
1%
#214570000000
0!
0%
#214575000000
1!
1%
#214580000000
0!
0%
#214585000000
1!
1%
#214590000000
0!
0%
#214595000000
1!
1%
#214600000000
0!
0%
#214605000000
1!
1%
#214610000000
0!
0%
#214615000000
1!
1%
#214620000000
0!
0%
#214625000000
1!
1%
#214630000000
0!
0%
#214635000000
1!
1%
#214640000000
0!
0%
#214645000000
1!
1%
#214650000000
0!
0%
#214655000000
1!
1%
#214660000000
0!
0%
#214665000000
1!
1%
#214670000000
0!
0%
#214675000000
1!
1%
#214680000000
0!
0%
#214685000000
1!
1%
#214690000000
0!
0%
#214695000000
1!
1%
#214700000000
0!
0%
#214705000000
1!
1%
#214710000000
0!
0%
#214715000000
1!
1%
#214720000000
0!
0%
#214725000000
1!
1%
#214730000000
0!
0%
#214735000000
1!
1%
#214740000000
0!
0%
#214745000000
1!
1%
#214750000000
0!
0%
#214755000000
1!
1%
#214760000000
0!
0%
#214765000000
1!
1%
#214770000000
0!
0%
#214775000000
1!
1%
#214780000000
0!
0%
#214785000000
1!
1%
#214790000000
0!
0%
#214795000000
1!
1%
#214800000000
0!
0%
#214805000000
1!
1%
#214810000000
0!
0%
#214815000000
1!
1%
#214820000000
0!
0%
#214825000000
1!
1%
#214830000000
0!
0%
#214835000000
1!
1%
#214840000000
0!
0%
#214845000000
1!
1%
#214850000000
0!
0%
#214855000000
1!
1%
#214860000000
0!
0%
#214865000000
1!
1%
#214870000000
0!
0%
#214875000000
1!
1%
#214880000000
0!
0%
#214885000000
1!
1%
#214890000000
0!
0%
#214895000000
1!
1%
#214900000000
0!
0%
#214905000000
1!
1%
#214910000000
0!
0%
#214915000000
1!
1%
#214920000000
0!
0%
#214925000000
1!
1%
#214930000000
0!
0%
#214935000000
1!
1%
#214940000000
0!
0%
#214945000000
1!
1%
#214950000000
0!
0%
#214955000000
1!
1%
#214960000000
0!
0%
#214965000000
1!
1%
#214970000000
0!
0%
#214975000000
1!
1%
#214980000000
0!
0%
#214985000000
1!
1%
#214990000000
0!
0%
#214995000000
1!
1%
#215000000000
0!
0%
#215005000000
1!
1%
#215010000000
0!
0%
#215015000000
1!
1%
#215020000000
0!
0%
#215025000000
1!
1%
#215030000000
0!
0%
#215035000000
1!
1%
#215040000000
0!
0%
#215045000000
1!
1%
#215050000000
0!
0%
#215055000000
1!
1%
#215060000000
0!
0%
#215065000000
1!
1%
#215070000000
0!
0%
#215075000000
1!
1%
#215080000000
0!
0%
#215085000000
1!
1%
#215090000000
0!
0%
#215095000000
1!
1%
#215100000000
0!
0%
#215105000000
1!
1%
#215110000000
0!
0%
#215115000000
1!
1%
#215120000000
0!
0%
#215125000000
1!
1%
#215130000000
0!
0%
#215135000000
1!
1%
#215140000000
0!
0%
#215145000000
1!
1%
#215150000000
0!
0%
#215155000000
1!
1%
#215160000000
0!
0%
#215165000000
1!
1%
#215170000000
0!
0%
#215175000000
1!
1%
#215180000000
0!
0%
#215185000000
1!
1%
#215190000000
0!
0%
#215195000000
1!
1%
#215200000000
0!
0%
#215205000000
1!
1%
#215210000000
0!
0%
#215215000000
1!
1%
#215220000000
0!
0%
#215225000000
1!
1%
#215230000000
0!
0%
#215235000000
1!
1%
#215240000000
0!
0%
#215245000000
1!
1%
#215250000000
0!
0%
#215255000000
1!
1%
#215260000000
0!
0%
#215265000000
1!
1%
#215270000000
0!
0%
#215275000000
1!
1%
#215280000000
0!
0%
#215285000000
1!
1%
#215290000000
0!
0%
#215295000000
1!
1%
#215300000000
0!
0%
#215305000000
1!
1%
#215310000000
0!
0%
#215315000000
1!
1%
#215320000000
0!
0%
#215325000000
1!
1%
#215330000000
0!
0%
#215335000000
1!
1%
#215340000000
0!
0%
#215345000000
1!
1%
#215350000000
0!
0%
#215355000000
1!
1%
#215360000000
0!
0%
#215365000000
1!
1%
#215370000000
0!
0%
#215375000000
1!
1%
#215380000000
0!
0%
#215385000000
1!
1%
#215390000000
0!
0%
#215395000000
1!
1%
#215400000000
0!
0%
#215405000000
1!
1%
#215410000000
0!
0%
#215415000000
1!
1%
#215420000000
0!
0%
#215425000000
1!
1%
#215430000000
0!
0%
#215435000000
1!
1%
#215440000000
0!
0%
#215445000000
1!
1%
#215450000000
0!
0%
#215455000000
1!
1%
#215460000000
0!
0%
#215465000000
1!
1%
#215470000000
0!
0%
#215475000000
1!
1%
#215480000000
0!
0%
#215485000000
1!
1%
#215490000000
0!
0%
#215495000000
1!
1%
#215500000000
0!
0%
#215505000000
1!
1%
#215510000000
0!
0%
#215515000000
1!
1%
#215520000000
0!
0%
#215525000000
1!
1%
#215530000000
0!
0%
#215535000000
1!
1%
#215540000000
0!
0%
#215545000000
1!
1%
#215550000000
0!
0%
#215555000000
1!
1%
#215560000000
0!
0%
#215565000000
1!
1%
#215570000000
0!
0%
#215575000000
1!
1%
#215580000000
0!
0%
#215585000000
1!
1%
#215590000000
0!
0%
#215595000000
1!
1%
#215600000000
0!
0%
#215605000000
1!
1%
#215610000000
0!
0%
#215615000000
1!
1%
#215620000000
0!
0%
#215625000000
1!
1%
#215630000000
0!
0%
#215635000000
1!
1%
#215640000000
0!
0%
#215645000000
1!
1%
#215650000000
0!
0%
#215655000000
1!
1%
#215660000000
0!
0%
#215665000000
1!
1%
#215670000000
0!
0%
#215675000000
1!
1%
#215680000000
0!
0%
#215685000000
1!
1%
#215690000000
0!
0%
#215695000000
1!
1%
#215700000000
0!
0%
#215705000000
1!
1%
#215710000000
0!
0%
#215715000000
1!
1%
#215720000000
0!
0%
#215725000000
1!
1%
#215730000000
0!
0%
#215735000000
1!
1%
#215740000000
0!
0%
#215745000000
1!
1%
#215750000000
0!
0%
#215755000000
1!
1%
#215760000000
0!
0%
#215765000000
1!
1%
#215770000000
0!
0%
#215775000000
1!
1%
#215780000000
0!
0%
#215785000000
1!
1%
#215790000000
0!
0%
#215795000000
1!
1%
#215800000000
0!
0%
#215805000000
1!
1%
#215810000000
0!
0%
#215815000000
1!
1%
#215820000000
0!
0%
#215825000000
1!
1%
#215830000000
0!
0%
#215835000000
1!
1%
#215840000000
0!
0%
#215845000000
1!
1%
#215850000000
0!
0%
#215855000000
1!
1%
#215860000000
0!
0%
#215865000000
1!
1%
#215870000000
0!
0%
#215875000000
1!
1%
#215880000000
0!
0%
#215885000000
1!
1%
#215890000000
0!
0%
#215895000000
1!
1%
#215900000000
0!
0%
#215905000000
1!
1%
#215910000000
0!
0%
#215915000000
1!
1%
#215920000000
0!
0%
#215925000000
1!
1%
#215930000000
0!
0%
#215935000000
1!
1%
#215940000000
0!
0%
#215945000000
1!
1%
#215950000000
0!
0%
#215955000000
1!
1%
#215960000000
0!
0%
#215965000000
1!
1%
#215970000000
0!
0%
#215975000000
1!
1%
#215980000000
0!
0%
#215985000000
1!
1%
#215990000000
0!
0%
#215995000000
1!
1%
#216000000000
0!
0%
#216005000000
1!
1%
#216010000000
0!
0%
#216015000000
1!
1%
#216020000000
0!
0%
#216025000000
1!
1%
#216030000000
0!
0%
#216035000000
1!
1%
#216040000000
0!
0%
#216045000000
1!
1%
#216050000000
0!
0%
#216055000000
1!
1%
#216060000000
0!
0%
#216065000000
1!
1%
#216070000000
0!
0%
#216075000000
1!
1%
#216080000000
0!
0%
#216085000000
1!
1%
#216090000000
0!
0%
#216095000000
1!
1%
#216100000000
0!
0%
#216105000000
1!
1%
#216110000000
0!
0%
#216115000000
1!
1%
#216120000000
0!
0%
#216125000000
1!
1%
#216130000000
0!
0%
#216135000000
1!
1%
#216140000000
0!
0%
#216145000000
1!
1%
#216150000000
0!
0%
#216155000000
1!
1%
#216160000000
0!
0%
#216165000000
1!
1%
#216170000000
0!
0%
#216175000000
1!
1%
#216180000000
0!
0%
#216185000000
1!
1%
#216190000000
0!
0%
#216195000000
1!
1%
#216200000000
0!
0%
#216205000000
1!
1%
#216210000000
0!
0%
#216215000000
1!
1%
#216220000000
0!
0%
#216225000000
1!
1%
#216230000000
0!
0%
#216235000000
1!
1%
#216240000000
0!
0%
#216245000000
1!
1%
#216250000000
0!
0%
#216255000000
1!
1%
#216260000000
0!
0%
#216265000000
1!
1%
#216270000000
0!
0%
#216275000000
1!
1%
#216280000000
0!
0%
#216285000000
1!
1%
#216290000000
0!
0%
#216295000000
1!
1%
#216300000000
0!
0%
#216305000000
1!
1%
#216310000000
0!
0%
#216315000000
1!
1%
#216320000000
0!
0%
#216325000000
1!
1%
#216330000000
0!
0%
#216335000000
1!
1%
#216340000000
0!
0%
#216345000000
1!
1%
#216350000000
0!
0%
#216355000000
1!
1%
#216360000000
0!
0%
#216365000000
1!
1%
#216370000000
0!
0%
#216375000000
1!
1%
#216380000000
0!
0%
#216385000000
1!
1%
#216390000000
0!
0%
#216395000000
1!
1%
#216400000000
0!
0%
#216405000000
1!
1%
#216410000000
0!
0%
#216415000000
1!
1%
#216420000000
0!
0%
#216425000000
1!
1%
#216430000000
0!
0%
#216435000000
1!
1%
#216440000000
0!
0%
#216445000000
1!
1%
#216450000000
0!
0%
#216455000000
1!
1%
#216460000000
0!
0%
#216465000000
1!
1%
#216470000000
0!
0%
#216475000000
1!
1%
#216480000000
0!
0%
#216485000000
1!
1%
#216490000000
0!
0%
#216495000000
1!
1%
#216500000000
0!
0%
#216505000000
1!
1%
#216510000000
0!
0%
#216515000000
1!
1%
#216520000000
0!
0%
#216525000000
1!
1%
#216530000000
0!
0%
#216535000000
1!
1%
#216540000000
0!
0%
#216545000000
1!
1%
#216550000000
0!
0%
#216555000000
1!
1%
#216560000000
0!
0%
#216565000000
1!
1%
#216570000000
0!
0%
#216575000000
1!
1%
#216580000000
0!
0%
#216585000000
1!
1%
#216590000000
0!
0%
#216595000000
1!
1%
#216600000000
0!
0%
#216605000000
1!
1%
#216610000000
0!
0%
#216615000000
1!
1%
#216620000000
0!
0%
#216625000000
1!
1%
#216630000000
0!
0%
#216635000000
1!
1%
#216640000000
0!
0%
#216645000000
1!
1%
#216650000000
0!
0%
#216655000000
1!
1%
#216660000000
0!
0%
#216665000000
1!
1%
#216670000000
0!
0%
#216675000000
1!
1%
#216680000000
0!
0%
#216685000000
1!
1%
#216690000000
0!
0%
#216695000000
1!
1%
#216700000000
0!
0%
#216705000000
1!
1%
#216710000000
0!
0%
#216715000000
1!
1%
#216720000000
0!
0%
#216725000000
1!
1%
#216730000000
0!
0%
#216735000000
1!
1%
#216740000000
0!
0%
#216745000000
1!
1%
#216750000000
0!
0%
#216755000000
1!
1%
#216760000000
0!
0%
#216765000000
1!
1%
#216770000000
0!
0%
#216775000000
1!
1%
#216780000000
0!
0%
#216785000000
1!
1%
#216790000000
0!
0%
#216795000000
1!
1%
#216800000000
0!
0%
#216805000000
1!
1%
#216810000000
0!
0%
#216815000000
1!
1%
#216820000000
0!
0%
#216825000000
1!
1%
#216830000000
0!
0%
#216835000000
1!
1%
#216840000000
0!
0%
#216845000000
1!
1%
#216850000000
0!
0%
#216855000000
1!
1%
#216860000000
0!
0%
#216865000000
1!
1%
#216870000000
0!
0%
#216875000000
1!
1%
#216880000000
0!
0%
#216885000000
1!
1%
#216890000000
0!
0%
#216895000000
1!
1%
#216900000000
0!
0%
#216905000000
1!
1%
#216910000000
0!
0%
#216915000000
1!
1%
#216920000000
0!
0%
#216925000000
1!
1%
#216930000000
0!
0%
#216935000000
1!
1%
#216940000000
0!
0%
#216945000000
1!
1%
#216950000000
0!
0%
#216955000000
1!
1%
#216960000000
0!
0%
#216965000000
1!
1%
#216970000000
0!
0%
#216975000000
1!
1%
#216980000000
0!
0%
#216985000000
1!
1%
#216990000000
0!
0%
#216995000000
1!
1%
#217000000000
0!
0%
#217005000000
1!
1%
#217010000000
0!
0%
#217015000000
1!
1%
#217020000000
0!
0%
#217025000000
1!
1%
#217030000000
0!
0%
#217035000000
1!
1%
#217040000000
0!
0%
#217045000000
1!
1%
#217050000000
0!
0%
#217055000000
1!
1%
#217060000000
0!
0%
#217065000000
1!
1%
#217070000000
0!
0%
#217075000000
1!
1%
#217080000000
0!
0%
#217085000000
1!
1%
#217090000000
0!
0%
#217095000000
1!
1%
#217100000000
0!
0%
#217105000000
1!
1%
#217110000000
0!
0%
#217115000000
1!
1%
#217120000000
0!
0%
#217125000000
1!
1%
#217130000000
0!
0%
#217135000000
1!
1%
#217140000000
0!
0%
#217145000000
1!
1%
#217150000000
0!
0%
#217155000000
1!
1%
#217160000000
0!
0%
#217165000000
1!
1%
#217170000000
0!
0%
#217175000000
1!
1%
#217180000000
0!
0%
#217185000000
1!
1%
#217190000000
0!
0%
#217195000000
1!
1%
#217200000000
0!
0%
#217205000000
1!
1%
#217210000000
0!
0%
#217215000000
1!
1%
#217220000000
0!
0%
#217225000000
1!
1%
#217230000000
0!
0%
#217235000000
1!
1%
#217240000000
0!
0%
#217245000000
1!
1%
#217250000000
0!
0%
#217255000000
1!
1%
#217260000000
0!
0%
#217265000000
1!
1%
#217270000000
0!
0%
#217275000000
1!
1%
#217280000000
0!
0%
#217285000000
1!
1%
#217290000000
0!
0%
#217295000000
1!
1%
#217300000000
0!
0%
#217305000000
1!
1%
#217310000000
0!
0%
#217315000000
1!
1%
#217320000000
0!
0%
#217325000000
1!
1%
#217330000000
0!
0%
#217335000000
1!
1%
#217340000000
0!
0%
#217345000000
1!
1%
#217350000000
0!
0%
#217355000000
1!
1%
#217360000000
0!
0%
#217365000000
1!
1%
#217370000000
0!
0%
#217375000000
1!
1%
#217380000000
0!
0%
#217385000000
1!
1%
#217390000000
0!
0%
#217395000000
1!
1%
#217400000000
0!
0%
#217405000000
1!
1%
#217410000000
0!
0%
#217415000000
1!
1%
#217420000000
0!
0%
#217425000000
1!
1%
#217430000000
0!
0%
#217435000000
1!
1%
#217440000000
0!
0%
#217445000000
1!
1%
#217450000000
0!
0%
#217455000000
1!
1%
#217460000000
0!
0%
#217465000000
1!
1%
#217470000000
0!
0%
#217475000000
1!
1%
#217480000000
0!
0%
#217485000000
1!
1%
#217490000000
0!
0%
#217495000000
1!
1%
#217500000000
0!
0%
#217505000000
1!
1%
#217510000000
0!
0%
#217515000000
1!
1%
#217520000000
0!
0%
#217525000000
1!
1%
#217530000000
0!
0%
#217535000000
1!
1%
#217540000000
0!
0%
#217545000000
1!
1%
#217550000000
0!
0%
#217555000000
1!
1%
#217560000000
0!
0%
#217565000000
1!
1%
#217570000000
0!
0%
#217575000000
1!
1%
#217580000000
0!
0%
#217585000000
1!
1%
#217590000000
0!
0%
#217595000000
1!
1%
#217600000000
0!
0%
#217605000000
1!
1%
#217610000000
0!
0%
#217615000000
1!
1%
#217620000000
0!
0%
#217625000000
1!
1%
#217630000000
0!
0%
#217635000000
1!
1%
#217640000000
0!
0%
#217645000000
1!
1%
#217650000000
0!
0%
#217655000000
1!
1%
#217660000000
0!
0%
#217665000000
1!
1%
#217670000000
0!
0%
#217675000000
1!
1%
#217680000000
0!
0%
#217685000000
1!
1%
#217690000000
0!
0%
#217695000000
1!
1%
#217700000000
0!
0%
#217705000000
1!
1%
#217710000000
0!
0%
#217715000000
1!
1%
#217720000000
0!
0%
#217725000000
1!
1%
#217730000000
0!
0%
#217735000000
1!
1%
#217740000000
0!
0%
#217745000000
1!
1%
#217750000000
0!
0%
#217755000000
1!
1%
#217760000000
0!
0%
#217765000000
1!
1%
#217770000000
0!
0%
#217775000000
1!
1%
#217780000000
0!
0%
#217785000000
1!
1%
#217790000000
0!
0%
#217795000000
1!
1%
#217800000000
0!
0%
#217805000000
1!
1%
#217810000000
0!
0%
#217815000000
1!
1%
#217820000000
0!
0%
#217825000000
1!
1%
#217830000000
0!
0%
#217835000000
1!
1%
#217840000000
0!
0%
#217845000000
1!
1%
#217850000000
0!
0%
#217855000000
1!
1%
#217860000000
0!
0%
#217865000000
1!
1%
#217870000000
0!
0%
#217875000000
1!
1%
#217880000000
0!
0%
#217885000000
1!
1%
#217890000000
0!
0%
#217895000000
1!
1%
#217900000000
0!
0%
#217905000000
1!
1%
#217910000000
0!
0%
#217915000000
1!
1%
#217920000000
0!
0%
#217925000000
1!
1%
#217930000000
0!
0%
#217935000000
1!
1%
#217940000000
0!
0%
#217945000000
1!
1%
#217950000000
0!
0%
#217955000000
1!
1%
#217960000000
0!
0%
#217965000000
1!
1%
#217970000000
0!
0%
#217975000000
1!
1%
#217980000000
0!
0%
#217985000000
1!
1%
#217990000000
0!
0%
#217995000000
1!
1%
#218000000000
0!
0%
#218005000000
1!
1%
#218010000000
0!
0%
#218015000000
1!
1%
#218020000000
0!
0%
#218025000000
1!
1%
#218030000000
0!
0%
#218035000000
1!
1%
#218040000000
0!
0%
#218045000000
1!
1%
#218050000000
0!
0%
#218055000000
1!
1%
#218060000000
0!
0%
#218065000000
1!
1%
#218070000000
0!
0%
#218075000000
1!
1%
#218080000000
0!
0%
#218085000000
1!
1%
#218090000000
0!
0%
#218095000000
1!
1%
#218100000000
0!
0%
#218105000000
1!
1%
#218110000000
0!
0%
#218115000000
1!
1%
#218120000000
0!
0%
#218125000000
1!
1%
#218130000000
0!
0%
#218135000000
1!
1%
#218140000000
0!
0%
#218145000000
1!
1%
#218150000000
0!
0%
#218155000000
1!
1%
#218160000000
0!
0%
#218165000000
1!
1%
#218170000000
0!
0%
#218175000000
1!
1%
#218180000000
0!
0%
#218185000000
1!
1%
#218190000000
0!
0%
#218195000000
1!
1%
#218200000000
0!
0%
#218205000000
1!
1%
#218210000000
0!
0%
#218215000000
1!
1%
#218220000000
0!
0%
#218225000000
1!
1%
#218230000000
0!
0%
#218235000000
1!
1%
#218240000000
0!
0%
#218245000000
1!
1%
#218250000000
0!
0%
#218255000000
1!
1%
#218260000000
0!
0%
#218265000000
1!
1%
#218270000000
0!
0%
#218275000000
1!
1%
#218280000000
0!
0%
#218285000000
1!
1%
#218290000000
0!
0%
#218295000000
1!
1%
#218300000000
0!
0%
#218305000000
1!
1%
#218310000000
0!
0%
#218315000000
1!
1%
#218320000000
0!
0%
#218325000000
1!
1%
#218330000000
0!
0%
#218335000000
1!
1%
#218340000000
0!
0%
#218345000000
1!
1%
#218350000000
0!
0%
#218355000000
1!
1%
#218360000000
0!
0%
#218365000000
1!
1%
#218370000000
0!
0%
#218375000000
1!
1%
#218380000000
0!
0%
#218385000000
1!
1%
#218390000000
0!
0%
#218395000000
1!
1%
#218400000000
0!
0%
#218405000000
1!
1%
#218410000000
0!
0%
#218415000000
1!
1%
#218420000000
0!
0%
#218425000000
1!
1%
#218430000000
0!
0%
#218435000000
1!
1%
#218440000000
0!
0%
#218445000000
1!
1%
#218450000000
0!
0%
#218455000000
1!
1%
#218460000000
0!
0%
#218465000000
1!
1%
#218470000000
0!
0%
#218475000000
1!
1%
#218480000000
0!
0%
#218485000000
1!
1%
#218490000000
0!
0%
#218495000000
1!
1%
#218500000000
0!
0%
#218505000000
1!
1%
#218510000000
0!
0%
#218515000000
1!
1%
#218520000000
0!
0%
#218525000000
1!
1%
#218530000000
0!
0%
#218535000000
1!
1%
#218540000000
0!
0%
#218545000000
1!
1%
#218550000000
0!
0%
#218555000000
1!
1%
#218560000000
0!
0%
#218565000000
1!
1%
#218570000000
0!
0%
#218575000000
1!
1%
#218580000000
0!
0%
#218585000000
1!
1%
#218590000000
0!
0%
#218595000000
1!
1%
#218600000000
0!
0%
#218605000000
1!
1%
#218610000000
0!
0%
#218615000000
1!
1%
#218620000000
0!
0%
#218625000000
1!
1%
#218630000000
0!
0%
#218635000000
1!
1%
#218640000000
0!
0%
#218645000000
1!
1%
#218650000000
0!
0%
#218655000000
1!
1%
#218660000000
0!
0%
#218665000000
1!
1%
#218670000000
0!
0%
#218675000000
1!
1%
#218680000000
0!
0%
#218685000000
1!
1%
#218690000000
0!
0%
#218695000000
1!
1%
#218700000000
0!
0%
#218705000000
1!
1%
#218710000000
0!
0%
#218715000000
1!
1%
#218720000000
0!
0%
#218725000000
1!
1%
#218730000000
0!
0%
#218735000000
1!
1%
#218740000000
0!
0%
#218745000000
1!
1%
#218750000000
0!
0%
#218755000000
1!
1%
#218760000000
0!
0%
#218765000000
1!
1%
#218770000000
0!
0%
#218775000000
1!
1%
#218780000000
0!
0%
#218785000000
1!
1%
#218790000000
0!
0%
#218795000000
1!
1%
#218800000000
0!
0%
#218805000000
1!
1%
#218810000000
0!
0%
#218815000000
1!
1%
#218820000000
0!
0%
#218825000000
1!
1%
#218830000000
0!
0%
#218835000000
1!
1%
#218840000000
0!
0%
#218845000000
1!
1%
#218850000000
0!
0%
#218855000000
1!
1%
#218860000000
0!
0%
#218865000000
1!
1%
#218870000000
0!
0%
#218875000000
1!
1%
#218880000000
0!
0%
#218885000000
1!
1%
#218890000000
0!
0%
#218895000000
1!
1%
#218900000000
0!
0%
#218905000000
1!
1%
#218910000000
0!
0%
#218915000000
1!
1%
#218920000000
0!
0%
#218925000000
1!
1%
#218930000000
0!
0%
#218935000000
1!
1%
#218940000000
0!
0%
#218945000000
1!
1%
#218950000000
0!
0%
#218955000000
1!
1%
#218960000000
0!
0%
#218965000000
1!
1%
#218970000000
0!
0%
#218975000000
1!
1%
#218980000000
0!
0%
#218985000000
1!
1%
#218990000000
0!
0%
#218995000000
1!
1%
#219000000000
0!
0%
#219005000000
1!
1%
#219010000000
0!
0%
#219015000000
1!
1%
#219020000000
0!
0%
#219025000000
1!
1%
#219030000000
0!
0%
#219035000000
1!
1%
#219040000000
0!
0%
#219045000000
1!
1%
#219050000000
0!
0%
#219055000000
1!
1%
#219060000000
0!
0%
#219065000000
1!
1%
#219070000000
0!
0%
#219075000000
1!
1%
#219080000000
0!
0%
#219085000000
1!
1%
#219090000000
0!
0%
#219095000000
1!
1%
#219100000000
0!
0%
#219105000000
1!
1%
#219110000000
0!
0%
#219115000000
1!
1%
#219120000000
0!
0%
#219125000000
1!
1%
#219130000000
0!
0%
#219135000000
1!
1%
#219140000000
0!
0%
#219145000000
1!
1%
#219150000000
0!
0%
#219155000000
1!
1%
#219160000000
0!
0%
#219165000000
1!
1%
#219170000000
0!
0%
#219175000000
1!
1%
#219180000000
0!
0%
#219185000000
1!
1%
#219190000000
0!
0%
#219195000000
1!
1%
#219200000000
0!
0%
#219205000000
1!
1%
#219210000000
0!
0%
#219215000000
1!
1%
#219220000000
0!
0%
#219225000000
1!
1%
#219230000000
0!
0%
#219235000000
1!
1%
#219240000000
0!
0%
#219245000000
1!
1%
#219250000000
0!
0%
#219255000000
1!
1%
#219260000000
0!
0%
#219265000000
1!
1%
#219270000000
0!
0%
#219275000000
1!
1%
#219280000000
0!
0%
#219285000000
1!
1%
#219290000000
0!
0%
#219295000000
1!
1%
#219300000000
0!
0%
#219305000000
1!
1%
#219310000000
0!
0%
#219315000000
1!
1%
#219320000000
0!
0%
#219325000000
1!
1%
#219330000000
0!
0%
#219335000000
1!
1%
#219340000000
0!
0%
#219345000000
1!
1%
#219350000000
0!
0%
#219355000000
1!
1%
#219360000000
0!
0%
#219365000000
1!
1%
#219370000000
0!
0%
#219375000000
1!
1%
#219380000000
0!
0%
#219385000000
1!
1%
#219390000000
0!
0%
#219395000000
1!
1%
#219400000000
0!
0%
#219405000000
1!
1%
#219410000000
0!
0%
#219415000000
1!
1%
#219420000000
0!
0%
#219425000000
1!
1%
#219430000000
0!
0%
#219435000000
1!
1%
#219440000000
0!
0%
#219445000000
1!
1%
#219450000000
0!
0%
#219455000000
1!
1%
#219460000000
0!
0%
#219465000000
1!
1%
#219470000000
0!
0%
#219475000000
1!
1%
#219480000000
0!
0%
#219485000000
1!
1%
#219490000000
0!
0%
#219495000000
1!
1%
#219500000000
0!
0%
#219505000000
1!
1%
#219510000000
0!
0%
#219515000000
1!
1%
#219520000000
0!
0%
#219525000000
1!
1%
#219530000000
0!
0%
#219535000000
1!
1%
#219540000000
0!
0%
#219545000000
1!
1%
#219550000000
0!
0%
#219555000000
1!
1%
#219560000000
0!
0%
#219565000000
1!
1%
#219570000000
0!
0%
#219575000000
1!
1%
#219580000000
0!
0%
#219585000000
1!
1%
#219590000000
0!
0%
#219595000000
1!
1%
#219600000000
0!
0%
#219605000000
1!
1%
#219610000000
0!
0%
#219615000000
1!
1%
#219620000000
0!
0%
#219625000000
1!
1%
#219630000000
0!
0%
#219635000000
1!
1%
#219640000000
0!
0%
#219645000000
1!
1%
#219650000000
0!
0%
#219655000000
1!
1%
#219660000000
0!
0%
#219665000000
1!
1%
#219670000000
0!
0%
#219675000000
1!
1%
#219680000000
0!
0%
#219685000000
1!
1%
#219690000000
0!
0%
#219695000000
1!
1%
#219700000000
0!
0%
#219705000000
1!
1%
#219710000000
0!
0%
#219715000000
1!
1%
#219720000000
0!
0%
#219725000000
1!
1%
#219730000000
0!
0%
#219735000000
1!
1%
#219740000000
0!
0%
#219745000000
1!
1%
#219750000000
0!
0%
#219755000000
1!
1%
#219760000000
0!
0%
#219765000000
1!
1%
#219770000000
0!
0%
#219775000000
1!
1%
#219780000000
0!
0%
#219785000000
1!
1%
#219790000000
0!
0%
#219795000000
1!
1%
#219800000000
0!
0%
#219805000000
1!
1%
#219810000000
0!
0%
#219815000000
1!
1%
#219820000000
0!
0%
#219825000000
1!
1%
#219830000000
0!
0%
#219835000000
1!
1%
#219840000000
0!
0%
#219845000000
1!
1%
#219850000000
0!
0%
#219855000000
1!
1%
#219860000000
0!
0%
#219865000000
1!
1%
#219870000000
0!
0%
#219875000000
1!
1%
#219880000000
0!
0%
#219885000000
1!
1%
#219890000000
0!
0%
#219895000000
1!
1%
#219900000000
0!
0%
#219905000000
1!
1%
#219910000000
0!
0%
#219915000000
1!
1%
#219920000000
0!
0%
#219925000000
1!
1%
#219930000000
0!
0%
#219935000000
1!
1%
#219940000000
0!
0%
#219945000000
1!
1%
#219950000000
0!
0%
#219955000000
1!
1%
#219960000000
0!
0%
#219965000000
1!
1%
#219970000000
0!
0%
#219975000000
1!
1%
#219980000000
0!
0%
#219985000000
1!
1%
#219990000000
0!
0%
#219995000000
1!
1%
#220000000000
0!
0%
#220005000000
1!
1%
#220010000000
0!
0%
#220015000000
1!
1%
#220020000000
0!
0%
#220025000000
1!
1%
#220030000000
0!
0%
#220035000000
1!
1%
#220040000000
0!
0%
#220045000000
1!
1%
#220050000000
0!
0%
#220055000000
1!
1%
#220060000000
0!
0%
#220065000000
1!
1%
#220070000000
0!
0%
#220075000000
1!
1%
#220080000000
0!
0%
#220085000000
1!
1%
#220090000000
0!
0%
#220095000000
1!
1%
#220100000000
0!
0%
#220105000000
1!
1%
#220110000000
0!
0%
#220115000000
1!
1%
#220120000000
0!
0%
#220125000000
1!
1%
#220130000000
0!
0%
#220135000000
1!
1%
#220140000000
0!
0%
#220145000000
1!
1%
#220150000000
0!
0%
#220155000000
1!
1%
#220160000000
0!
0%
#220165000000
1!
1%
#220170000000
0!
0%
#220175000000
1!
1%
#220180000000
0!
0%
#220185000000
1!
1%
#220190000000
0!
0%
#220195000000
1!
1%
#220200000000
0!
0%
#220205000000
1!
1%
#220210000000
0!
0%
#220215000000
1!
1%
#220220000000
0!
0%
#220225000000
1!
1%
#220230000000
0!
0%
#220235000000
1!
1%
#220240000000
0!
0%
#220245000000
1!
1%
#220250000000
0!
0%
#220255000000
1!
1%
#220260000000
0!
0%
#220265000000
1!
1%
#220270000000
0!
0%
#220275000000
1!
1%
#220280000000
0!
0%
#220285000000
1!
1%
#220290000000
0!
0%
#220295000000
1!
1%
#220300000000
0!
0%
#220305000000
1!
1%
#220310000000
0!
0%
#220315000000
1!
1%
#220320000000
0!
0%
#220325000000
1!
1%
#220330000000
0!
0%
#220335000000
1!
1%
#220340000000
0!
0%
#220345000000
1!
1%
#220350000000
0!
0%
#220355000000
1!
1%
#220360000000
0!
0%
#220365000000
1!
1%
#220370000000
0!
0%
#220375000000
1!
1%
#220380000000
0!
0%
#220385000000
1!
1%
#220390000000
0!
0%
#220395000000
1!
1%
#220400000000
0!
0%
#220405000000
1!
1%
#220410000000
0!
0%
#220415000000
1!
1%
#220420000000
0!
0%
#220425000000
1!
1%
#220430000000
0!
0%
#220435000000
1!
1%
#220440000000
0!
0%
#220445000000
1!
1%
#220450000000
0!
0%
#220455000000
1!
1%
#220460000000
0!
0%
#220465000000
1!
1%
#220470000000
0!
0%
#220475000000
1!
1%
#220480000000
0!
0%
#220485000000
1!
1%
#220490000000
0!
0%
#220495000000
1!
1%
#220500000000
0!
0%
#220505000000
1!
1%
#220510000000
0!
0%
#220515000000
1!
1%
#220520000000
0!
0%
#220525000000
1!
1%
#220530000000
0!
0%
#220535000000
1!
1%
#220540000000
0!
0%
#220545000000
1!
1%
#220550000000
0!
0%
#220555000000
1!
1%
#220560000000
0!
0%
#220565000000
1!
1%
#220570000000
0!
0%
#220575000000
1!
1%
#220580000000
0!
0%
#220585000000
1!
1%
#220590000000
0!
0%
#220595000000
1!
1%
#220600000000
0!
0%
#220605000000
1!
1%
#220610000000
0!
0%
#220615000000
1!
1%
#220620000000
0!
0%
#220625000000
1!
1%
#220630000000
0!
0%
#220635000000
1!
1%
#220640000000
0!
0%
#220645000000
1!
1%
#220650000000
0!
0%
#220655000000
1!
1%
#220660000000
0!
0%
#220665000000
1!
1%
#220670000000
0!
0%
#220675000000
1!
1%
#220680000000
0!
0%
#220685000000
1!
1%
#220690000000
0!
0%
#220695000000
1!
1%
#220700000000
0!
0%
#220705000000
1!
1%
#220710000000
0!
0%
#220715000000
1!
1%
#220720000000
0!
0%
#220725000000
1!
1%
#220730000000
0!
0%
#220735000000
1!
1%
#220740000000
0!
0%
#220745000000
1!
1%
#220750000000
0!
0%
#220755000000
1!
1%
#220760000000
0!
0%
#220765000000
1!
1%
#220770000000
0!
0%
#220775000000
1!
1%
#220780000000
0!
0%
#220785000000
1!
1%
#220790000000
0!
0%
#220795000000
1!
1%
#220800000000
0!
0%
#220805000000
1!
1%
#220810000000
0!
0%
#220815000000
1!
1%
#220820000000
0!
0%
#220825000000
1!
1%
#220830000000
0!
0%
#220835000000
1!
1%
#220840000000
0!
0%
#220845000000
1!
1%
#220850000000
0!
0%
#220855000000
1!
1%
#220860000000
0!
0%
#220865000000
1!
1%
#220870000000
0!
0%
#220875000000
1!
1%
#220880000000
0!
0%
#220885000000
1!
1%
#220890000000
0!
0%
#220895000000
1!
1%
#220900000000
0!
0%
#220905000000
1!
1%
#220910000000
0!
0%
#220915000000
1!
1%
#220920000000
0!
0%
#220925000000
1!
1%
#220930000000
0!
0%
#220935000000
1!
1%
#220940000000
0!
0%
#220945000000
1!
1%
#220950000000
0!
0%
#220955000000
1!
1%
#220960000000
0!
0%
#220965000000
1!
1%
#220970000000
0!
0%
#220975000000
1!
1%
#220980000000
0!
0%
#220985000000
1!
1%
#220990000000
0!
0%
#220995000000
1!
1%
#221000000000
0!
0%
#221005000000
1!
1%
#221010000000
0!
0%
#221015000000
1!
1%
#221020000000
0!
0%
#221025000000
1!
1%
#221030000000
0!
0%
#221035000000
1!
1%
#221040000000
0!
0%
#221045000000
1!
1%
#221050000000
0!
0%
#221055000000
1!
1%
#221060000000
0!
0%
#221065000000
1!
1%
#221070000000
0!
0%
#221075000000
1!
1%
#221080000000
0!
0%
#221085000000
1!
1%
#221090000000
0!
0%
#221095000000
1!
1%
#221100000000
0!
0%
#221105000000
1!
1%
#221110000000
0!
0%
#221115000000
1!
1%
#221120000000
0!
0%
#221125000000
1!
1%
#221130000000
0!
0%
#221135000000
1!
1%
#221140000000
0!
0%
#221145000000
1!
1%
#221150000000
0!
0%
#221155000000
1!
1%
#221160000000
0!
0%
#221165000000
1!
1%
#221170000000
0!
0%
#221175000000
1!
1%
#221180000000
0!
0%
#221185000000
1!
1%
#221190000000
0!
0%
#221195000000
1!
1%
#221200000000
0!
0%
#221205000000
1!
1%
#221210000000
0!
0%
#221215000000
1!
1%
#221220000000
0!
0%
#221225000000
1!
1%
#221230000000
0!
0%
#221235000000
1!
1%
#221240000000
0!
0%
#221245000000
1!
1%
#221250000000
0!
0%
#221255000000
1!
1%
#221260000000
0!
0%
#221265000000
1!
1%
#221270000000
0!
0%
#221275000000
1!
1%
#221280000000
0!
0%
#221285000000
1!
1%
#221290000000
0!
0%
#221295000000
1!
1%
#221300000000
0!
0%
#221305000000
1!
1%
#221310000000
0!
0%
#221315000000
1!
1%
#221320000000
0!
0%
#221325000000
1!
1%
#221330000000
0!
0%
#221335000000
1!
1%
#221340000000
0!
0%
#221345000000
1!
1%
#221350000000
0!
0%
#221355000000
1!
1%
#221360000000
0!
0%
#221365000000
1!
1%
#221370000000
0!
0%
#221375000000
1!
1%
#221380000000
0!
0%
#221385000000
1!
1%
#221390000000
0!
0%
#221395000000
1!
1%
#221400000000
0!
0%
#221405000000
1!
1%
#221410000000
0!
0%
#221415000000
1!
1%
#221420000000
0!
0%
#221425000000
1!
1%
#221430000000
0!
0%
#221435000000
1!
1%
#221440000000
0!
0%
#221445000000
1!
1%
#221450000000
0!
0%
#221455000000
1!
1%
#221460000000
0!
0%
#221465000000
1!
1%
#221470000000
0!
0%
#221475000000
1!
1%
#221480000000
0!
0%
#221485000000
1!
1%
#221490000000
0!
0%
#221495000000
1!
1%
#221500000000
0!
0%
#221505000000
1!
1%
#221510000000
0!
0%
#221515000000
1!
1%
#221520000000
0!
0%
#221525000000
1!
1%
#221530000000
0!
0%
#221535000000
1!
1%
#221540000000
0!
0%
#221545000000
1!
1%
#221550000000
0!
0%
#221555000000
1!
1%
#221560000000
0!
0%
#221565000000
1!
1%
#221570000000
0!
0%
#221575000000
1!
1%
#221580000000
0!
0%
#221585000000
1!
1%
#221590000000
0!
0%
#221595000000
1!
1%
#221600000000
0!
0%
#221605000000
1!
1%
#221610000000
0!
0%
#221615000000
1!
1%
#221620000000
0!
0%
#221625000000
1!
1%
#221630000000
0!
0%
#221635000000
1!
1%
#221640000000
0!
0%
#221645000000
1!
1%
#221650000000
0!
0%
#221655000000
1!
1%
#221660000000
0!
0%
#221665000000
1!
1%
#221670000000
0!
0%
#221675000000
1!
1%
#221680000000
0!
0%
#221685000000
1!
1%
#221690000000
0!
0%
#221695000000
1!
1%
#221700000000
0!
0%
#221705000000
1!
1%
#221710000000
0!
0%
#221715000000
1!
1%
#221720000000
0!
0%
#221725000000
1!
1%
#221730000000
0!
0%
#221735000000
1!
1%
#221740000000
0!
0%
#221745000000
1!
1%
#221750000000
0!
0%
#221755000000
1!
1%
#221760000000
0!
0%
#221765000000
1!
1%
#221770000000
0!
0%
#221775000000
1!
1%
#221780000000
0!
0%
#221785000000
1!
1%
#221790000000
0!
0%
#221795000000
1!
1%
#221800000000
0!
0%
#221805000000
1!
1%
#221810000000
0!
0%
#221815000000
1!
1%
#221820000000
0!
0%
#221825000000
1!
1%
#221830000000
0!
0%
#221835000000
1!
1%
#221840000000
0!
0%
#221845000000
1!
1%
#221850000000
0!
0%
#221855000000
1!
1%
#221860000000
0!
0%
#221865000000
1!
1%
#221870000000
0!
0%
#221875000000
1!
1%
#221880000000
0!
0%
#221885000000
1!
1%
#221890000000
0!
0%
#221895000000
1!
1%
#221900000000
0!
0%
#221905000000
1!
1%
#221910000000
0!
0%
#221915000000
1!
1%
#221920000000
0!
0%
#221925000000
1!
1%
#221930000000
0!
0%
#221935000000
1!
1%
#221940000000
0!
0%
#221945000000
1!
1%
#221950000000
0!
0%
#221955000000
1!
1%
#221960000000
0!
0%
#221965000000
1!
1%
#221970000000
0!
0%
#221975000000
1!
1%
#221980000000
0!
0%
#221985000000
1!
1%
#221990000000
0!
0%
#221995000000
1!
1%
#222000000000
0!
0%
#222005000000
1!
1%
#222010000000
0!
0%
#222015000000
1!
1%
#222020000000
0!
0%
#222025000000
1!
1%
#222030000000
0!
0%
#222035000000
1!
1%
#222040000000
0!
0%
#222045000000
1!
1%
#222050000000
0!
0%
#222055000000
1!
1%
#222060000000
0!
0%
#222065000000
1!
1%
#222070000000
0!
0%
#222075000000
1!
1%
#222080000000
0!
0%
#222085000000
1!
1%
#222090000000
0!
0%
#222095000000
1!
1%
#222100000000
0!
0%
#222105000000
1!
1%
#222110000000
0!
0%
#222115000000
1!
1%
#222120000000
0!
0%
#222125000000
1!
1%
#222130000000
0!
0%
#222135000000
1!
1%
#222140000000
0!
0%
#222145000000
1!
1%
#222150000000
0!
0%
#222155000000
1!
1%
#222160000000
0!
0%
#222165000000
1!
1%
#222170000000
0!
0%
#222175000000
1!
1%
#222180000000
0!
0%
#222185000000
1!
1%
#222190000000
0!
0%
#222195000000
1!
1%
#222200000000
0!
0%
#222205000000
1!
1%
#222210000000
0!
0%
#222215000000
1!
1%
#222220000000
0!
0%
#222225000000
1!
1%
#222230000000
0!
0%
#222235000000
1!
1%
#222240000000
0!
0%
#222245000000
1!
1%
#222250000000
0!
0%
#222255000000
1!
1%
#222260000000
0!
0%
#222265000000
1!
1%
#222270000000
0!
0%
#222275000000
1!
1%
#222280000000
0!
0%
#222285000000
1!
1%
#222290000000
0!
0%
#222295000000
1!
1%
#222300000000
0!
0%
#222305000000
1!
1%
#222310000000
0!
0%
#222315000000
1!
1%
#222320000000
0!
0%
#222325000000
1!
1%
#222330000000
0!
0%
#222335000000
1!
1%
#222340000000
0!
0%
#222345000000
1!
1%
#222350000000
0!
0%
#222355000000
1!
1%
#222360000000
0!
0%
#222365000000
1!
1%
#222370000000
0!
0%
#222375000000
1!
1%
#222380000000
0!
0%
#222385000000
1!
1%
#222390000000
0!
0%
#222395000000
1!
1%
#222400000000
0!
0%
#222405000000
1!
1%
#222410000000
0!
0%
#222415000000
1!
1%
#222420000000
0!
0%
#222425000000
1!
1%
#222430000000
0!
0%
#222435000000
1!
1%
#222440000000
0!
0%
#222445000000
1!
1%
#222450000000
0!
0%
#222455000000
1!
1%
#222460000000
0!
0%
#222465000000
1!
1%
#222470000000
0!
0%
#222475000000
1!
1%
#222480000000
0!
0%
#222485000000
1!
1%
#222490000000
0!
0%
#222495000000
1!
1%
#222500000000
0!
0%
#222505000000
1!
1%
#222510000000
0!
0%
#222515000000
1!
1%
#222520000000
0!
0%
#222525000000
1!
1%
#222530000000
0!
0%
#222535000000
1!
1%
#222540000000
0!
0%
#222545000000
1!
1%
#222550000000
0!
0%
#222555000000
1!
1%
#222560000000
0!
0%
#222565000000
1!
1%
#222570000000
0!
0%
#222575000000
1!
1%
#222580000000
0!
0%
#222585000000
1!
1%
#222590000000
0!
0%
#222595000000
1!
1%
#222600000000
0!
0%
#222605000000
1!
1%
#222610000000
0!
0%
#222615000000
1!
1%
#222620000000
0!
0%
#222625000000
1!
1%
#222630000000
0!
0%
#222635000000
1!
1%
#222640000000
0!
0%
#222645000000
1!
1%
#222650000000
0!
0%
#222655000000
1!
1%
#222660000000
0!
0%
#222665000000
1!
1%
#222670000000
0!
0%
#222675000000
1!
1%
#222680000000
0!
0%
#222685000000
1!
1%
#222690000000
0!
0%
#222695000000
1!
1%
#222700000000
0!
0%
#222705000000
1!
1%
#222710000000
0!
0%
#222715000000
1!
1%
#222720000000
0!
0%
#222725000000
1!
1%
#222730000000
0!
0%
#222735000000
1!
1%
#222740000000
0!
0%
#222745000000
1!
1%
#222750000000
0!
0%
#222755000000
1!
1%
#222760000000
0!
0%
#222765000000
1!
1%
#222770000000
0!
0%
#222775000000
1!
1%
#222780000000
0!
0%
#222785000000
1!
1%
#222790000000
0!
0%
#222795000000
1!
1%
#222800000000
0!
0%
#222805000000
1!
1%
#222810000000
0!
0%
#222815000000
1!
1%
#222820000000
0!
0%
#222825000000
1!
1%
#222830000000
0!
0%
#222835000000
1!
1%
#222840000000
0!
0%
#222845000000
1!
1%
#222850000000
0!
0%
#222855000000
1!
1%
#222860000000
0!
0%
#222865000000
1!
1%
#222870000000
0!
0%
#222875000000
1!
1%
#222880000000
0!
0%
#222885000000
1!
1%
#222890000000
0!
0%
#222895000000
1!
1%
#222900000000
0!
0%
#222905000000
1!
1%
#222910000000
0!
0%
#222915000000
1!
1%
#222920000000
0!
0%
#222925000000
1!
1%
#222930000000
0!
0%
#222935000000
1!
1%
#222940000000
0!
0%
#222945000000
1!
1%
#222950000000
0!
0%
#222955000000
1!
1%
#222960000000
0!
0%
#222965000000
1!
1%
#222970000000
0!
0%
#222975000000
1!
1%
#222980000000
0!
0%
#222985000000
1!
1%
#222990000000
0!
0%
#222995000000
1!
1%
#223000000000
0!
0%
#223005000000
1!
1%
#223010000000
0!
0%
#223015000000
1!
1%
#223020000000
0!
0%
#223025000000
1!
1%
#223030000000
0!
0%
#223035000000
1!
1%
#223040000000
0!
0%
#223045000000
1!
1%
#223050000000
0!
0%
#223055000000
1!
1%
#223060000000
0!
0%
#223065000000
1!
1%
#223070000000
0!
0%
#223075000000
1!
1%
#223080000000
0!
0%
#223085000000
1!
1%
#223090000000
0!
0%
#223095000000
1!
1%
#223100000000
0!
0%
#223105000000
1!
1%
#223110000000
0!
0%
#223115000000
1!
1%
#223120000000
0!
0%
#223125000000
1!
1%
#223130000000
0!
0%
#223135000000
1!
1%
#223140000000
0!
0%
#223145000000
1!
1%
#223150000000
0!
0%
#223155000000
1!
1%
#223160000000
0!
0%
#223165000000
1!
1%
#223170000000
0!
0%
#223175000000
1!
1%
#223180000000
0!
0%
#223185000000
1!
1%
#223190000000
0!
0%
#223195000000
1!
1%
#223200000000
0!
0%
#223205000000
1!
1%
#223210000000
0!
0%
#223215000000
1!
1%
#223220000000
0!
0%
#223225000000
1!
1%
#223230000000
0!
0%
#223235000000
1!
1%
#223240000000
0!
0%
#223245000000
1!
1%
#223250000000
0!
0%
#223255000000
1!
1%
#223260000000
0!
0%
#223265000000
1!
1%
#223270000000
0!
0%
#223275000000
1!
1%
#223280000000
0!
0%
#223285000000
1!
1%
#223290000000
0!
0%
#223295000000
1!
1%
#223300000000
0!
0%
#223305000000
1!
1%
#223310000000
0!
0%
#223315000000
1!
1%
#223320000000
0!
0%
#223325000000
1!
1%
#223330000000
0!
0%
#223335000000
1!
1%
#223340000000
0!
0%
#223345000000
1!
1%
#223350000000
0!
0%
#223355000000
1!
1%
#223360000000
0!
0%
#223365000000
1!
1%
#223370000000
0!
0%
#223375000000
1!
1%
#223380000000
0!
0%
#223385000000
1!
1%
#223390000000
0!
0%
#223395000000
1!
1%
#223400000000
0!
0%
#223405000000
1!
1%
#223410000000
0!
0%
#223415000000
1!
1%
#223420000000
0!
0%
#223425000000
1!
1%
#223430000000
0!
0%
#223435000000
1!
1%
#223440000000
0!
0%
#223445000000
1!
1%
#223450000000
0!
0%
#223455000000
1!
1%
#223460000000
0!
0%
#223465000000
1!
1%
#223470000000
0!
0%
#223475000000
1!
1%
#223480000000
0!
0%
#223485000000
1!
1%
#223490000000
0!
0%
#223495000000
1!
1%
#223500000000
0!
0%
#223505000000
1!
1%
#223510000000
0!
0%
#223515000000
1!
1%
#223520000000
0!
0%
#223525000000
1!
1%
#223530000000
0!
0%
#223535000000
1!
1%
#223540000000
0!
0%
#223545000000
1!
1%
#223550000000
0!
0%
#223555000000
1!
1%
#223560000000
0!
0%
#223565000000
1!
1%
#223570000000
0!
0%
#223575000000
1!
1%
#223580000000
0!
0%
#223585000000
1!
1%
#223590000000
0!
0%
#223595000000
1!
1%
#223600000000
0!
0%
#223605000000
1!
1%
#223610000000
0!
0%
#223615000000
1!
1%
#223620000000
0!
0%
#223625000000
1!
1%
#223630000000
0!
0%
#223635000000
1!
1%
#223640000000
0!
0%
#223645000000
1!
1%
#223650000000
0!
0%
#223655000000
1!
1%
#223660000000
0!
0%
#223665000000
1!
1%
#223670000000
0!
0%
#223675000000
1!
1%
#223680000000
0!
0%
#223685000000
1!
1%
#223690000000
0!
0%
#223695000000
1!
1%
#223700000000
0!
0%
#223705000000
1!
1%
#223710000000
0!
0%
#223715000000
1!
1%
#223720000000
0!
0%
#223725000000
1!
1%
#223730000000
0!
0%
#223735000000
1!
1%
#223740000000
0!
0%
#223745000000
1!
1%
#223750000000
0!
0%
#223755000000
1!
1%
#223760000000
0!
0%
#223765000000
1!
1%
#223770000000
0!
0%
#223775000000
1!
1%
#223780000000
0!
0%
#223785000000
1!
1%
#223790000000
0!
0%
#223795000000
1!
1%
#223800000000
0!
0%
#223805000000
1!
1%
#223810000000
0!
0%
#223815000000
1!
1%
#223820000000
0!
0%
#223825000000
1!
1%
#223830000000
0!
0%
#223835000000
1!
1%
#223840000000
0!
0%
#223845000000
1!
1%
#223850000000
0!
0%
#223855000000
1!
1%
#223860000000
0!
0%
#223865000000
1!
1%
#223870000000
0!
0%
#223875000000
1!
1%
#223880000000
0!
0%
#223885000000
1!
1%
#223890000000
0!
0%
#223895000000
1!
1%
#223900000000
0!
0%
#223905000000
1!
1%
#223910000000
0!
0%
#223915000000
1!
1%
#223920000000
0!
0%
#223925000000
1!
1%
#223930000000
0!
0%
#223935000000
1!
1%
#223940000000
0!
0%
#223945000000
1!
1%
#223950000000
0!
0%
#223955000000
1!
1%
#223960000000
0!
0%
#223965000000
1!
1%
#223970000000
0!
0%
#223975000000
1!
1%
#223980000000
0!
0%
#223985000000
1!
1%
#223990000000
0!
0%
#223995000000
1!
1%
#224000000000
0!
0%
#224005000000
1!
1%
#224010000000
0!
0%
#224015000000
1!
1%
#224020000000
0!
0%
#224025000000
1!
1%
#224030000000
0!
0%
#224035000000
1!
1%
#224040000000
0!
0%
#224045000000
1!
1%
#224050000000
0!
0%
#224055000000
1!
1%
#224060000000
0!
0%
#224065000000
1!
1%
#224070000000
0!
0%
#224075000000
1!
1%
#224080000000
0!
0%
#224085000000
1!
1%
#224090000000
0!
0%
#224095000000
1!
1%
#224100000000
0!
0%
#224105000000
1!
1%
#224110000000
0!
0%
#224115000000
1!
1%
#224120000000
0!
0%
#224125000000
1!
1%
#224130000000
0!
0%
#224135000000
1!
1%
#224140000000
0!
0%
#224145000000
1!
1%
#224150000000
0!
0%
#224155000000
1!
1%
#224160000000
0!
0%
#224165000000
1!
1%
#224170000000
0!
0%
#224175000000
1!
1%
#224180000000
0!
0%
#224185000000
1!
1%
#224190000000
0!
0%
#224195000000
1!
1%
#224200000000
0!
0%
#224205000000
1!
1%
#224210000000
0!
0%
#224215000000
1!
1%
#224220000000
0!
0%
#224225000000
1!
1%
#224230000000
0!
0%
#224235000000
1!
1%
#224240000000
0!
0%
#224245000000
1!
1%
#224250000000
0!
0%
#224255000000
1!
1%
#224260000000
0!
0%
#224265000000
1!
1%
#224270000000
0!
0%
#224275000000
1!
1%
#224280000000
0!
0%
#224285000000
1!
1%
#224290000000
0!
0%
#224295000000
1!
1%
#224300000000
0!
0%
#224305000000
1!
1%
#224310000000
0!
0%
#224315000000
1!
1%
#224320000000
0!
0%
#224325000000
1!
1%
#224330000000
0!
0%
#224335000000
1!
1%
#224340000000
0!
0%
#224345000000
1!
1%
#224350000000
0!
0%
#224355000000
1!
1%
#224360000000
0!
0%
#224365000000
1!
1%
#224370000000
0!
0%
#224375000000
1!
1%
#224380000000
0!
0%
#224385000000
1!
1%
#224390000000
0!
0%
#224395000000
1!
1%
#224400000000
0!
0%
#224405000000
1!
1%
#224410000000
0!
0%
#224415000000
1!
1%
#224420000000
0!
0%
#224425000000
1!
1%
#224430000000
0!
0%
#224435000000
1!
1%
#224440000000
0!
0%
#224445000000
1!
1%
#224450000000
0!
0%
#224455000000
1!
1%
#224460000000
0!
0%
#224465000000
1!
1%
#224470000000
0!
0%
#224475000000
1!
1%
#224480000000
0!
0%
#224485000000
1!
1%
#224490000000
0!
0%
#224495000000
1!
1%
#224500000000
0!
0%
#224505000000
1!
1%
#224510000000
0!
0%
#224515000000
1!
1%
#224520000000
0!
0%
#224525000000
1!
1%
#224530000000
0!
0%
#224535000000
1!
1%
#224540000000
0!
0%
#224545000000
1!
1%
#224550000000
0!
0%
#224555000000
1!
1%
#224560000000
0!
0%
#224565000000
1!
1%
#224570000000
0!
0%
#224575000000
1!
1%
#224580000000
0!
0%
#224585000000
1!
1%
#224590000000
0!
0%
#224595000000
1!
1%
#224600000000
0!
0%
#224605000000
1!
1%
#224610000000
0!
0%
#224615000000
1!
1%
#224620000000
0!
0%
#224625000000
1!
1%
#224630000000
0!
0%
#224635000000
1!
1%
#224640000000
0!
0%
#224645000000
1!
1%
#224650000000
0!
0%
#224655000000
1!
1%
#224660000000
0!
0%
#224665000000
1!
1%
#224670000000
0!
0%
#224675000000
1!
1%
#224680000000
0!
0%
#224685000000
1!
1%
#224690000000
0!
0%
#224695000000
1!
1%
#224700000000
0!
0%
#224705000000
1!
1%
#224710000000
0!
0%
#224715000000
1!
1%
#224720000000
0!
0%
#224725000000
1!
1%
#224730000000
0!
0%
#224735000000
1!
1%
#224740000000
0!
0%
#224745000000
1!
1%
#224750000000
0!
0%
#224755000000
1!
1%
#224760000000
0!
0%
#224765000000
1!
1%
#224770000000
0!
0%
#224775000000
1!
1%
#224780000000
0!
0%
#224785000000
1!
1%
#224790000000
0!
0%
#224795000000
1!
1%
#224800000000
0!
0%
#224805000000
1!
1%
#224810000000
0!
0%
#224815000000
1!
1%
#224820000000
0!
0%
#224825000000
1!
1%
#224830000000
0!
0%
#224835000000
1!
1%
#224840000000
0!
0%
#224845000000
1!
1%
#224850000000
0!
0%
#224855000000
1!
1%
#224860000000
0!
0%
#224865000000
1!
1%
#224870000000
0!
0%
#224875000000
1!
1%
#224880000000
0!
0%
#224885000000
1!
1%
#224890000000
0!
0%
#224895000000
1!
1%
#224900000000
0!
0%
#224905000000
1!
1%
#224910000000
0!
0%
#224915000000
1!
1%
#224920000000
0!
0%
#224925000000
1!
1%
#224930000000
0!
0%
#224935000000
1!
1%
#224940000000
0!
0%
#224945000000
1!
1%
#224950000000
0!
0%
#224955000000
1!
1%
#224960000000
0!
0%
#224965000000
1!
1%
#224970000000
0!
0%
#224975000000
1!
1%
#224980000000
0!
0%
#224985000000
1!
1%
#224990000000
0!
0%
#224995000000
1!
1%
#225000000000
0!
0%
#225005000000
1!
1%
#225010000000
0!
0%
#225015000000
1!
1%
#225020000000
0!
0%
#225025000000
1!
1%
#225030000000
0!
0%
#225035000000
1!
1%
#225040000000
0!
0%
#225045000000
1!
1%
#225050000000
0!
0%
#225055000000
1!
1%
#225060000000
0!
0%
#225065000000
1!
1%
#225070000000
0!
0%
#225075000000
1!
1%
#225080000000
0!
0%
#225085000000
1!
1%
#225090000000
0!
0%
#225095000000
1!
1%
#225100000000
0!
0%
#225105000000
1!
1%
#225110000000
0!
0%
#225115000000
1!
1%
#225120000000
0!
0%
#225125000000
1!
1%
#225130000000
0!
0%
#225135000000
1!
1%
#225140000000
0!
0%
#225145000000
1!
1%
#225150000000
0!
0%
#225155000000
1!
1%
#225160000000
0!
0%
#225165000000
1!
1%
#225170000000
0!
0%
#225175000000
1!
1%
#225180000000
0!
0%
#225185000000
1!
1%
#225190000000
0!
0%
#225195000000
1!
1%
#225200000000
0!
0%
#225205000000
1!
1%
#225210000000
0!
0%
#225215000000
1!
1%
#225220000000
0!
0%
#225225000000
1!
1%
#225230000000
0!
0%
#225235000000
1!
1%
#225240000000
0!
0%
#225245000000
1!
1%
#225250000000
0!
0%
#225255000000
1!
1%
#225260000000
0!
0%
#225265000000
1!
1%
#225270000000
0!
0%
#225275000000
1!
1%
#225280000000
0!
0%
#225285000000
1!
1%
#225290000000
0!
0%
#225295000000
1!
1%
#225300000000
0!
0%
#225305000000
1!
1%
#225310000000
0!
0%
#225315000000
1!
1%
#225320000000
0!
0%
#225325000000
1!
1%
#225330000000
0!
0%
#225335000000
1!
1%
#225340000000
0!
0%
#225345000000
1!
1%
#225350000000
0!
0%
#225355000000
1!
1%
#225360000000
0!
0%
#225365000000
1!
1%
#225370000000
0!
0%
#225375000000
1!
1%
#225380000000
0!
0%
#225385000000
1!
1%
#225390000000
0!
0%
#225395000000
1!
1%
#225400000000
0!
0%
#225405000000
1!
1%
#225410000000
0!
0%
#225415000000
1!
1%
#225420000000
0!
0%
#225425000000
1!
1%
#225430000000
0!
0%
#225435000000
1!
1%
#225440000000
0!
0%
#225445000000
1!
1%
#225450000000
0!
0%
#225455000000
1!
1%
#225460000000
0!
0%
#225465000000
1!
1%
#225470000000
0!
0%
#225475000000
1!
1%
#225480000000
0!
0%
#225485000000
1!
1%
#225490000000
0!
0%
#225495000000
1!
1%
#225500000000
0!
0%
#225505000000
1!
1%
#225510000000
0!
0%
#225515000000
1!
1%
#225520000000
0!
0%
#225525000000
1!
1%
#225530000000
0!
0%
#225535000000
1!
1%
#225540000000
0!
0%
#225545000000
1!
1%
#225550000000
0!
0%
#225555000000
1!
1%
#225560000000
0!
0%
#225565000000
1!
1%
#225570000000
0!
0%
#225575000000
1!
1%
#225580000000
0!
0%
#225585000000
1!
1%
#225590000000
0!
0%
#225595000000
1!
1%
#225600000000
0!
0%
#225605000000
1!
1%
#225610000000
0!
0%
#225615000000
1!
1%
#225620000000
0!
0%
#225625000000
1!
1%
#225630000000
0!
0%
#225635000000
1!
1%
#225640000000
0!
0%
#225645000000
1!
1%
#225650000000
0!
0%
#225655000000
1!
1%
#225660000000
0!
0%
#225665000000
1!
1%
#225670000000
0!
0%
#225675000000
1!
1%
#225680000000
0!
0%
#225685000000
1!
1%
#225690000000
0!
0%
#225695000000
1!
1%
#225700000000
0!
0%
#225705000000
1!
1%
#225710000000
0!
0%
#225715000000
1!
1%
#225720000000
0!
0%
#225725000000
1!
1%
#225730000000
0!
0%
#225735000000
1!
1%
#225740000000
0!
0%
#225745000000
1!
1%
#225750000000
0!
0%
#225755000000
1!
1%
#225760000000
0!
0%
#225765000000
1!
1%
#225770000000
0!
0%
#225775000000
1!
1%
#225780000000
0!
0%
#225785000000
1!
1%
#225790000000
0!
0%
#225795000000
1!
1%
#225800000000
0!
0%
#225805000000
1!
1%
#225810000000
0!
0%
#225815000000
1!
1%
#225820000000
0!
0%
#225825000000
1!
1%
#225830000000
0!
0%
#225835000000
1!
1%
#225840000000
0!
0%
#225845000000
1!
1%
#225850000000
0!
0%
#225855000000
1!
1%
#225860000000
0!
0%
#225865000000
1!
1%
#225870000000
0!
0%
#225875000000
1!
1%
#225880000000
0!
0%
#225885000000
1!
1%
#225890000000
0!
0%
#225895000000
1!
1%
#225900000000
0!
0%
#225905000000
1!
1%
#225910000000
0!
0%
#225915000000
1!
1%
#225920000000
0!
0%
#225925000000
1!
1%
#225930000000
0!
0%
#225935000000
1!
1%
#225940000000
0!
0%
#225945000000
1!
1%
#225950000000
0!
0%
#225955000000
1!
1%
#225960000000
0!
0%
#225965000000
1!
1%
#225970000000
0!
0%
#225975000000
1!
1%
#225980000000
0!
0%
#225985000000
1!
1%
#225990000000
0!
0%
#225995000000
1!
1%
#226000000000
0!
0%
#226005000000
1!
1%
#226010000000
0!
0%
#226015000000
1!
1%
#226020000000
0!
0%
#226025000000
1!
1%
#226030000000
0!
0%
#226035000000
1!
1%
#226040000000
0!
0%
#226045000000
1!
1%
#226050000000
0!
0%
#226055000000
1!
1%
#226060000000
0!
0%
#226065000000
1!
1%
#226070000000
0!
0%
#226075000000
1!
1%
#226080000000
0!
0%
#226085000000
1!
1%
#226090000000
0!
0%
#226095000000
1!
1%
#226100000000
0!
0%
#226105000000
1!
1%
#226110000000
0!
0%
#226115000000
1!
1%
#226120000000
0!
0%
#226125000000
1!
1%
#226130000000
0!
0%
#226135000000
1!
1%
#226140000000
0!
0%
#226145000000
1!
1%
#226150000000
0!
0%
#226155000000
1!
1%
#226160000000
0!
0%
#226165000000
1!
1%
#226170000000
0!
0%
#226175000000
1!
1%
#226180000000
0!
0%
#226185000000
1!
1%
#226190000000
0!
0%
#226195000000
1!
1%
#226200000000
0!
0%
#226205000000
1!
1%
#226210000000
0!
0%
#226215000000
1!
1%
#226220000000
0!
0%
#226225000000
1!
1%
#226230000000
0!
0%
#226235000000
1!
1%
#226240000000
0!
0%
#226245000000
1!
1%
#226250000000
0!
0%
#226255000000
1!
1%
#226260000000
0!
0%
#226265000000
1!
1%
#226270000000
0!
0%
#226275000000
1!
1%
#226280000000
0!
0%
#226285000000
1!
1%
#226290000000
0!
0%
#226295000000
1!
1%
#226300000000
0!
0%
#226305000000
1!
1%
#226310000000
0!
0%
#226315000000
1!
1%
#226320000000
0!
0%
#226325000000
1!
1%
#226330000000
0!
0%
#226335000000
1!
1%
#226340000000
0!
0%
#226345000000
1!
1%
#226350000000
0!
0%
#226355000000
1!
1%
#226360000000
0!
0%
#226365000000
1!
1%
#226370000000
0!
0%
#226375000000
1!
1%
#226380000000
0!
0%
#226385000000
1!
1%
#226390000000
0!
0%
#226395000000
1!
1%
#226400000000
0!
0%
#226405000000
1!
1%
#226410000000
0!
0%
#226415000000
1!
1%
#226420000000
0!
0%
#226425000000
1!
1%
#226430000000
0!
0%
#226435000000
1!
1%
#226440000000
0!
0%
#226445000000
1!
1%
#226450000000
0!
0%
#226455000000
1!
1%
#226460000000
0!
0%
#226465000000
1!
1%
#226470000000
0!
0%
#226475000000
1!
1%
#226480000000
0!
0%
#226485000000
1!
1%
#226490000000
0!
0%
#226495000000
1!
1%
#226500000000
0!
0%
#226505000000
1!
1%
#226510000000
0!
0%
#226515000000
1!
1%
#226520000000
0!
0%
#226525000000
1!
1%
#226530000000
0!
0%
#226535000000
1!
1%
#226540000000
0!
0%
#226545000000
1!
1%
#226550000000
0!
0%
#226555000000
1!
1%
#226560000000
0!
0%
#226565000000
1!
1%
#226570000000
0!
0%
#226575000000
1!
1%
#226580000000
0!
0%
#226585000000
1!
1%
#226590000000
0!
0%
#226595000000
1!
1%
#226600000000
0!
0%
#226605000000
1!
1%
#226610000000
0!
0%
#226615000000
1!
1%
#226620000000
0!
0%
#226625000000
1!
1%
#226630000000
0!
0%
#226635000000
1!
1%
#226640000000
0!
0%
#226645000000
1!
1%
#226650000000
0!
0%
#226655000000
1!
1%
#226660000000
0!
0%
#226665000000
1!
1%
#226670000000
0!
0%
#226675000000
1!
1%
#226680000000
0!
0%
#226685000000
1!
1%
#226690000000
0!
0%
#226695000000
1!
1%
#226700000000
0!
0%
#226705000000
1!
1%
#226710000000
0!
0%
#226715000000
1!
1%
#226720000000
0!
0%
#226725000000
1!
1%
#226730000000
0!
0%
#226735000000
1!
1%
#226740000000
0!
0%
#226745000000
1!
1%
#226750000000
0!
0%
#226755000000
1!
1%
#226760000000
0!
0%
#226765000000
1!
1%
#226770000000
0!
0%
#226775000000
1!
1%
#226780000000
0!
0%
#226785000000
1!
1%
#226790000000
0!
0%
#226795000000
1!
1%
#226800000000
0!
0%
#226805000000
1!
1%
#226810000000
0!
0%
#226815000000
1!
1%
#226820000000
0!
0%
#226825000000
1!
1%
#226830000000
0!
0%
#226835000000
1!
1%
#226840000000
0!
0%
#226845000000
1!
1%
#226850000000
0!
0%
#226855000000
1!
1%
#226860000000
0!
0%
#226865000000
1!
1%
#226870000000
0!
0%
#226875000000
1!
1%
#226880000000
0!
0%
#226885000000
1!
1%
#226890000000
0!
0%
#226895000000
1!
1%
#226900000000
0!
0%
#226905000000
1!
1%
#226910000000
0!
0%
#226915000000
1!
1%
#226920000000
0!
0%
#226925000000
1!
1%
#226930000000
0!
0%
#226935000000
1!
1%
#226940000000
0!
0%
#226945000000
1!
1%
#226950000000
0!
0%
#226955000000
1!
1%
#226960000000
0!
0%
#226965000000
1!
1%
#226970000000
0!
0%
#226975000000
1!
1%
#226980000000
0!
0%
#226985000000
1!
1%
#226990000000
0!
0%
#226995000000
1!
1%
#227000000000
0!
0%
#227005000000
1!
1%
#227010000000
0!
0%
#227015000000
1!
1%
#227020000000
0!
0%
#227025000000
1!
1%
#227030000000
0!
0%
#227035000000
1!
1%
#227040000000
0!
0%
#227045000000
1!
1%
#227050000000
0!
0%
#227055000000
1!
1%
#227060000000
0!
0%
#227065000000
1!
1%
#227070000000
0!
0%
#227075000000
1!
1%
#227080000000
0!
0%
#227085000000
1!
1%
#227090000000
0!
0%
#227095000000
1!
1%
#227100000000
0!
0%
#227105000000
1!
1%
#227110000000
0!
0%
#227115000000
1!
1%
#227120000000
0!
0%
#227125000000
1!
1%
#227130000000
0!
0%
#227135000000
1!
1%
#227140000000
0!
0%
#227145000000
1!
1%
#227150000000
0!
0%
#227155000000
1!
1%
#227160000000
0!
0%
#227165000000
1!
1%
#227170000000
0!
0%
#227175000000
1!
1%
#227180000000
0!
0%
#227185000000
1!
1%
#227190000000
0!
0%
#227195000000
1!
1%
#227200000000
0!
0%
#227205000000
1!
1%
#227210000000
0!
0%
#227215000000
1!
1%
#227220000000
0!
0%
#227225000000
1!
1%
#227230000000
0!
0%
#227235000000
1!
1%
#227240000000
0!
0%
#227245000000
1!
1%
#227250000000
0!
0%
#227255000000
1!
1%
#227260000000
0!
0%
#227265000000
1!
1%
#227270000000
0!
0%
#227275000000
1!
1%
#227280000000
0!
0%
#227285000000
1!
1%
#227290000000
0!
0%
#227295000000
1!
1%
#227300000000
0!
0%
#227305000000
1!
1%
#227310000000
0!
0%
#227315000000
1!
1%
#227320000000
0!
0%
#227325000000
1!
1%
#227330000000
0!
0%
#227335000000
1!
1%
#227340000000
0!
0%
#227345000000
1!
1%
#227350000000
0!
0%
#227355000000
1!
1%
#227360000000
0!
0%
#227365000000
1!
1%
#227370000000
0!
0%
#227375000000
1!
1%
#227380000000
0!
0%
#227385000000
1!
1%
#227390000000
0!
0%
#227395000000
1!
1%
#227400000000
0!
0%
#227405000000
1!
1%
#227410000000
0!
0%
#227415000000
1!
1%
#227420000000
0!
0%
#227425000000
1!
1%
#227430000000
0!
0%
#227435000000
1!
1%
#227440000000
0!
0%
#227445000000
1!
1%
#227450000000
0!
0%
#227455000000
1!
1%
#227460000000
0!
0%
#227465000000
1!
1%
#227470000000
0!
0%
#227475000000
1!
1%
#227480000000
0!
0%
#227485000000
1!
1%
#227490000000
0!
0%
#227495000000
1!
1%
#227500000000
0!
0%
#227505000000
1!
1%
#227510000000
0!
0%
#227515000000
1!
1%
#227520000000
0!
0%
#227525000000
1!
1%
#227530000000
0!
0%
#227535000000
1!
1%
#227540000000
0!
0%
#227545000000
1!
1%
#227550000000
0!
0%
#227555000000
1!
1%
#227560000000
0!
0%
#227565000000
1!
1%
#227570000000
0!
0%
#227575000000
1!
1%
#227580000000
0!
0%
#227585000000
1!
1%
#227590000000
0!
0%
#227595000000
1!
1%
#227600000000
0!
0%
#227605000000
1!
1%
#227610000000
0!
0%
#227615000000
1!
1%
#227620000000
0!
0%
#227625000000
1!
1%
#227630000000
0!
0%
#227635000000
1!
1%
#227640000000
0!
0%
#227645000000
1!
1%
#227650000000
0!
0%
#227655000000
1!
1%
#227660000000
0!
0%
#227665000000
1!
1%
#227670000000
0!
0%
#227675000000
1!
1%
#227680000000
0!
0%
#227685000000
1!
1%
#227690000000
0!
0%
#227695000000
1!
1%
#227700000000
0!
0%
#227705000000
1!
1%
#227710000000
0!
0%
#227715000000
1!
1%
#227720000000
0!
0%
#227725000000
1!
1%
#227730000000
0!
0%
#227735000000
1!
1%
#227740000000
0!
0%
#227745000000
1!
1%
#227750000000
0!
0%
#227755000000
1!
1%
#227760000000
0!
0%
#227765000000
1!
1%
#227770000000
0!
0%
#227775000000
1!
1%
#227780000000
0!
0%
#227785000000
1!
1%
#227790000000
0!
0%
#227795000000
1!
1%
#227800000000
0!
0%
#227805000000
1!
1%
#227810000000
0!
0%
#227815000000
1!
1%
#227820000000
0!
0%
#227825000000
1!
1%
#227830000000
0!
0%
#227835000000
1!
1%
#227840000000
0!
0%
#227845000000
1!
1%
#227850000000
0!
0%
#227855000000
1!
1%
#227860000000
0!
0%
#227865000000
1!
1%
#227870000000
0!
0%
#227875000000
1!
1%
#227880000000
0!
0%
#227885000000
1!
1%
#227890000000
0!
0%
#227895000000
1!
1%
#227900000000
0!
0%
#227905000000
1!
1%
#227910000000
0!
0%
#227915000000
1!
1%
#227920000000
0!
0%
#227925000000
1!
1%
#227930000000
0!
0%
#227935000000
1!
1%
#227940000000
0!
0%
#227945000000
1!
1%
#227950000000
0!
0%
#227955000000
1!
1%
#227960000000
0!
0%
#227965000000
1!
1%
#227970000000
0!
0%
#227975000000
1!
1%
#227980000000
0!
0%
#227985000000
1!
1%
#227990000000
0!
0%
#227995000000
1!
1%
#228000000000
0!
0%
#228005000000
1!
1%
#228010000000
0!
0%
#228015000000
1!
1%
#228020000000
0!
0%
#228025000000
1!
1%
#228030000000
0!
0%
#228035000000
1!
1%
#228040000000
0!
0%
#228045000000
1!
1%
#228050000000
0!
0%
#228055000000
1!
1%
#228060000000
0!
0%
#228065000000
1!
1%
#228070000000
0!
0%
#228075000000
1!
1%
#228080000000
0!
0%
#228085000000
1!
1%
#228090000000
0!
0%
#228095000000
1!
1%
#228100000000
0!
0%
#228105000000
1!
1%
#228110000000
0!
0%
#228115000000
1!
1%
#228120000000
0!
0%
#228125000000
1!
1%
#228130000000
0!
0%
#228135000000
1!
1%
#228140000000
0!
0%
#228145000000
1!
1%
#228150000000
0!
0%
#228155000000
1!
1%
#228160000000
0!
0%
#228165000000
1!
1%
#228170000000
0!
0%
#228175000000
1!
1%
#228180000000
0!
0%
#228185000000
1!
1%
#228190000000
0!
0%
#228195000000
1!
1%
#228200000000
0!
0%
#228205000000
1!
1%
#228210000000
0!
0%
#228215000000
1!
1%
#228220000000
0!
0%
#228225000000
1!
1%
#228230000000
0!
0%
#228235000000
1!
1%
#228240000000
0!
0%
#228245000000
1!
1%
#228250000000
0!
0%
#228255000000
1!
1%
#228260000000
0!
0%
#228265000000
1!
1%
#228270000000
0!
0%
#228275000000
1!
1%
#228280000000
0!
0%
#228285000000
1!
1%
#228290000000
0!
0%
#228295000000
1!
1%
#228300000000
0!
0%
#228305000000
1!
1%
#228310000000
0!
0%
#228315000000
1!
1%
#228320000000
0!
0%
#228325000000
1!
1%
#228330000000
0!
0%
#228335000000
1!
1%
#228340000000
0!
0%
#228345000000
1!
1%
#228350000000
0!
0%
#228355000000
1!
1%
#228360000000
0!
0%
#228365000000
1!
1%
#228370000000
0!
0%
#228375000000
1!
1%
#228380000000
0!
0%
#228385000000
1!
1%
#228390000000
0!
0%
#228395000000
1!
1%
#228400000000
0!
0%
#228405000000
1!
1%
#228410000000
0!
0%
#228415000000
1!
1%
#228420000000
0!
0%
#228425000000
1!
1%
#228430000000
0!
0%
#228435000000
1!
1%
#228440000000
0!
0%
#228445000000
1!
1%
#228450000000
0!
0%
#228455000000
1!
1%
#228460000000
0!
0%
#228465000000
1!
1%
#228470000000
0!
0%
#228475000000
1!
1%
#228480000000
0!
0%
#228485000000
1!
1%
#228490000000
0!
0%
#228495000000
1!
1%
#228500000000
0!
0%
#228505000000
1!
1%
#228510000000
0!
0%
#228515000000
1!
1%
#228520000000
0!
0%
#228525000000
1!
1%
#228530000000
0!
0%
#228535000000
1!
1%
#228540000000
0!
0%
#228545000000
1!
1%
#228550000000
0!
0%
#228555000000
1!
1%
#228560000000
0!
0%
#228565000000
1!
1%
#228570000000
0!
0%
#228575000000
1!
1%
#228580000000
0!
0%
#228585000000
1!
1%
#228590000000
0!
0%
#228595000000
1!
1%
#228600000000
0!
0%
#228605000000
1!
1%
#228610000000
0!
0%
#228615000000
1!
1%
#228620000000
0!
0%
#228625000000
1!
1%
#228630000000
0!
0%
#228635000000
1!
1%
#228640000000
0!
0%
#228645000000
1!
1%
#228650000000
0!
0%
#228655000000
1!
1%
#228660000000
0!
0%
#228665000000
1!
1%
#228670000000
0!
0%
#228675000000
1!
1%
#228680000000
0!
0%
#228685000000
1!
1%
#228690000000
0!
0%
#228695000000
1!
1%
#228700000000
0!
0%
#228705000000
1!
1%
#228710000000
0!
0%
#228715000000
1!
1%
#228720000000
0!
0%
#228725000000
1!
1%
#228730000000
0!
0%
#228735000000
1!
1%
#228740000000
0!
0%
#228745000000
1!
1%
#228750000000
0!
0%
#228755000000
1!
1%
#228760000000
0!
0%
#228765000000
1!
1%
#228770000000
0!
0%
#228775000000
1!
1%
#228780000000
0!
0%
#228785000000
1!
1%
#228790000000
0!
0%
#228795000000
1!
1%
#228800000000
0!
0%
#228805000000
1!
1%
#228810000000
0!
0%
#228815000000
1!
1%
#228820000000
0!
0%
#228825000000
1!
1%
#228830000000
0!
0%
#228835000000
1!
1%
#228840000000
0!
0%
#228845000000
1!
1%
#228850000000
0!
0%
#228855000000
1!
1%
#228860000000
0!
0%
#228865000000
1!
1%
#228870000000
0!
0%
#228875000000
1!
1%
#228880000000
0!
0%
#228885000000
1!
1%
#228890000000
0!
0%
#228895000000
1!
1%
#228900000000
0!
0%
#228905000000
1!
1%
#228910000000
0!
0%
#228915000000
1!
1%
#228920000000
0!
0%
#228925000000
1!
1%
#228930000000
0!
0%
#228935000000
1!
1%
#228940000000
0!
0%
#228945000000
1!
1%
#228950000000
0!
0%
#228955000000
1!
1%
#228960000000
0!
0%
#228965000000
1!
1%
#228970000000
0!
0%
#228975000000
1!
1%
#228980000000
0!
0%
#228985000000
1!
1%
#228990000000
0!
0%
#228995000000
1!
1%
#229000000000
0!
0%
#229005000000
1!
1%
#229010000000
0!
0%
#229015000000
1!
1%
#229020000000
0!
0%
#229025000000
1!
1%
#229030000000
0!
0%
#229035000000
1!
1%
#229040000000
0!
0%
#229045000000
1!
1%
#229050000000
0!
0%
#229055000000
1!
1%
#229060000000
0!
0%
#229065000000
1!
1%
#229070000000
0!
0%
#229075000000
1!
1%
#229080000000
0!
0%
#229085000000
1!
1%
#229090000000
0!
0%
#229095000000
1!
1%
#229100000000
0!
0%
#229105000000
1!
1%
#229110000000
0!
0%
#229115000000
1!
1%
#229120000000
0!
0%
#229125000000
1!
1%
#229130000000
0!
0%
#229135000000
1!
1%
#229140000000
0!
0%
#229145000000
1!
1%
#229150000000
0!
0%
#229155000000
1!
1%
#229160000000
0!
0%
#229165000000
1!
1%
#229170000000
0!
0%
#229175000000
1!
1%
#229180000000
0!
0%
#229185000000
1!
1%
#229190000000
0!
0%
#229195000000
1!
1%
#229200000000
0!
0%
#229205000000
1!
1%
#229210000000
0!
0%
#229215000000
1!
1%
#229220000000
0!
0%
#229225000000
1!
1%
#229230000000
0!
0%
#229235000000
1!
1%
#229240000000
0!
0%
#229245000000
1!
1%
#229250000000
0!
0%
#229255000000
1!
1%
#229260000000
0!
0%
#229265000000
1!
1%
#229270000000
0!
0%
#229275000000
1!
1%
#229280000000
0!
0%
#229285000000
1!
1%
#229290000000
0!
0%
#229295000000
1!
1%
#229300000000
0!
0%
#229305000000
1!
1%
#229310000000
0!
0%
#229315000000
1!
1%
#229320000000
0!
0%
#229325000000
1!
1%
#229330000000
0!
0%
#229335000000
1!
1%
#229340000000
0!
0%
#229345000000
1!
1%
#229350000000
0!
0%
#229355000000
1!
1%
#229360000000
0!
0%
#229365000000
1!
1%
#229370000000
0!
0%
#229375000000
1!
1%
#229380000000
0!
0%
#229385000000
1!
1%
#229390000000
0!
0%
#229395000000
1!
1%
#229400000000
0!
0%
#229405000000
1!
1%
#229410000000
0!
0%
#229415000000
1!
1%
#229420000000
0!
0%
#229425000000
1!
1%
#229430000000
0!
0%
#229435000000
1!
1%
#229440000000
0!
0%
#229445000000
1!
1%
#229450000000
0!
0%
#229455000000
1!
1%
#229460000000
0!
0%
#229465000000
1!
1%
#229470000000
0!
0%
#229475000000
1!
1%
#229480000000
0!
0%
#229485000000
1!
1%
#229490000000
0!
0%
#229495000000
1!
1%
#229500000000
0!
0%
#229505000000
1!
1%
#229510000000
0!
0%
#229515000000
1!
1%
#229520000000
0!
0%
#229525000000
1!
1%
#229530000000
0!
0%
#229535000000
1!
1%
#229540000000
0!
0%
#229545000000
1!
1%
#229550000000
0!
0%
#229555000000
1!
1%
#229560000000
0!
0%
#229565000000
1!
1%
#229570000000
0!
0%
#229575000000
1!
1%
#229580000000
0!
0%
#229585000000
1!
1%
#229590000000
0!
0%
#229595000000
1!
1%
#229600000000
0!
0%
#229605000000
1!
1%
#229610000000
0!
0%
#229615000000
1!
1%
#229620000000
0!
0%
#229625000000
1!
1%
#229630000000
0!
0%
#229635000000
1!
1%
#229640000000
0!
0%
#229645000000
1!
1%
#229650000000
0!
0%
#229655000000
1!
1%
#229660000000
0!
0%
#229665000000
1!
1%
#229670000000
0!
0%
#229675000000
1!
1%
#229680000000
0!
0%
#229685000000
1!
1%
#229690000000
0!
0%
#229695000000
1!
1%
#229700000000
0!
0%
#229705000000
1!
1%
#229710000000
0!
0%
#229715000000
1!
1%
#229720000000
0!
0%
#229725000000
1!
1%
#229730000000
0!
0%
#229735000000
1!
1%
#229740000000
0!
0%
#229745000000
1!
1%
#229750000000
0!
0%
#229755000000
1!
1%
#229760000000
0!
0%
#229765000000
1!
1%
#229770000000
0!
0%
#229775000000
1!
1%
#229780000000
0!
0%
#229785000000
1!
1%
#229790000000
0!
0%
#229795000000
1!
1%
#229800000000
0!
0%
#229805000000
1!
1%
#229810000000
0!
0%
#229815000000
1!
1%
#229820000000
0!
0%
#229825000000
1!
1%
#229830000000
0!
0%
#229835000000
1!
1%
#229840000000
0!
0%
#229845000000
1!
1%
#229850000000
0!
0%
#229855000000
1!
1%
#229860000000
0!
0%
#229865000000
1!
1%
#229870000000
0!
0%
#229875000000
1!
1%
#229880000000
0!
0%
#229885000000
1!
1%
#229890000000
0!
0%
#229895000000
1!
1%
#229900000000
0!
0%
#229905000000
1!
1%
#229910000000
0!
0%
#229915000000
1!
1%
#229920000000
0!
0%
#229925000000
1!
1%
#229930000000
0!
0%
#229935000000
1!
1%
#229940000000
0!
0%
#229945000000
1!
1%
#229950000000
0!
0%
#229955000000
1!
1%
#229960000000
0!
0%
#229965000000
1!
1%
#229970000000
0!
0%
#229975000000
1!
1%
#229980000000
0!
0%
#229985000000
1!
1%
#229990000000
0!
0%
#229995000000
1!
1%
#230000000000
0!
0%
#230005000000
1!
1%
#230010000000
0!
0%
#230015000000
1!
1%
#230020000000
0!
0%
#230025000000
1!
1%
#230030000000
0!
0%
#230035000000
1!
1%
#230040000000
0!
0%
#230045000000
1!
1%
#230050000000
0!
0%
#230055000000
1!
1%
#230060000000
0!
0%
#230065000000
1!
1%
#230070000000
0!
0%
#230075000000
1!
1%
#230080000000
0!
0%
#230085000000
1!
1%
#230090000000
0!
0%
#230095000000
1!
1%
#230100000000
0!
0%
#230105000000
1!
1%
#230110000000
0!
0%
#230115000000
1!
1%
#230120000000
0!
0%
#230125000000
1!
1%
#230130000000
0!
0%
#230135000000
1!
1%
#230140000000
0!
0%
#230145000000
1!
1%
#230150000000
0!
0%
#230155000000
1!
1%
#230160000000
0!
0%
#230165000000
1!
1%
#230170000000
0!
0%
#230175000000
1!
1%
#230180000000
0!
0%
#230185000000
1!
1%
#230190000000
0!
0%
#230195000000
1!
1%
#230200000000
0!
0%
#230205000000
1!
1%
#230210000000
0!
0%
#230215000000
1!
1%
#230220000000
0!
0%
#230225000000
1!
1%
#230230000000
0!
0%
#230235000000
1!
1%
#230240000000
0!
0%
#230245000000
1!
1%
#230250000000
0!
0%
#230255000000
1!
1%
#230260000000
0!
0%
#230265000000
1!
1%
#230270000000
0!
0%
#230275000000
1!
1%
#230280000000
0!
0%
#230285000000
1!
1%
#230290000000
0!
0%
#230295000000
1!
1%
#230300000000
0!
0%
#230305000000
1!
1%
#230310000000
0!
0%
#230315000000
1!
1%
#230320000000
0!
0%
#230325000000
1!
1%
#230330000000
0!
0%
#230335000000
1!
1%
#230340000000
0!
0%
#230345000000
1!
1%
#230350000000
0!
0%
#230355000000
1!
1%
#230360000000
0!
0%
#230365000000
1!
1%
#230370000000
0!
0%
#230375000000
1!
1%
#230380000000
0!
0%
#230385000000
1!
1%
#230390000000
0!
0%
#230395000000
1!
1%
#230400000000
0!
0%
#230405000000
1!
1%
#230410000000
0!
0%
#230415000000
1!
1%
#230420000000
0!
0%
#230425000000
1!
1%
#230430000000
0!
0%
#230435000000
1!
1%
#230440000000
0!
0%
#230445000000
1!
1%
#230450000000
0!
0%
#230455000000
1!
1%
#230460000000
0!
0%
#230465000000
1!
1%
#230470000000
0!
0%
#230475000000
1!
1%
#230480000000
0!
0%
#230485000000
1!
1%
#230490000000
0!
0%
#230495000000
1!
1%
#230500000000
0!
0%
#230505000000
1!
1%
#230510000000
0!
0%
#230515000000
1!
1%
#230520000000
0!
0%
#230525000000
1!
1%
#230530000000
0!
0%
#230535000000
1!
1%
#230540000000
0!
0%
#230545000000
1!
1%
#230550000000
0!
0%
#230555000000
1!
1%
#230560000000
0!
0%
#230565000000
1!
1%
#230570000000
0!
0%
#230575000000
1!
1%
#230580000000
0!
0%
#230585000000
1!
1%
#230590000000
0!
0%
#230595000000
1!
1%
#230600000000
0!
0%
#230605000000
1!
1%
#230610000000
0!
0%
#230615000000
1!
1%
#230620000000
0!
0%
#230625000000
1!
1%
#230630000000
0!
0%
#230635000000
1!
1%
#230640000000
0!
0%
#230645000000
1!
1%
#230650000000
0!
0%
#230655000000
1!
1%
#230660000000
0!
0%
#230665000000
1!
1%
#230670000000
0!
0%
#230675000000
1!
1%
#230680000000
0!
0%
#230685000000
1!
1%
#230690000000
0!
0%
#230695000000
1!
1%
#230700000000
0!
0%
#230705000000
1!
1%
#230710000000
0!
0%
#230715000000
1!
1%
#230720000000
0!
0%
#230725000000
1!
1%
#230730000000
0!
0%
#230735000000
1!
1%
#230740000000
0!
0%
#230745000000
1!
1%
#230750000000
0!
0%
#230755000000
1!
1%
#230760000000
0!
0%
#230765000000
1!
1%
#230770000000
0!
0%
#230775000000
1!
1%
#230780000000
0!
0%
#230785000000
1!
1%
#230790000000
0!
0%
#230795000000
1!
1%
#230800000000
0!
0%
#230805000000
1!
1%
#230810000000
0!
0%
#230815000000
1!
1%
#230820000000
0!
0%
#230825000000
1!
1%
#230830000000
0!
0%
#230835000000
1!
1%
#230840000000
0!
0%
#230845000000
1!
1%
#230850000000
0!
0%
#230855000000
1!
1%
#230860000000
0!
0%
#230865000000
1!
1%
#230870000000
0!
0%
#230875000000
1!
1%
#230880000000
0!
0%
#230885000000
1!
1%
#230890000000
0!
0%
#230895000000
1!
1%
#230900000000
0!
0%
#230905000000
1!
1%
#230910000000
0!
0%
#230915000000
1!
1%
#230920000000
0!
0%
#230925000000
1!
1%
#230930000000
0!
0%
#230935000000
1!
1%
#230940000000
0!
0%
#230945000000
1!
1%
#230950000000
0!
0%
#230955000000
1!
1%
#230960000000
0!
0%
#230965000000
1!
1%
#230970000000
0!
0%
#230975000000
1!
1%
#230980000000
0!
0%
#230985000000
1!
1%
#230990000000
0!
0%
#230995000000
1!
1%
#231000000000
0!
0%
#231005000000
1!
1%
#231010000000
0!
0%
#231015000000
1!
1%
#231020000000
0!
0%
#231025000000
1!
1%
#231030000000
0!
0%
#231035000000
1!
1%
#231040000000
0!
0%
#231045000000
1!
1%
#231050000000
0!
0%
#231055000000
1!
1%
#231060000000
0!
0%
#231065000000
1!
1%
#231070000000
0!
0%
#231075000000
1!
1%
#231080000000
0!
0%
#231085000000
1!
1%
#231090000000
0!
0%
#231095000000
1!
1%
#231100000000
0!
0%
#231105000000
1!
1%
#231110000000
0!
0%
#231115000000
1!
1%
#231120000000
0!
0%
#231125000000
1!
1%
#231130000000
0!
0%
#231135000000
1!
1%
#231140000000
0!
0%
#231145000000
1!
1%
#231150000000
0!
0%
#231155000000
1!
1%
#231160000000
0!
0%
#231165000000
1!
1%
#231170000000
0!
0%
#231175000000
1!
1%
#231180000000
0!
0%
#231185000000
1!
1%
#231190000000
0!
0%
#231195000000
1!
1%
#231200000000
0!
0%
#231205000000
1!
1%
#231210000000
0!
0%
#231215000000
1!
1%
#231220000000
0!
0%
#231225000000
1!
1%
#231230000000
0!
0%
#231235000000
1!
1%
#231240000000
0!
0%
#231245000000
1!
1%
#231250000000
0!
0%
#231255000000
1!
1%
#231260000000
0!
0%
#231265000000
1!
1%
#231270000000
0!
0%
#231275000000
1!
1%
#231280000000
0!
0%
#231285000000
1!
1%
#231290000000
0!
0%
#231295000000
1!
1%
#231300000000
0!
0%
#231305000000
1!
1%
#231310000000
0!
0%
#231315000000
1!
1%
#231320000000
0!
0%
#231325000000
1!
1%
#231330000000
0!
0%
#231335000000
1!
1%
#231340000000
0!
0%
#231345000000
1!
1%
#231350000000
0!
0%
#231355000000
1!
1%
#231360000000
0!
0%
#231365000000
1!
1%
#231370000000
0!
0%
#231375000000
1!
1%
#231380000000
0!
0%
#231385000000
1!
1%
#231390000000
0!
0%
#231395000000
1!
1%
#231400000000
0!
0%
#231405000000
1!
1%
#231410000000
0!
0%
#231415000000
1!
1%
#231420000000
0!
0%
#231425000000
1!
1%
#231430000000
0!
0%
#231435000000
1!
1%
#231440000000
0!
0%
#231445000000
1!
1%
#231450000000
0!
0%
#231455000000
1!
1%
#231460000000
0!
0%
#231465000000
1!
1%
#231470000000
0!
0%
#231475000000
1!
1%
#231480000000
0!
0%
#231485000000
1!
1%
#231490000000
0!
0%
#231495000000
1!
1%
#231500000000
0!
0%
#231505000000
1!
1%
#231510000000
0!
0%
#231515000000
1!
1%
#231520000000
0!
0%
#231525000000
1!
1%
#231530000000
0!
0%
#231535000000
1!
1%
#231540000000
0!
0%
#231545000000
1!
1%
#231550000000
0!
0%
#231555000000
1!
1%
#231560000000
0!
0%
#231565000000
1!
1%
#231570000000
0!
0%
#231575000000
1!
1%
#231580000000
0!
0%
#231585000000
1!
1%
#231590000000
0!
0%
#231595000000
1!
1%
#231600000000
0!
0%
#231605000000
1!
1%
#231610000000
0!
0%
#231615000000
1!
1%
#231620000000
0!
0%
#231625000000
1!
1%
#231630000000
0!
0%
#231635000000
1!
1%
#231640000000
0!
0%
#231645000000
1!
1%
#231650000000
0!
0%
#231655000000
1!
1%
#231660000000
0!
0%
#231665000000
1!
1%
#231670000000
0!
0%
#231675000000
1!
1%
#231680000000
0!
0%
#231685000000
1!
1%
#231690000000
0!
0%
#231695000000
1!
1%
#231700000000
0!
0%
#231705000000
1!
1%
#231710000000
0!
0%
#231715000000
1!
1%
#231720000000
0!
0%
#231725000000
1!
1%
#231730000000
0!
0%
#231735000000
1!
1%
#231740000000
0!
0%
#231745000000
1!
1%
#231750000000
0!
0%
#231755000000
1!
1%
#231760000000
0!
0%
#231765000000
1!
1%
#231770000000
0!
0%
#231775000000
1!
1%
#231780000000
0!
0%
#231785000000
1!
1%
#231790000000
0!
0%
#231795000000
1!
1%
#231800000000
0!
0%
#231805000000
1!
1%
#231810000000
0!
0%
#231815000000
1!
1%
#231820000000
0!
0%
#231825000000
1!
1%
#231830000000
0!
0%
#231835000000
1!
1%
#231840000000
0!
0%
#231845000000
1!
1%
#231850000000
0!
0%
#231855000000
1!
1%
#231860000000
0!
0%
#231865000000
1!
1%
#231870000000
0!
0%
#231875000000
1!
1%
#231880000000
0!
0%
#231885000000
1!
1%
#231890000000
0!
0%
#231895000000
1!
1%
#231900000000
0!
0%
#231905000000
1!
1%
#231910000000
0!
0%
#231915000000
1!
1%
#231920000000
0!
0%
#231925000000
1!
1%
#231930000000
0!
0%
#231935000000
1!
1%
#231940000000
0!
0%
#231945000000
1!
1%
#231950000000
0!
0%
#231955000000
1!
1%
#231960000000
0!
0%
#231965000000
1!
1%
#231970000000
0!
0%
#231975000000
1!
1%
#231980000000
0!
0%
#231985000000
1!
1%
#231990000000
0!
0%
#231995000000
1!
1%
#232000000000
0!
0%
#232005000000
1!
1%
#232010000000
0!
0%
#232015000000
1!
1%
#232020000000
0!
0%
#232025000000
1!
1%
#232030000000
0!
0%
#232035000000
1!
1%
#232040000000
0!
0%
#232045000000
1!
1%
#232050000000
0!
0%
#232055000000
1!
1%
#232060000000
0!
0%
#232065000000
1!
1%
#232070000000
0!
0%
#232075000000
1!
1%
#232080000000
0!
0%
#232085000000
1!
1%
#232090000000
0!
0%
#232095000000
1!
1%
#232100000000
0!
0%
#232105000000
1!
1%
#232110000000
0!
0%
#232115000000
1!
1%
#232120000000
0!
0%
#232125000000
1!
1%
#232130000000
0!
0%
#232135000000
1!
1%
#232140000000
0!
0%
#232145000000
1!
1%
#232150000000
0!
0%
#232155000000
1!
1%
#232160000000
0!
0%
#232165000000
1!
1%
#232170000000
0!
0%
#232175000000
1!
1%
#232180000000
0!
0%
#232185000000
1!
1%
#232190000000
0!
0%
#232195000000
1!
1%
#232200000000
0!
0%
#232205000000
1!
1%
#232210000000
0!
0%
#232215000000
1!
1%
#232220000000
0!
0%
#232225000000
1!
1%
#232230000000
0!
0%
#232235000000
1!
1%
#232240000000
0!
0%
#232245000000
1!
1%
#232250000000
0!
0%
#232255000000
1!
1%
#232260000000
0!
0%
#232265000000
1!
1%
#232270000000
0!
0%
#232275000000
1!
1%
#232280000000
0!
0%
#232285000000
1!
1%
#232290000000
0!
0%
#232295000000
1!
1%
#232300000000
0!
0%
#232305000000
1!
1%
#232310000000
0!
0%
#232315000000
1!
1%
#232320000000
0!
0%
#232325000000
1!
1%
#232330000000
0!
0%
#232335000000
1!
1%
#232340000000
0!
0%
#232345000000
1!
1%
#232350000000
0!
0%
#232355000000
1!
1%
#232360000000
0!
0%
#232365000000
1!
1%
#232370000000
0!
0%
#232375000000
1!
1%
#232380000000
0!
0%
#232385000000
1!
1%
#232390000000
0!
0%
#232395000000
1!
1%
#232400000000
0!
0%
#232405000000
1!
1%
#232410000000
0!
0%
#232415000000
1!
1%
#232420000000
0!
0%
#232425000000
1!
1%
#232430000000
0!
0%
#232435000000
1!
1%
#232440000000
0!
0%
#232445000000
1!
1%
#232450000000
0!
0%
#232455000000
1!
1%
#232460000000
0!
0%
#232465000000
1!
1%
#232470000000
0!
0%
#232475000000
1!
1%
#232480000000
0!
0%
#232485000000
1!
1%
#232490000000
0!
0%
#232495000000
1!
1%
#232500000000
0!
0%
#232505000000
1!
1%
#232510000000
0!
0%
#232515000000
1!
1%
#232520000000
0!
0%
#232525000000
1!
1%
#232530000000
0!
0%
#232535000000
1!
1%
#232540000000
0!
0%
#232545000000
1!
1%
#232550000000
0!
0%
#232555000000
1!
1%
#232560000000
0!
0%
#232565000000
1!
1%
#232570000000
0!
0%
#232575000000
1!
1%
#232580000000
0!
0%
#232585000000
1!
1%
#232590000000
0!
0%
#232595000000
1!
1%
#232600000000
0!
0%
#232605000000
1!
1%
#232610000000
0!
0%
#232615000000
1!
1%
#232620000000
0!
0%
#232625000000
1!
1%
#232630000000
0!
0%
#232635000000
1!
1%
#232640000000
0!
0%
#232645000000
1!
1%
#232650000000
0!
0%
#232655000000
1!
1%
#232660000000
0!
0%
#232665000000
1!
1%
#232670000000
0!
0%
#232675000000
1!
1%
#232680000000
0!
0%
#232685000000
1!
1%
#232690000000
0!
0%
#232695000000
1!
1%
#232700000000
0!
0%
#232705000000
1!
1%
#232710000000
0!
0%
#232715000000
1!
1%
#232720000000
0!
0%
#232725000000
1!
1%
#232730000000
0!
0%
#232735000000
1!
1%
#232740000000
0!
0%
#232745000000
1!
1%
#232750000000
0!
0%
#232755000000
1!
1%
#232760000000
0!
0%
#232765000000
1!
1%
#232770000000
0!
0%
#232775000000
1!
1%
#232780000000
0!
0%
#232785000000
1!
1%
#232790000000
0!
0%
#232795000000
1!
1%
#232800000000
0!
0%
#232805000000
1!
1%
#232810000000
0!
0%
#232815000000
1!
1%
#232820000000
0!
0%
#232825000000
1!
1%
#232830000000
0!
0%
#232835000000
1!
1%
#232840000000
0!
0%
#232845000000
1!
1%
#232850000000
0!
0%
#232855000000
1!
1%
#232860000000
0!
0%
#232865000000
1!
1%
#232870000000
0!
0%
#232875000000
1!
1%
#232880000000
0!
0%
#232885000000
1!
1%
#232890000000
0!
0%
#232895000000
1!
1%
#232900000000
0!
0%
#232905000000
1!
1%
#232910000000
0!
0%
#232915000000
1!
1%
#232920000000
0!
0%
#232925000000
1!
1%
#232930000000
0!
0%
#232935000000
1!
1%
#232940000000
0!
0%
#232945000000
1!
1%
#232950000000
0!
0%
#232955000000
1!
1%
#232960000000
0!
0%
#232965000000
1!
1%
#232970000000
0!
0%
#232975000000
1!
1%
#232980000000
0!
0%
#232985000000
1!
1%
#232990000000
0!
0%
#232995000000
1!
1%
#233000000000
0!
0%
#233005000000
1!
1%
#233010000000
0!
0%
#233015000000
1!
1%
#233020000000
0!
0%
#233025000000
1!
1%
#233030000000
0!
0%
#233035000000
1!
1%
#233040000000
0!
0%
#233045000000
1!
1%
#233050000000
0!
0%
#233055000000
1!
1%
#233060000000
0!
0%
#233065000000
1!
1%
#233070000000
0!
0%
#233075000000
1!
1%
#233080000000
0!
0%
#233085000000
1!
1%
#233090000000
0!
0%
#233095000000
1!
1%
#233100000000
0!
0%
#233105000000
1!
1%
#233110000000
0!
0%
#233115000000
1!
1%
#233120000000
0!
0%
#233125000000
1!
1%
#233130000000
0!
0%
#233135000000
1!
1%
#233140000000
0!
0%
#233145000000
1!
1%
#233150000000
0!
0%
#233155000000
1!
1%
#233160000000
0!
0%
#233165000000
1!
1%
#233170000000
0!
0%
#233175000000
1!
1%
#233180000000
0!
0%
#233185000000
1!
1%
#233190000000
0!
0%
#233195000000
1!
1%
#233200000000
0!
0%
#233205000000
1!
1%
#233210000000
0!
0%
#233215000000
1!
1%
#233220000000
0!
0%
#233225000000
1!
1%
#233230000000
0!
0%
#233235000000
1!
1%
#233240000000
0!
0%
#233245000000
1!
1%
#233250000000
0!
0%
#233255000000
1!
1%
#233260000000
0!
0%
#233265000000
1!
1%
#233270000000
0!
0%
#233275000000
1!
1%
#233280000000
0!
0%
#233285000000
1!
1%
#233290000000
0!
0%
#233295000000
1!
1%
#233300000000
0!
0%
#233305000000
1!
1%
#233310000000
0!
0%
#233315000000
1!
1%
#233320000000
0!
0%
#233325000000
1!
1%
#233330000000
0!
0%
#233335000000
1!
1%
#233340000000
0!
0%
#233345000000
1!
1%
#233350000000
0!
0%
#233355000000
1!
1%
#233360000000
0!
0%
#233365000000
1!
1%
#233370000000
0!
0%
#233375000000
1!
1%
#233380000000
0!
0%
#233385000000
1!
1%
#233390000000
0!
0%
#233395000000
1!
1%
#233400000000
0!
0%
#233405000000
1!
1%
#233410000000
0!
0%
#233415000000
1!
1%
#233420000000
0!
0%
#233425000000
1!
1%
#233430000000
0!
0%
#233435000000
1!
1%
#233440000000
0!
0%
#233445000000
1!
1%
#233450000000
0!
0%
#233455000000
1!
1%
#233460000000
0!
0%
#233465000000
1!
1%
#233470000000
0!
0%
#233475000000
1!
1%
#233480000000
0!
0%
#233485000000
1!
1%
#233490000000
0!
0%
#233495000000
1!
1%
#233500000000
0!
0%
#233505000000
1!
1%
#233510000000
0!
0%
#233515000000
1!
1%
#233520000000
0!
0%
#233525000000
1!
1%
#233530000000
0!
0%
#233535000000
1!
1%
#233540000000
0!
0%
#233545000000
1!
1%
#233550000000
0!
0%
#233555000000
1!
1%
#233560000000
0!
0%
#233565000000
1!
1%
#233570000000
0!
0%
#233575000000
1!
1%
#233580000000
0!
0%
#233585000000
1!
1%
#233590000000
0!
0%
#233595000000
1!
1%
#233600000000
0!
0%
#233605000000
1!
1%
#233610000000
0!
0%
#233615000000
1!
1%
#233620000000
0!
0%
#233625000000
1!
1%
#233630000000
0!
0%
#233635000000
1!
1%
#233640000000
0!
0%
#233645000000
1!
1%
#233650000000
0!
0%
#233655000000
1!
1%
#233660000000
0!
0%
#233665000000
1!
1%
#233670000000
0!
0%
#233675000000
1!
1%
#233680000000
0!
0%
#233685000000
1!
1%
#233690000000
0!
0%
#233695000000
1!
1%
#233700000000
0!
0%
#233705000000
1!
1%
#233710000000
0!
0%
#233715000000
1!
1%
#233720000000
0!
0%
#233725000000
1!
1%
#233730000000
0!
0%
#233735000000
1!
1%
#233740000000
0!
0%
#233745000000
1!
1%
#233750000000
0!
0%
#233755000000
1!
1%
#233760000000
0!
0%
#233765000000
1!
1%
#233770000000
0!
0%
#233775000000
1!
1%
#233780000000
0!
0%
#233785000000
1!
1%
#233790000000
0!
0%
#233795000000
1!
1%
#233800000000
0!
0%
#233805000000
1!
1%
#233810000000
0!
0%
#233815000000
1!
1%
#233820000000
0!
0%
#233825000000
1!
1%
#233830000000
0!
0%
#233835000000
1!
1%
#233840000000
0!
0%
#233845000000
1!
1%
#233850000000
0!
0%
#233855000000
1!
1%
#233860000000
0!
0%
#233865000000
1!
1%
#233870000000
0!
0%
#233875000000
1!
1%
#233880000000
0!
0%
#233885000000
1!
1%
#233890000000
0!
0%
#233895000000
1!
1%
#233900000000
0!
0%
#233905000000
1!
1%
#233910000000
0!
0%
#233915000000
1!
1%
#233920000000
0!
0%
#233925000000
1!
1%
#233930000000
0!
0%
#233935000000
1!
1%
#233940000000
0!
0%
#233945000000
1!
1%
#233950000000
0!
0%
#233955000000
1!
1%
#233960000000
0!
0%
#233965000000
1!
1%
#233970000000
0!
0%
#233975000000
1!
1%
#233980000000
0!
0%
#233985000000
1!
1%
#233990000000
0!
0%
#233995000000
1!
1%
#234000000000
0!
0%
#234005000000
1!
1%
#234010000000
0!
0%
#234015000000
1!
1%
#234020000000
0!
0%
#234025000000
1!
1%
#234030000000
0!
0%
#234035000000
1!
1%
#234040000000
0!
0%
#234045000000
1!
1%
#234050000000
0!
0%
#234055000000
1!
1%
#234060000000
0!
0%
#234065000000
1!
1%
#234070000000
0!
0%
#234075000000
1!
1%
#234080000000
0!
0%
#234085000000
1!
1%
#234090000000
0!
0%
#234095000000
1!
1%
#234100000000
0!
0%
#234105000000
1!
1%
#234110000000
0!
0%
#234115000000
1!
1%
#234120000000
0!
0%
#234125000000
1!
1%
#234130000000
0!
0%
#234135000000
1!
1%
#234140000000
0!
0%
#234145000000
1!
1%
#234150000000
0!
0%
#234155000000
1!
1%
#234160000000
0!
0%
#234165000000
1!
1%
#234170000000
0!
0%
#234175000000
1!
1%
#234180000000
0!
0%
#234185000000
1!
1%
#234190000000
0!
0%
#234195000000
1!
1%
#234200000000
0!
0%
#234205000000
1!
1%
#234210000000
0!
0%
#234215000000
1!
1%
#234220000000
0!
0%
#234225000000
1!
1%
#234230000000
0!
0%
#234235000000
1!
1%
#234240000000
0!
0%
#234245000000
1!
1%
#234250000000
0!
0%
#234255000000
1!
1%
#234260000000
0!
0%
#234265000000
1!
1%
#234270000000
0!
0%
#234275000000
1!
1%
#234280000000
0!
0%
#234285000000
1!
1%
#234290000000
0!
0%
#234295000000
1!
1%
#234300000000
0!
0%
#234305000000
1!
1%
#234310000000
0!
0%
#234315000000
1!
1%
#234320000000
0!
0%
#234325000000
1!
1%
#234330000000
0!
0%
#234335000000
1!
1%
#234340000000
0!
0%
#234345000000
1!
1%
#234350000000
0!
0%
#234355000000
1!
1%
#234360000000
0!
0%
#234365000000
1!
1%
#234370000000
0!
0%
#234375000000
1!
1%
#234380000000
0!
0%
#234385000000
1!
1%
#234390000000
0!
0%
#234395000000
1!
1%
#234400000000
0!
0%
#234405000000
1!
1%
#234410000000
0!
0%
#234415000000
1!
1%
#234420000000
0!
0%
#234425000000
1!
1%
#234430000000
0!
0%
#234435000000
1!
1%
#234440000000
0!
0%
#234445000000
1!
1%
#234450000000
0!
0%
#234455000000
1!
1%
#234460000000
0!
0%
#234465000000
1!
1%
#234470000000
0!
0%
#234475000000
1!
1%
#234480000000
0!
0%
#234485000000
1!
1%
#234490000000
0!
0%
#234495000000
1!
1%
#234500000000
0!
0%
#234505000000
1!
1%
#234510000000
0!
0%
#234515000000
1!
1%
#234520000000
0!
0%
#234525000000
1!
1%
#234530000000
0!
0%
#234535000000
1!
1%
#234540000000
0!
0%
#234545000000
1!
1%
#234550000000
0!
0%
#234555000000
1!
1%
#234560000000
0!
0%
#234565000000
1!
1%
#234570000000
0!
0%
#234575000000
1!
1%
#234580000000
0!
0%
#234585000000
1!
1%
#234590000000
0!
0%
#234595000000
1!
1%
#234600000000
0!
0%
#234605000000
1!
1%
#234610000000
0!
0%
#234615000000
1!
1%
#234620000000
0!
0%
#234625000000
1!
1%
#234630000000
0!
0%
#234635000000
1!
1%
#234640000000
0!
0%
#234645000000
1!
1%
#234650000000
0!
0%
#234655000000
1!
1%
#234660000000
0!
0%
#234665000000
1!
1%
#234670000000
0!
0%
#234675000000
1!
1%
#234680000000
0!
0%
#234685000000
1!
1%
#234690000000
0!
0%
#234695000000
1!
1%
#234700000000
0!
0%
#234705000000
1!
1%
#234710000000
0!
0%
#234715000000
1!
1%
#234720000000
0!
0%
#234725000000
1!
1%
#234730000000
0!
0%
#234735000000
1!
1%
#234740000000
0!
0%
#234745000000
1!
1%
#234750000000
0!
0%
#234755000000
1!
1%
#234760000000
0!
0%
#234765000000
1!
1%
#234770000000
0!
0%
#234775000000
1!
1%
#234780000000
0!
0%
#234785000000
1!
1%
#234790000000
0!
0%
#234795000000
1!
1%
#234800000000
0!
0%
#234805000000
1!
1%
#234810000000
0!
0%
#234815000000
1!
1%
#234820000000
0!
0%
#234825000000
1!
1%
#234830000000
0!
0%
#234835000000
1!
1%
#234840000000
0!
0%
#234845000000
1!
1%
#234850000000
0!
0%
#234855000000
1!
1%
#234860000000
0!
0%
#234865000000
1!
1%
#234870000000
0!
0%
#234875000000
1!
1%
#234880000000
0!
0%
#234885000000
1!
1%
#234890000000
0!
0%
#234895000000
1!
1%
#234900000000
0!
0%
#234905000000
1!
1%
#234910000000
0!
0%
#234915000000
1!
1%
#234920000000
0!
0%
#234925000000
1!
1%
#234930000000
0!
0%
#234935000000
1!
1%
#234940000000
0!
0%
#234945000000
1!
1%
#234950000000
0!
0%
#234955000000
1!
1%
#234960000000
0!
0%
#234965000000
1!
1%
#234970000000
0!
0%
#234975000000
1!
1%
#234980000000
0!
0%
#234985000000
1!
1%
#234990000000
0!
0%
#234995000000
1!
1%
#235000000000
0!
0%
#235005000000
1!
1%
#235010000000
0!
0%
#235015000000
1!
1%
#235020000000
0!
0%
#235025000000
1!
1%
#235030000000
0!
0%
#235035000000
1!
1%
#235040000000
0!
0%
#235045000000
1!
1%
#235050000000
0!
0%
#235055000000
1!
1%
#235060000000
0!
0%
#235065000000
1!
1%
#235070000000
0!
0%
#235075000000
1!
1%
#235080000000
0!
0%
#235085000000
1!
1%
#235090000000
0!
0%
#235095000000
1!
1%
#235100000000
0!
0%
#235105000000
1!
1%
#235110000000
0!
0%
#235115000000
1!
1%
#235120000000
0!
0%
#235125000000
1!
1%
#235130000000
0!
0%
#235135000000
1!
1%
#235140000000
0!
0%
#235145000000
1!
1%
#235150000000
0!
0%
#235155000000
1!
1%
#235160000000
0!
0%
#235165000000
1!
1%
#235170000000
0!
0%
#235175000000
1!
1%
#235180000000
0!
0%
#235185000000
1!
1%
#235190000000
0!
0%
#235195000000
1!
1%
#235200000000
0!
0%
#235205000000
1!
1%
#235210000000
0!
0%
#235215000000
1!
1%
#235220000000
0!
0%
#235225000000
1!
1%
#235230000000
0!
0%
#235235000000
1!
1%
#235240000000
0!
0%
#235245000000
1!
1%
#235250000000
0!
0%
#235255000000
1!
1%
#235260000000
0!
0%
#235265000000
1!
1%
#235270000000
0!
0%
#235275000000
1!
1%
#235280000000
0!
0%
#235285000000
1!
1%
#235290000000
0!
0%
#235295000000
1!
1%
#235300000000
0!
0%
#235305000000
1!
1%
#235310000000
0!
0%
#235315000000
1!
1%
#235320000000
0!
0%
#235325000000
1!
1%
#235330000000
0!
0%
#235335000000
1!
1%
#235340000000
0!
0%
#235345000000
1!
1%
#235350000000
0!
0%
#235355000000
1!
1%
#235360000000
0!
0%
#235365000000
1!
1%
#235370000000
0!
0%
#235375000000
1!
1%
#235380000000
0!
0%
#235385000000
1!
1%
#235390000000
0!
0%
#235395000000
1!
1%
#235400000000
0!
0%
#235405000000
1!
1%
#235410000000
0!
0%
#235415000000
1!
1%
#235420000000
0!
0%
#235425000000
1!
1%
#235430000000
0!
0%
#235435000000
1!
1%
#235440000000
0!
0%
#235445000000
1!
1%
#235450000000
0!
0%
#235455000000
1!
1%
#235460000000
0!
0%
#235465000000
1!
1%
#235470000000
0!
0%
#235475000000
1!
1%
#235480000000
0!
0%
#235485000000
1!
1%
#235490000000
0!
0%
#235495000000
1!
1%
#235500000000
0!
0%
#235505000000
1!
1%
#235510000000
0!
0%
#235515000000
1!
1%
#235520000000
0!
0%
#235525000000
1!
1%
#235530000000
0!
0%
#235535000000
1!
1%
#235540000000
0!
0%
#235545000000
1!
1%
#235550000000
0!
0%
#235555000000
1!
1%
#235560000000
0!
0%
#235565000000
1!
1%
#235570000000
0!
0%
#235575000000
1!
1%
#235580000000
0!
0%
#235585000000
1!
1%
#235590000000
0!
0%
#235595000000
1!
1%
#235600000000
0!
0%
#235605000000
1!
1%
#235610000000
0!
0%
#235615000000
1!
1%
#235620000000
0!
0%
#235625000000
1!
1%
#235630000000
0!
0%
#235635000000
1!
1%
#235640000000
0!
0%
#235645000000
1!
1%
#235650000000
0!
0%
#235655000000
1!
1%
#235660000000
0!
0%
#235665000000
1!
1%
#235670000000
0!
0%
#235675000000
1!
1%
#235680000000
0!
0%
#235685000000
1!
1%
#235690000000
0!
0%
#235695000000
1!
1%
#235700000000
0!
0%
#235705000000
1!
1%
#235710000000
0!
0%
#235715000000
1!
1%
#235720000000
0!
0%
#235725000000
1!
1%
#235730000000
0!
0%
#235735000000
1!
1%
#235740000000
0!
0%
#235745000000
1!
1%
#235750000000
0!
0%
#235755000000
1!
1%
#235760000000
0!
0%
#235765000000
1!
1%
#235770000000
0!
0%
#235775000000
1!
1%
#235780000000
0!
0%
#235785000000
1!
1%
#235790000000
0!
0%
#235795000000
1!
1%
#235800000000
0!
0%
#235805000000
1!
1%
#235810000000
0!
0%
#235815000000
1!
1%
#235820000000
0!
0%
#235825000000
1!
1%
#235830000000
0!
0%
#235835000000
1!
1%
#235840000000
0!
0%
#235845000000
1!
1%
#235850000000
0!
0%
#235855000000
1!
1%
#235860000000
0!
0%
#235865000000
1!
1%
#235870000000
0!
0%
#235875000000
1!
1%
#235880000000
0!
0%
#235885000000
1!
1%
#235890000000
0!
0%
#235895000000
1!
1%
#235900000000
0!
0%
#235905000000
1!
1%
#235910000000
0!
0%
#235915000000
1!
1%
#235920000000
0!
0%
#235925000000
1!
1%
#235930000000
0!
0%
#235935000000
1!
1%
#235940000000
0!
0%
#235945000000
1!
1%
#235950000000
0!
0%
#235955000000
1!
1%
#235960000000
0!
0%
#235965000000
1!
1%
#235970000000
0!
0%
#235975000000
1!
1%
#235980000000
0!
0%
#235985000000
1!
1%
#235990000000
0!
0%
#235995000000
1!
1%
#236000000000
0!
0%
#236005000000
1!
1%
#236010000000
0!
0%
#236015000000
1!
1%
#236020000000
0!
0%
#236025000000
1!
1%
#236030000000
0!
0%
#236035000000
1!
1%
#236040000000
0!
0%
#236045000000
1!
1%
#236050000000
0!
0%
#236055000000
1!
1%
#236060000000
0!
0%
#236065000000
1!
1%
#236070000000
0!
0%
#236075000000
1!
1%
#236080000000
0!
0%
#236085000000
1!
1%
#236090000000
0!
0%
#236095000000
1!
1%
#236100000000
0!
0%
#236105000000
1!
1%
#236110000000
0!
0%
#236115000000
1!
1%
#236120000000
0!
0%
#236125000000
1!
1%
#236130000000
0!
0%
#236135000000
1!
1%
#236140000000
0!
0%
#236145000000
1!
1%
#236150000000
0!
0%
#236155000000
1!
1%
#236160000000
0!
0%
#236165000000
1!
1%
#236170000000
0!
0%
#236175000000
1!
1%
#236180000000
0!
0%
#236185000000
1!
1%
#236190000000
0!
0%
#236195000000
1!
1%
#236200000000
0!
0%
#236205000000
1!
1%
#236210000000
0!
0%
#236215000000
1!
1%
#236220000000
0!
0%
#236225000000
1!
1%
#236230000000
0!
0%
#236235000000
1!
1%
#236240000000
0!
0%
#236245000000
1!
1%
#236250000000
0!
0%
#236255000000
1!
1%
#236260000000
0!
0%
#236265000000
1!
1%
#236270000000
0!
0%
#236275000000
1!
1%
#236280000000
0!
0%
#236285000000
1!
1%
#236290000000
0!
0%
#236295000000
1!
1%
#236300000000
0!
0%
#236305000000
1!
1%
#236310000000
0!
0%
#236315000000
1!
1%
#236320000000
0!
0%
#236325000000
1!
1%
#236330000000
0!
0%
#236335000000
1!
1%
#236340000000
0!
0%
#236345000000
1!
1%
#236350000000
0!
0%
#236355000000
1!
1%
#236360000000
0!
0%
#236365000000
1!
1%
#236370000000
0!
0%
#236375000000
1!
1%
#236380000000
0!
0%
#236385000000
1!
1%
#236390000000
0!
0%
#236395000000
1!
1%
#236400000000
0!
0%
#236405000000
1!
1%
#236410000000
0!
0%
#236415000000
1!
1%
#236420000000
0!
0%
#236425000000
1!
1%
#236430000000
0!
0%
#236435000000
1!
1%
#236440000000
0!
0%
#236445000000
1!
1%
#236450000000
0!
0%
#236455000000
1!
1%
#236460000000
0!
0%
#236465000000
1!
1%
#236470000000
0!
0%
#236475000000
1!
1%
#236480000000
0!
0%
#236485000000
1!
1%
#236490000000
0!
0%
#236495000000
1!
1%
#236500000000
0!
0%
#236505000000
1!
1%
#236510000000
0!
0%
#236515000000
1!
1%
#236520000000
0!
0%
#236525000000
1!
1%
#236530000000
0!
0%
#236535000000
1!
1%
#236540000000
0!
0%
#236545000000
1!
1%
#236550000000
0!
0%
#236555000000
1!
1%
#236560000000
0!
0%
#236565000000
1!
1%
#236570000000
0!
0%
#236575000000
1!
1%
#236580000000
0!
0%
#236585000000
1!
1%
#236590000000
0!
0%
#236595000000
1!
1%
#236600000000
0!
0%
#236605000000
1!
1%
#236610000000
0!
0%
#236615000000
1!
1%
#236620000000
0!
0%
#236625000000
1!
1%
#236630000000
0!
0%
#236635000000
1!
1%
#236640000000
0!
0%
#236645000000
1!
1%
#236650000000
0!
0%
#236655000000
1!
1%
#236660000000
0!
0%
#236665000000
1!
1%
#236670000000
0!
0%
#236675000000
1!
1%
#236680000000
0!
0%
#236685000000
1!
1%
#236690000000
0!
0%
#236695000000
1!
1%
#236700000000
0!
0%
#236705000000
1!
1%
#236710000000
0!
0%
#236715000000
1!
1%
#236720000000
0!
0%
#236725000000
1!
1%
#236730000000
0!
0%
#236735000000
1!
1%
#236740000000
0!
0%
#236745000000
1!
1%
#236750000000
0!
0%
#236755000000
1!
1%
#236760000000
0!
0%
#236765000000
1!
1%
#236770000000
0!
0%
#236775000000
1!
1%
#236780000000
0!
0%
#236785000000
1!
1%
#236790000000
0!
0%
#236795000000
1!
1%
#236800000000
0!
0%
#236805000000
1!
1%
#236810000000
0!
0%
#236815000000
1!
1%
#236820000000
0!
0%
#236825000000
1!
1%
#236830000000
0!
0%
#236835000000
1!
1%
#236840000000
0!
0%
#236845000000
1!
1%
#236850000000
0!
0%
#236855000000
1!
1%
#236860000000
0!
0%
#236865000000
1!
1%
#236870000000
0!
0%
#236875000000
1!
1%
#236880000000
0!
0%
#236885000000
1!
1%
#236890000000
0!
0%
#236895000000
1!
1%
#236900000000
0!
0%
#236905000000
1!
1%
#236910000000
0!
0%
#236915000000
1!
1%
#236920000000
0!
0%
#236925000000
1!
1%
#236930000000
0!
0%
#236935000000
1!
1%
#236940000000
0!
0%
#236945000000
1!
1%
#236950000000
0!
0%
#236955000000
1!
1%
#236960000000
0!
0%
#236965000000
1!
1%
#236970000000
0!
0%
#236975000000
1!
1%
#236980000000
0!
0%
#236985000000
1!
1%
#236990000000
0!
0%
#236995000000
1!
1%
#237000000000
0!
0%
#237005000000
1!
1%
#237010000000
0!
0%
#237015000000
1!
1%
#237020000000
0!
0%
#237025000000
1!
1%
#237030000000
0!
0%
#237035000000
1!
1%
#237040000000
0!
0%
#237045000000
1!
1%
#237050000000
0!
0%
#237055000000
1!
1%
#237060000000
0!
0%
#237065000000
1!
1%
#237070000000
0!
0%
#237075000000
1!
1%
#237080000000
0!
0%
#237085000000
1!
1%
#237090000000
0!
0%
#237095000000
1!
1%
#237100000000
0!
0%
#237105000000
1!
1%
#237110000000
0!
0%
#237115000000
1!
1%
#237120000000
0!
0%
#237125000000
1!
1%
#237130000000
0!
0%
#237135000000
1!
1%
#237140000000
0!
0%
#237145000000
1!
1%
#237150000000
0!
0%
#237155000000
1!
1%
#237160000000
0!
0%
#237165000000
1!
1%
#237170000000
0!
0%
#237175000000
1!
1%
#237180000000
0!
0%
#237185000000
1!
1%
#237190000000
0!
0%
#237195000000
1!
1%
#237200000000
0!
0%
#237205000000
1!
1%
#237210000000
0!
0%
#237215000000
1!
1%
#237220000000
0!
0%
#237225000000
1!
1%
#237230000000
0!
0%
#237235000000
1!
1%
#237240000000
0!
0%
#237245000000
1!
1%
#237250000000
0!
0%
#237255000000
1!
1%
#237260000000
0!
0%
#237265000000
1!
1%
#237270000000
0!
0%
#237275000000
1!
1%
#237280000000
0!
0%
#237285000000
1!
1%
#237290000000
0!
0%
#237295000000
1!
1%
#237300000000
0!
0%
#237305000000
1!
1%
#237310000000
0!
0%
#237315000000
1!
1%
#237320000000
0!
0%
#237325000000
1!
1%
#237330000000
0!
0%
#237335000000
1!
1%
#237340000000
0!
0%
#237345000000
1!
1%
#237350000000
0!
0%
#237355000000
1!
1%
#237360000000
0!
0%
#237365000000
1!
1%
#237370000000
0!
0%
#237375000000
1!
1%
#237380000000
0!
0%
#237385000000
1!
1%
#237390000000
0!
0%
#237395000000
1!
1%
#237400000000
0!
0%
#237405000000
1!
1%
#237410000000
0!
0%
#237415000000
1!
1%
#237420000000
0!
0%
#237425000000
1!
1%
#237430000000
0!
0%
#237435000000
1!
1%
#237440000000
0!
0%
#237445000000
1!
1%
#237450000000
0!
0%
#237455000000
1!
1%
#237460000000
0!
0%
#237465000000
1!
1%
#237470000000
0!
0%
#237475000000
1!
1%
#237480000000
0!
0%
#237485000000
1!
1%
#237490000000
0!
0%
#237495000000
1!
1%
#237500000000
0!
0%
#237505000000
1!
1%
#237510000000
0!
0%
#237515000000
1!
1%
#237520000000
0!
0%
#237525000000
1!
1%
#237530000000
0!
0%
#237535000000
1!
1%
#237540000000
0!
0%
#237545000000
1!
1%
#237550000000
0!
0%
#237555000000
1!
1%
#237560000000
0!
0%
#237565000000
1!
1%
#237570000000
0!
0%
#237575000000
1!
1%
#237580000000
0!
0%
#237585000000
1!
1%
#237590000000
0!
0%
#237595000000
1!
1%
#237600000000
0!
0%
#237605000000
1!
1%
#237610000000
0!
0%
#237615000000
1!
1%
#237620000000
0!
0%
#237625000000
1!
1%
#237630000000
0!
0%
#237635000000
1!
1%
#237640000000
0!
0%
#237645000000
1!
1%
#237650000000
0!
0%
#237655000000
1!
1%
#237660000000
0!
0%
#237665000000
1!
1%
#237670000000
0!
0%
#237675000000
1!
1%
#237680000000
0!
0%
#237685000000
1!
1%
#237690000000
0!
0%
#237695000000
1!
1%
#237700000000
0!
0%
#237705000000
1!
1%
#237710000000
0!
0%
#237715000000
1!
1%
#237720000000
0!
0%
#237725000000
1!
1%
#237730000000
0!
0%
#237735000000
1!
1%
#237740000000
0!
0%
#237745000000
1!
1%
#237750000000
0!
0%
#237755000000
1!
1%
#237760000000
0!
0%
#237765000000
1!
1%
#237770000000
0!
0%
#237775000000
1!
1%
#237780000000
0!
0%
#237785000000
1!
1%
#237790000000
0!
0%
#237795000000
1!
1%
#237800000000
0!
0%
#237805000000
1!
1%
#237810000000
0!
0%
#237815000000
1!
1%
#237820000000
0!
0%
#237825000000
1!
1%
#237830000000
0!
0%
#237835000000
1!
1%
#237840000000
0!
0%
#237845000000
1!
1%
#237850000000
0!
0%
#237855000000
1!
1%
#237860000000
0!
0%
#237865000000
1!
1%
#237870000000
0!
0%
#237875000000
1!
1%
#237880000000
0!
0%
#237885000000
1!
1%
#237890000000
0!
0%
#237895000000
1!
1%
#237900000000
0!
0%
#237905000000
1!
1%
#237910000000
0!
0%
#237915000000
1!
1%
#237920000000
0!
0%
#237925000000
1!
1%
#237930000000
0!
0%
#237935000000
1!
1%
#237940000000
0!
0%
#237945000000
1!
1%
#237950000000
0!
0%
#237955000000
1!
1%
#237960000000
0!
0%
#237965000000
1!
1%
#237970000000
0!
0%
#237975000000
1!
1%
#237980000000
0!
0%
#237985000000
1!
1%
#237990000000
0!
0%
#237995000000
1!
1%
#238000000000
0!
0%
#238005000000
1!
1%
#238010000000
0!
0%
#238015000000
1!
1%
#238020000000
0!
0%
#238025000000
1!
1%
#238030000000
0!
0%
#238035000000
1!
1%
#238040000000
0!
0%
#238045000000
1!
1%
#238050000000
0!
0%
#238055000000
1!
1%
#238060000000
0!
0%
#238065000000
1!
1%
#238070000000
0!
0%
#238075000000
1!
1%
#238080000000
0!
0%
#238085000000
1!
1%
#238090000000
0!
0%
#238095000000
1!
1%
#238100000000
0!
0%
#238105000000
1!
1%
#238110000000
0!
0%
#238115000000
1!
1%
#238120000000
0!
0%
#238125000000
1!
1%
#238130000000
0!
0%
#238135000000
1!
1%
#238140000000
0!
0%
#238145000000
1!
1%
#238150000000
0!
0%
#238155000000
1!
1%
#238160000000
0!
0%
#238165000000
1!
1%
#238170000000
0!
0%
#238175000000
1!
1%
#238180000000
0!
0%
#238185000000
1!
1%
#238190000000
0!
0%
#238195000000
1!
1%
#238200000000
0!
0%
#238205000000
1!
1%
#238210000000
0!
0%
#238215000000
1!
1%
#238220000000
0!
0%
#238225000000
1!
1%
#238230000000
0!
0%
#238235000000
1!
1%
#238240000000
0!
0%
#238245000000
1!
1%
#238250000000
0!
0%
#238255000000
1!
1%
#238260000000
0!
0%
#238265000000
1!
1%
#238270000000
0!
0%
#238275000000
1!
1%
#238280000000
0!
0%
#238285000000
1!
1%
#238290000000
0!
0%
#238295000000
1!
1%
#238300000000
0!
0%
#238305000000
1!
1%
#238310000000
0!
0%
#238315000000
1!
1%
#238320000000
0!
0%
#238325000000
1!
1%
#238330000000
0!
0%
#238335000000
1!
1%
#238340000000
0!
0%
#238345000000
1!
1%
#238350000000
0!
0%
#238355000000
1!
1%
#238360000000
0!
0%
#238365000000
1!
1%
#238370000000
0!
0%
#238375000000
1!
1%
#238380000000
0!
0%
#238385000000
1!
1%
#238390000000
0!
0%
#238395000000
1!
1%
#238400000000
0!
0%
#238405000000
1!
1%
#238410000000
0!
0%
#238415000000
1!
1%
#238420000000
0!
0%
#238425000000
1!
1%
#238430000000
0!
0%
#238435000000
1!
1%
#238440000000
0!
0%
#238445000000
1!
1%
#238450000000
0!
0%
#238455000000
1!
1%
#238460000000
0!
0%
#238465000000
1!
1%
#238470000000
0!
0%
#238475000000
1!
1%
#238480000000
0!
0%
#238485000000
1!
1%
#238490000000
0!
0%
#238495000000
1!
1%
#238500000000
0!
0%
#238505000000
1!
1%
#238510000000
0!
0%
#238515000000
1!
1%
#238520000000
0!
0%
#238525000000
1!
1%
#238530000000
0!
0%
#238535000000
1!
1%
#238540000000
0!
0%
#238545000000
1!
1%
#238550000000
0!
0%
#238555000000
1!
1%
#238560000000
0!
0%
#238565000000
1!
1%
#238570000000
0!
0%
#238575000000
1!
1%
#238580000000
0!
0%
#238585000000
1!
1%
#238590000000
0!
0%
#238595000000
1!
1%
#238600000000
0!
0%
#238605000000
1!
1%
#238610000000
0!
0%
#238615000000
1!
1%
#238620000000
0!
0%
#238625000000
1!
1%
#238630000000
0!
0%
#238635000000
1!
1%
#238640000000
0!
0%
#238645000000
1!
1%
#238650000000
0!
0%
#238655000000
1!
1%
#238660000000
0!
0%
#238665000000
1!
1%
#238670000000
0!
0%
#238675000000
1!
1%
#238680000000
0!
0%
#238685000000
1!
1%
#238690000000
0!
0%
#238695000000
1!
1%
#238700000000
0!
0%
#238705000000
1!
1%
#238710000000
0!
0%
#238715000000
1!
1%
#238720000000
0!
0%
#238725000000
1!
1%
#238730000000
0!
0%
#238735000000
1!
1%
#238740000000
0!
0%
#238745000000
1!
1%
#238750000000
0!
0%
#238755000000
1!
1%
#238760000000
0!
0%
#238765000000
1!
1%
#238770000000
0!
0%
#238775000000
1!
1%
#238780000000
0!
0%
#238785000000
1!
1%
#238790000000
0!
0%
#238795000000
1!
1%
#238800000000
0!
0%
#238805000000
1!
1%
#238810000000
0!
0%
#238815000000
1!
1%
#238820000000
0!
0%
#238825000000
1!
1%
#238830000000
0!
0%
#238835000000
1!
1%
#238840000000
0!
0%
#238845000000
1!
1%
#238850000000
0!
0%
#238855000000
1!
1%
#238860000000
0!
0%
#238865000000
1!
1%
#238870000000
0!
0%
#238875000000
1!
1%
#238880000000
0!
0%
#238885000000
1!
1%
#238890000000
0!
0%
#238895000000
1!
1%
#238900000000
0!
0%
#238905000000
1!
1%
#238910000000
0!
0%
#238915000000
1!
1%
#238920000000
0!
0%
#238925000000
1!
1%
#238930000000
0!
0%
#238935000000
1!
1%
#238940000000
0!
0%
#238945000000
1!
1%
#238950000000
0!
0%
#238955000000
1!
1%
#238960000000
0!
0%
#238965000000
1!
1%
#238970000000
0!
0%
#238975000000
1!
1%
#238980000000
0!
0%
#238985000000
1!
1%
#238990000000
0!
0%
#238995000000
1!
1%
#239000000000
0!
0%
#239005000000
1!
1%
#239010000000
0!
0%
#239015000000
1!
1%
#239020000000
0!
0%
#239025000000
1!
1%
#239030000000
0!
0%
#239035000000
1!
1%
#239040000000
0!
0%
#239045000000
1!
1%
#239050000000
0!
0%
#239055000000
1!
1%
#239060000000
0!
0%
#239065000000
1!
1%
#239070000000
0!
0%
#239075000000
1!
1%
#239080000000
0!
0%
#239085000000
1!
1%
#239090000000
0!
0%
#239095000000
1!
1%
#239100000000
0!
0%
#239105000000
1!
1%
#239110000000
0!
0%
#239115000000
1!
1%
#239120000000
0!
0%
#239125000000
1!
1%
#239130000000
0!
0%
#239135000000
1!
1%
#239140000000
0!
0%
#239145000000
1!
1%
#239150000000
0!
0%
#239155000000
1!
1%
#239160000000
0!
0%
#239165000000
1!
1%
#239170000000
0!
0%
#239175000000
1!
1%
#239180000000
0!
0%
#239185000000
1!
1%
#239190000000
0!
0%
#239195000000
1!
1%
#239200000000
0!
0%
#239205000000
1!
1%
#239210000000
0!
0%
#239215000000
1!
1%
#239220000000
0!
0%
#239225000000
1!
1%
#239230000000
0!
0%
#239235000000
1!
1%
#239240000000
0!
0%
#239245000000
1!
1%
#239250000000
0!
0%
#239255000000
1!
1%
#239260000000
0!
0%
#239265000000
1!
1%
#239270000000
0!
0%
#239275000000
1!
1%
#239280000000
0!
0%
#239285000000
1!
1%
#239290000000
0!
0%
#239295000000
1!
1%
#239300000000
0!
0%
#239305000000
1!
1%
#239310000000
0!
0%
#239315000000
1!
1%
#239320000000
0!
0%
#239325000000
1!
1%
#239330000000
0!
0%
#239335000000
1!
1%
#239340000000
0!
0%
#239345000000
1!
1%
#239350000000
0!
0%
#239355000000
1!
1%
#239360000000
0!
0%
#239365000000
1!
1%
#239370000000
0!
0%
#239375000000
1!
1%
#239380000000
0!
0%
#239385000000
1!
1%
#239390000000
0!
0%
#239395000000
1!
1%
#239400000000
0!
0%
#239405000000
1!
1%
#239410000000
0!
0%
#239415000000
1!
1%
#239420000000
0!
0%
#239425000000
1!
1%
#239430000000
0!
0%
#239435000000
1!
1%
#239440000000
0!
0%
#239445000000
1!
1%
#239450000000
0!
0%
#239455000000
1!
1%
#239460000000
0!
0%
#239465000000
1!
1%
#239470000000
0!
0%
#239475000000
1!
1%
#239480000000
0!
0%
#239485000000
1!
1%
#239490000000
0!
0%
#239495000000
1!
1%
#239500000000
0!
0%
#239505000000
1!
1%
#239510000000
0!
0%
#239515000000
1!
1%
#239520000000
0!
0%
#239525000000
1!
1%
#239530000000
0!
0%
#239535000000
1!
1%
#239540000000
0!
0%
#239545000000
1!
1%
#239550000000
0!
0%
#239555000000
1!
1%
#239560000000
0!
0%
#239565000000
1!
1%
#239570000000
0!
0%
#239575000000
1!
1%
#239580000000
0!
0%
#239585000000
1!
1%
#239590000000
0!
0%
#239595000000
1!
1%
#239600000000
0!
0%
#239605000000
1!
1%
#239610000000
0!
0%
#239615000000
1!
1%
#239620000000
0!
0%
#239625000000
1!
1%
#239630000000
0!
0%
#239635000000
1!
1%
#239640000000
0!
0%
#239645000000
1!
1%
#239650000000
0!
0%
#239655000000
1!
1%
#239660000000
0!
0%
#239665000000
1!
1%
#239670000000
0!
0%
#239675000000
1!
1%
#239680000000
0!
0%
#239685000000
1!
1%
#239690000000
0!
0%
#239695000000
1!
1%
#239700000000
0!
0%
#239705000000
1!
1%
#239710000000
0!
0%
#239715000000
1!
1%
#239720000000
0!
0%
#239725000000
1!
1%
#239730000000
0!
0%
#239735000000
1!
1%
#239740000000
0!
0%
#239745000000
1!
1%
#239750000000
0!
0%
#239755000000
1!
1%
#239760000000
0!
0%
#239765000000
1!
1%
#239770000000
0!
0%
#239775000000
1!
1%
#239780000000
0!
0%
#239785000000
1!
1%
#239790000000
0!
0%
#239795000000
1!
1%
#239800000000
0!
0%
#239805000000
1!
1%
#239810000000
0!
0%
#239815000000
1!
1%
#239820000000
0!
0%
#239825000000
1!
1%
#239830000000
0!
0%
#239835000000
1!
1%
#239840000000
0!
0%
#239845000000
1!
1%
#239850000000
0!
0%
#239855000000
1!
1%
#239860000000
0!
0%
#239865000000
1!
1%
#239870000000
0!
0%
#239875000000
1!
1%
#239880000000
0!
0%
#239885000000
1!
1%
#239890000000
0!
0%
#239895000000
1!
1%
#239900000000
0!
0%
#239905000000
1!
1%
#239910000000
0!
0%
#239915000000
1!
1%
#239920000000
0!
0%
#239925000000
1!
1%
#239930000000
0!
0%
#239935000000
1!
1%
#239940000000
0!
0%
#239945000000
1!
1%
#239950000000
0!
0%
#239955000000
1!
1%
#239960000000
0!
0%
#239965000000
1!
1%
#239970000000
0!
0%
#239975000000
1!
1%
#239980000000
0!
0%
#239985000000
1!
1%
#239990000000
0!
0%
#239995000000
1!
1%
#240000000000
0!
0%
#240005000000
1!
1%
#240010000000
0!
0%
#240015000000
1!
1%
#240020000000
0!
0%
#240025000000
1!
1%
#240030000000
0!
0%
#240035000000
1!
1%
#240040000000
0!
0%
#240045000000
1!
1%
#240050000000
0!
0%
#240055000000
1!
1%
#240060000000
0!
0%
#240065000000
1!
1%
#240070000000
0!
0%
#240075000000
1!
1%
#240080000000
0!
0%
#240085000000
1!
1%
#240090000000
0!
0%
#240095000000
1!
1%
#240100000000
0!
0%
#240105000000
1!
1%
#240110000000
0!
0%
#240115000000
1!
1%
#240120000000
0!
0%
#240125000000
1!
1%
#240130000000
0!
0%
#240135000000
1!
1%
#240140000000
0!
0%
#240145000000
1!
1%
#240150000000
0!
0%
#240155000000
1!
1%
#240160000000
0!
0%
#240165000000
1!
1%
#240170000000
0!
0%
#240175000000
1!
1%
#240180000000
0!
0%
#240185000000
1!
1%
#240190000000
0!
0%
#240195000000
1!
1%
#240200000000
0!
0%
#240205000000
1!
1%
#240210000000
0!
0%
#240215000000
1!
1%
#240220000000
0!
0%
#240225000000
1!
1%
#240230000000
0!
0%
#240235000000
1!
1%
#240240000000
0!
0%
#240245000000
1!
1%
#240250000000
0!
0%
#240255000000
1!
1%
#240260000000
0!
0%
#240265000000
1!
1%
#240270000000
0!
0%
#240275000000
1!
1%
#240280000000
0!
0%
#240285000000
1!
1%
#240290000000
0!
0%
#240295000000
1!
1%
#240300000000
0!
0%
#240305000000
1!
1%
#240310000000
0!
0%
#240315000000
1!
1%
#240320000000
0!
0%
#240325000000
1!
1%
#240330000000
0!
0%
#240335000000
1!
1%
#240340000000
0!
0%
#240345000000
1!
1%
#240350000000
0!
0%
#240355000000
1!
1%
#240360000000
0!
0%
#240365000000
1!
1%
#240370000000
0!
0%
#240375000000
1!
1%
#240380000000
0!
0%
#240385000000
1!
1%
#240390000000
0!
0%
#240395000000
1!
1%
#240400000000
0!
0%
#240405000000
1!
1%
#240410000000
0!
0%
#240415000000
1!
1%
#240420000000
0!
0%
#240425000000
1!
1%
#240430000000
0!
0%
#240435000000
1!
1%
#240440000000
0!
0%
#240445000000
1!
1%
#240450000000
0!
0%
#240455000000
1!
1%
#240460000000
0!
0%
#240465000000
1!
1%
#240470000000
0!
0%
#240475000000
1!
1%
#240480000000
0!
0%
#240485000000
1!
1%
#240490000000
0!
0%
#240495000000
1!
1%
#240500000000
0!
0%
#240505000000
1!
1%
#240510000000
0!
0%
#240515000000
1!
1%
#240520000000
0!
0%
#240525000000
1!
1%
#240530000000
0!
0%
#240535000000
1!
1%
#240540000000
0!
0%
#240545000000
1!
1%
#240550000000
0!
0%
#240555000000
1!
1%
#240560000000
0!
0%
#240565000000
1!
1%
#240570000000
0!
0%
#240575000000
1!
1%
#240580000000
0!
0%
#240585000000
1!
1%
#240590000000
0!
0%
#240595000000
1!
1%
#240600000000
0!
0%
#240605000000
1!
1%
#240610000000
0!
0%
#240615000000
1!
1%
#240620000000
0!
0%
#240625000000
1!
1%
#240630000000
0!
0%
#240635000000
1!
1%
#240640000000
0!
0%
#240645000000
1!
1%
#240650000000
0!
0%
#240655000000
1!
1%
#240660000000
0!
0%
#240665000000
1!
1%
#240670000000
0!
0%
#240675000000
1!
1%
#240680000000
0!
0%
#240685000000
1!
1%
#240690000000
0!
0%
#240695000000
1!
1%
#240700000000
0!
0%
#240705000000
1!
1%
#240710000000
0!
0%
#240715000000
1!
1%
#240720000000
0!
0%
#240725000000
1!
1%
#240730000000
0!
0%
#240735000000
1!
1%
#240740000000
0!
0%
#240745000000
1!
1%
#240750000000
0!
0%
#240755000000
1!
1%
#240760000000
0!
0%
#240765000000
1!
1%
#240770000000
0!
0%
#240775000000
1!
1%
#240780000000
0!
0%
#240785000000
1!
1%
#240790000000
0!
0%
#240795000000
1!
1%
#240800000000
0!
0%
#240805000000
1!
1%
#240810000000
0!
0%
#240815000000
1!
1%
#240820000000
0!
0%
#240825000000
1!
1%
#240830000000
0!
0%
#240835000000
1!
1%
#240840000000
0!
0%
#240845000000
1!
1%
#240850000000
0!
0%
#240855000000
1!
1%
#240860000000
0!
0%
#240865000000
1!
1%
#240870000000
0!
0%
#240875000000
1!
1%
#240880000000
0!
0%
#240885000000
1!
1%
#240890000000
0!
0%
#240895000000
1!
1%
#240900000000
0!
0%
#240905000000
1!
1%
#240910000000
0!
0%
#240915000000
1!
1%
#240920000000
0!
0%
#240925000000
1!
1%
#240930000000
0!
0%
#240935000000
1!
1%
#240940000000
0!
0%
#240945000000
1!
1%
#240950000000
0!
0%
#240955000000
1!
1%
#240960000000
0!
0%
#240965000000
1!
1%
#240970000000
0!
0%
#240975000000
1!
1%
#240980000000
0!
0%
#240985000000
1!
1%
#240990000000
0!
0%
#240995000000
1!
1%
#241000000000
0!
0%
#241005000000
1!
1%
#241010000000
0!
0%
#241015000000
1!
1%
#241020000000
0!
0%
#241025000000
1!
1%
#241030000000
0!
0%
#241035000000
1!
1%
#241040000000
0!
0%
#241045000000
1!
1%
#241050000000
0!
0%
#241055000000
1!
1%
#241060000000
0!
0%
#241065000000
1!
1%
#241070000000
0!
0%
#241075000000
1!
1%
#241080000000
0!
0%
#241085000000
1!
1%
#241090000000
0!
0%
#241095000000
1!
1%
#241100000000
0!
0%
#241105000000
1!
1%
#241110000000
0!
0%
#241115000000
1!
1%
#241120000000
0!
0%
#241125000000
1!
1%
#241130000000
0!
0%
#241135000000
1!
1%
#241140000000
0!
0%
#241145000000
1!
1%
#241150000000
0!
0%
#241155000000
1!
1%
#241160000000
0!
0%
#241165000000
1!
1%
#241170000000
0!
0%
#241175000000
1!
1%
#241180000000
0!
0%
#241185000000
1!
1%
#241190000000
0!
0%
#241195000000
1!
1%
#241200000000
0!
0%
#241205000000
1!
1%
#241210000000
0!
0%
#241215000000
1!
1%
#241220000000
0!
0%
#241225000000
1!
1%
#241230000000
0!
0%
#241235000000
1!
1%
#241240000000
0!
0%
#241245000000
1!
1%
#241250000000
0!
0%
#241255000000
1!
1%
#241260000000
0!
0%
#241265000000
1!
1%
#241270000000
0!
0%
#241275000000
1!
1%
#241280000000
0!
0%
#241285000000
1!
1%
#241290000000
0!
0%
#241295000000
1!
1%
#241300000000
0!
0%
#241305000000
1!
1%
#241310000000
0!
0%
#241315000000
1!
1%
#241320000000
0!
0%
#241325000000
1!
1%
#241330000000
0!
0%
#241335000000
1!
1%
#241340000000
0!
0%
#241345000000
1!
1%
#241350000000
0!
0%
#241355000000
1!
1%
#241360000000
0!
0%
#241365000000
1!
1%
#241370000000
0!
0%
#241375000000
1!
1%
#241380000000
0!
0%
#241385000000
1!
1%
#241390000000
0!
0%
#241395000000
1!
1%
#241400000000
0!
0%
#241405000000
1!
1%
#241410000000
0!
0%
#241415000000
1!
1%
#241420000000
0!
0%
#241425000000
1!
1%
#241430000000
0!
0%
#241435000000
1!
1%
#241440000000
0!
0%
#241445000000
1!
1%
#241450000000
0!
0%
#241455000000
1!
1%
#241460000000
0!
0%
#241465000000
1!
1%
#241470000000
0!
0%
#241475000000
1!
1%
#241480000000
0!
0%
#241485000000
1!
1%
#241490000000
0!
0%
#241495000000
1!
1%
#241500000000
0!
0%
#241505000000
1!
1%
#241510000000
0!
0%
#241515000000
1!
1%
#241520000000
0!
0%
#241525000000
1!
1%
#241530000000
0!
0%
#241535000000
1!
1%
#241540000000
0!
0%
#241545000000
1!
1%
#241550000000
0!
0%
#241555000000
1!
1%
#241560000000
0!
0%
#241565000000
1!
1%
#241570000000
0!
0%
#241575000000
1!
1%
#241580000000
0!
0%
#241585000000
1!
1%
#241590000000
0!
0%
#241595000000
1!
1%
#241600000000
0!
0%
#241605000000
1!
1%
#241610000000
0!
0%
#241615000000
1!
1%
#241620000000
0!
0%
#241625000000
1!
1%
#241630000000
0!
0%
#241635000000
1!
1%
#241640000000
0!
0%
#241645000000
1!
1%
#241650000000
0!
0%
#241655000000
1!
1%
#241660000000
0!
0%
#241665000000
1!
1%
#241670000000
0!
0%
#241675000000
1!
1%
#241680000000
0!
0%
#241685000000
1!
1%
#241690000000
0!
0%
#241695000000
1!
1%
#241700000000
0!
0%
#241705000000
1!
1%
#241710000000
0!
0%
#241715000000
1!
1%
#241720000000
0!
0%
#241725000000
1!
1%
#241730000000
0!
0%
#241735000000
1!
1%
#241740000000
0!
0%
#241745000000
1!
1%
#241750000000
0!
0%
#241755000000
1!
1%
#241760000000
0!
0%
#241765000000
1!
1%
#241770000000
0!
0%
#241775000000
1!
1%
#241780000000
0!
0%
#241785000000
1!
1%
#241790000000
0!
0%
#241795000000
1!
1%
#241800000000
0!
0%
#241805000000
1!
1%
#241810000000
0!
0%
#241815000000
1!
1%
#241820000000
0!
0%
#241825000000
1!
1%
#241830000000
0!
0%
#241835000000
1!
1%
#241840000000
0!
0%
#241845000000
1!
1%
#241850000000
0!
0%
#241855000000
1!
1%
#241860000000
0!
0%
#241865000000
1!
1%
#241870000000
0!
0%
#241875000000
1!
1%
#241880000000
0!
0%
#241885000000
1!
1%
#241890000000
0!
0%
#241895000000
1!
1%
#241900000000
0!
0%
#241905000000
1!
1%
#241910000000
0!
0%
#241915000000
1!
1%
#241920000000
0!
0%
#241925000000
1!
1%
#241930000000
0!
0%
#241935000000
1!
1%
#241940000000
0!
0%
#241945000000
1!
1%
#241950000000
0!
0%
#241955000000
1!
1%
#241960000000
0!
0%
#241965000000
1!
1%
#241970000000
0!
0%
#241975000000
1!
1%
#241980000000
0!
0%
#241985000000
1!
1%
#241990000000
0!
0%
#241995000000
1!
1%
#242000000000
0!
0%
#242005000000
1!
1%
#242010000000
0!
0%
#242015000000
1!
1%
#242020000000
0!
0%
#242025000000
1!
1%
#242030000000
0!
0%
#242035000000
1!
1%
#242040000000
0!
0%
#242045000000
1!
1%
#242050000000
0!
0%
#242055000000
1!
1%
#242060000000
0!
0%
#242065000000
1!
1%
#242070000000
0!
0%
#242075000000
1!
1%
#242080000000
0!
0%
#242085000000
1!
1%
#242090000000
0!
0%
#242095000000
1!
1%
#242100000000
0!
0%
#242105000000
1!
1%
#242110000000
0!
0%
#242115000000
1!
1%
#242120000000
0!
0%
#242125000000
1!
1%
#242130000000
0!
0%
#242135000000
1!
1%
#242140000000
0!
0%
#242145000000
1!
1%
#242150000000
0!
0%
#242155000000
1!
1%
#242160000000
0!
0%
#242165000000
1!
1%
#242170000000
0!
0%
#242175000000
1!
1%
#242180000000
0!
0%
#242185000000
1!
1%
#242190000000
0!
0%
#242195000000
1!
1%
#242200000000
0!
0%
#242205000000
1!
1%
#242210000000
0!
0%
#242215000000
1!
1%
#242220000000
0!
0%
#242225000000
1!
1%
#242230000000
0!
0%
#242235000000
1!
1%
#242240000000
0!
0%
#242245000000
1!
1%
#242250000000
0!
0%
#242255000000
1!
1%
#242260000000
0!
0%
#242265000000
1!
1%
#242270000000
0!
0%
#242275000000
1!
1%
#242280000000
0!
0%
#242285000000
1!
1%
#242290000000
0!
0%
#242295000000
1!
1%
#242300000000
0!
0%
#242305000000
1!
1%
#242310000000
0!
0%
#242315000000
1!
1%
#242320000000
0!
0%
#242325000000
1!
1%
#242330000000
0!
0%
#242335000000
1!
1%
#242340000000
0!
0%
#242345000000
1!
1%
#242350000000
0!
0%
#242355000000
1!
1%
#242360000000
0!
0%
#242365000000
1!
1%
#242370000000
0!
0%
#242375000000
1!
1%
#242380000000
0!
0%
#242385000000
1!
1%
#242390000000
0!
0%
#242395000000
1!
1%
#242400000000
0!
0%
#242405000000
1!
1%
#242410000000
0!
0%
#242415000000
1!
1%
#242420000000
0!
0%
#242425000000
1!
1%
#242430000000
0!
0%
#242435000000
1!
1%
#242440000000
0!
0%
#242445000000
1!
1%
#242450000000
0!
0%
#242455000000
1!
1%
#242460000000
0!
0%
#242465000000
1!
1%
#242470000000
0!
0%
#242475000000
1!
1%
#242480000000
0!
0%
#242485000000
1!
1%
#242490000000
0!
0%
#242495000000
1!
1%
#242500000000
0!
0%
#242505000000
1!
1%
#242510000000
0!
0%
#242515000000
1!
1%
#242520000000
0!
0%
#242525000000
1!
1%
#242530000000
0!
0%
#242535000000
1!
1%
#242540000000
0!
0%
#242545000000
1!
1%
#242550000000
0!
0%
#242555000000
1!
1%
#242560000000
0!
0%
#242565000000
1!
1%
#242570000000
0!
0%
#242575000000
1!
1%
#242580000000
0!
0%
#242585000000
1!
1%
#242590000000
0!
0%
#242595000000
1!
1%
#242600000000
0!
0%
#242605000000
1!
1%
#242610000000
0!
0%
#242615000000
1!
1%
#242620000000
0!
0%
#242625000000
1!
1%
#242630000000
0!
0%
#242635000000
1!
1%
#242640000000
0!
0%
#242645000000
1!
1%
#242650000000
0!
0%
#242655000000
1!
1%
#242660000000
0!
0%
#242665000000
1!
1%
#242670000000
0!
0%
#242675000000
1!
1%
#242680000000
0!
0%
#242685000000
1!
1%
#242690000000
0!
0%
#242695000000
1!
1%
#242700000000
0!
0%
#242705000000
1!
1%
#242710000000
0!
0%
#242715000000
1!
1%
#242720000000
0!
0%
#242725000000
1!
1%
#242730000000
0!
0%
#242735000000
1!
1%
#242740000000
0!
0%
#242745000000
1!
1%
#242750000000
0!
0%
#242755000000
1!
1%
#242760000000
0!
0%
#242765000000
1!
1%
#242770000000
0!
0%
#242775000000
1!
1%
#242780000000
0!
0%
#242785000000
1!
1%
#242790000000
0!
0%
#242795000000
1!
1%
#242800000000
0!
0%
#242805000000
1!
1%
#242810000000
0!
0%
#242815000000
1!
1%
#242820000000
0!
0%
#242825000000
1!
1%
#242830000000
0!
0%
#242835000000
1!
1%
#242840000000
0!
0%
#242845000000
1!
1%
#242850000000
0!
0%
#242855000000
1!
1%
#242860000000
0!
0%
#242865000000
1!
1%
#242870000000
0!
0%
#242875000000
1!
1%
#242880000000
0!
0%
#242885000000
1!
1%
#242890000000
0!
0%
#242895000000
1!
1%
#242900000000
0!
0%
#242905000000
1!
1%
#242910000000
0!
0%
#242915000000
1!
1%
#242920000000
0!
0%
#242925000000
1!
1%
#242930000000
0!
0%
#242935000000
1!
1%
#242940000000
0!
0%
#242945000000
1!
1%
#242950000000
0!
0%
#242955000000
1!
1%
#242960000000
0!
0%
#242965000000
1!
1%
#242970000000
0!
0%
#242975000000
1!
1%
#242980000000
0!
0%
#242985000000
1!
1%
#242990000000
0!
0%
#242995000000
1!
1%
#243000000000
0!
0%
#243005000000
1!
1%
#243010000000
0!
0%
#243015000000
1!
1%
#243020000000
0!
0%
#243025000000
1!
1%
#243030000000
0!
0%
#243035000000
1!
1%
#243040000000
0!
0%
#243045000000
1!
1%
#243050000000
0!
0%
#243055000000
1!
1%
#243060000000
0!
0%
#243065000000
1!
1%
#243070000000
0!
0%
#243075000000
1!
1%
#243080000000
0!
0%
#243085000000
1!
1%
#243090000000
0!
0%
#243095000000
1!
1%
#243100000000
0!
0%
#243105000000
1!
1%
#243110000000
0!
0%
#243115000000
1!
1%
#243120000000
0!
0%
#243125000000
1!
1%
#243130000000
0!
0%
#243135000000
1!
1%
#243140000000
0!
0%
#243145000000
1!
1%
#243150000000
0!
0%
#243155000000
1!
1%
#243160000000
0!
0%
#243165000000
1!
1%
#243170000000
0!
0%
#243175000000
1!
1%
#243180000000
0!
0%
#243185000000
1!
1%
#243190000000
0!
0%
#243195000000
1!
1%
#243200000000
0!
0%
#243205000000
1!
1%
#243210000000
0!
0%
#243215000000
1!
1%
#243220000000
0!
0%
#243225000000
1!
1%
#243230000000
0!
0%
#243235000000
1!
1%
#243240000000
0!
0%
#243245000000
1!
1%
#243250000000
0!
0%
#243255000000
1!
1%
#243260000000
0!
0%
#243265000000
1!
1%
#243270000000
0!
0%
#243275000000
1!
1%
#243280000000
0!
0%
#243285000000
1!
1%
#243290000000
0!
0%
#243295000000
1!
1%
#243300000000
0!
0%
#243305000000
1!
1%
#243310000000
0!
0%
#243315000000
1!
1%
#243320000000
0!
0%
#243325000000
1!
1%
#243330000000
0!
0%
#243335000000
1!
1%
#243340000000
0!
0%
#243345000000
1!
1%
#243350000000
0!
0%
#243355000000
1!
1%
#243360000000
0!
0%
#243365000000
1!
1%
#243370000000
0!
0%
#243375000000
1!
1%
#243380000000
0!
0%
#243385000000
1!
1%
#243390000000
0!
0%
#243395000000
1!
1%
#243400000000
0!
0%
#243405000000
1!
1%
#243410000000
0!
0%
#243415000000
1!
1%
#243420000000
0!
0%
#243425000000
1!
1%
#243430000000
0!
0%
#243435000000
1!
1%
#243440000000
0!
0%
#243445000000
1!
1%
#243450000000
0!
0%
#243455000000
1!
1%
#243460000000
0!
0%
#243465000000
1!
1%
#243470000000
0!
0%
#243475000000
1!
1%
#243480000000
0!
0%
#243485000000
1!
1%
#243490000000
0!
0%
#243495000000
1!
1%
#243500000000
0!
0%
#243505000000
1!
1%
#243510000000
0!
0%
#243515000000
1!
1%
#243520000000
0!
0%
#243525000000
1!
1%
#243530000000
0!
0%
#243535000000
1!
1%
#243540000000
0!
0%
#243545000000
1!
1%
#243550000000
0!
0%
#243555000000
1!
1%
#243560000000
0!
0%
#243565000000
1!
1%
#243570000000
0!
0%
#243575000000
1!
1%
#243580000000
0!
0%
#243585000000
1!
1%
#243590000000
0!
0%
#243595000000
1!
1%
#243600000000
0!
0%
#243605000000
1!
1%
#243610000000
0!
0%
#243615000000
1!
1%
#243620000000
0!
0%
#243625000000
1!
1%
#243630000000
0!
0%
#243635000000
1!
1%
#243640000000
0!
0%
#243645000000
1!
1%
#243650000000
0!
0%
#243655000000
1!
1%
#243660000000
0!
0%
#243665000000
1!
1%
#243670000000
0!
0%
#243675000000
1!
1%
#243680000000
0!
0%
#243685000000
1!
1%
#243690000000
0!
0%
#243695000000
1!
1%
#243700000000
0!
0%
#243705000000
1!
1%
#243710000000
0!
0%
#243715000000
1!
1%
#243720000000
0!
0%
#243725000000
1!
1%
#243730000000
0!
0%
#243735000000
1!
1%
#243740000000
0!
0%
#243745000000
1!
1%
#243750000000
0!
0%
#243755000000
1!
1%
#243760000000
0!
0%
#243765000000
1!
1%
#243770000000
0!
0%
#243775000000
1!
1%
#243780000000
0!
0%
#243785000000
1!
1%
#243790000000
0!
0%
#243795000000
1!
1%
#243800000000
0!
0%
#243805000000
1!
1%
#243810000000
0!
0%
#243815000000
1!
1%
#243820000000
0!
0%
#243825000000
1!
1%
#243830000000
0!
0%
#243835000000
1!
1%
#243840000000
0!
0%
#243845000000
1!
1%
#243850000000
0!
0%
#243855000000
1!
1%
#243860000000
0!
0%
#243865000000
1!
1%
#243870000000
0!
0%
#243875000000
1!
1%
#243880000000
0!
0%
#243885000000
1!
1%
#243890000000
0!
0%
#243895000000
1!
1%
#243900000000
0!
0%
#243905000000
1!
1%
#243910000000
0!
0%
#243915000000
1!
1%
#243920000000
0!
0%
#243925000000
1!
1%
#243930000000
0!
0%
#243935000000
1!
1%
#243940000000
0!
0%
#243945000000
1!
1%
#243950000000
0!
0%
#243955000000
1!
1%
#243960000000
0!
0%
#243965000000
1!
1%
#243970000000
0!
0%
#243975000000
1!
1%
#243980000000
0!
0%
#243985000000
1!
1%
#243990000000
0!
0%
#243995000000
1!
1%
#244000000000
0!
0%
#244005000000
1!
1%
#244010000000
0!
0%
#244015000000
1!
1%
#244020000000
0!
0%
#244025000000
1!
1%
#244030000000
0!
0%
#244035000000
1!
1%
#244040000000
0!
0%
#244045000000
1!
1%
#244050000000
0!
0%
#244055000000
1!
1%
#244060000000
0!
0%
#244065000000
1!
1%
#244070000000
0!
0%
#244075000000
1!
1%
#244080000000
0!
0%
#244085000000
1!
1%
#244090000000
0!
0%
#244095000000
1!
1%
#244100000000
0!
0%
#244105000000
1!
1%
#244110000000
0!
0%
#244115000000
1!
1%
#244120000000
0!
0%
#244125000000
1!
1%
#244130000000
0!
0%
#244135000000
1!
1%
#244140000000
0!
0%
#244145000000
1!
1%
#244150000000
0!
0%
#244155000000
1!
1%
#244160000000
0!
0%
#244165000000
1!
1%
#244170000000
0!
0%
#244175000000
1!
1%
#244180000000
0!
0%
#244185000000
1!
1%
#244190000000
0!
0%
#244195000000
1!
1%
#244200000000
0!
0%
#244205000000
1!
1%
#244210000000
0!
0%
#244215000000
1!
1%
#244220000000
0!
0%
#244225000000
1!
1%
#244230000000
0!
0%
#244235000000
1!
1%
#244240000000
0!
0%
#244245000000
1!
1%
#244250000000
0!
0%
#244255000000
1!
1%
#244260000000
0!
0%
#244265000000
1!
1%
#244270000000
0!
0%
#244275000000
1!
1%
#244280000000
0!
0%
#244285000000
1!
1%
#244290000000
0!
0%
#244295000000
1!
1%
#244300000000
0!
0%
#244305000000
1!
1%
#244310000000
0!
0%
#244315000000
1!
1%
#244320000000
0!
0%
#244325000000
1!
1%
#244330000000
0!
0%
#244335000000
1!
1%
#244340000000
0!
0%
#244345000000
1!
1%
#244350000000
0!
0%
#244355000000
1!
1%
#244360000000
0!
0%
#244365000000
1!
1%
#244370000000
0!
0%
#244375000000
1!
1%
#244380000000
0!
0%
#244385000000
1!
1%
#244390000000
0!
0%
#244395000000
1!
1%
#244400000000
0!
0%
#244405000000
1!
1%
#244410000000
0!
0%
#244415000000
1!
1%
#244420000000
0!
0%
#244425000000
1!
1%
#244430000000
0!
0%
#244435000000
1!
1%
#244440000000
0!
0%
#244445000000
1!
1%
#244450000000
0!
0%
#244455000000
1!
1%
#244460000000
0!
0%
#244465000000
1!
1%
#244470000000
0!
0%
#244475000000
1!
1%
#244480000000
0!
0%
#244485000000
1!
1%
#244490000000
0!
0%
#244495000000
1!
1%
#244500000000
0!
0%
#244505000000
1!
1%
#244510000000
0!
0%
#244515000000
1!
1%
#244520000000
0!
0%
#244525000000
1!
1%
#244530000000
0!
0%
#244535000000
1!
1%
#244540000000
0!
0%
#244545000000
1!
1%
#244550000000
0!
0%
#244555000000
1!
1%
#244560000000
0!
0%
#244565000000
1!
1%
#244570000000
0!
0%
#244575000000
1!
1%
#244580000000
0!
0%
#244585000000
1!
1%
#244590000000
0!
0%
#244595000000
1!
1%
#244600000000
0!
0%
#244605000000
1!
1%
#244610000000
0!
0%
#244615000000
1!
1%
#244620000000
0!
0%
#244625000000
1!
1%
#244630000000
0!
0%
#244635000000
1!
1%
#244640000000
0!
0%
#244645000000
1!
1%
#244650000000
0!
0%
#244655000000
1!
1%
#244660000000
0!
0%
#244665000000
1!
1%
#244670000000
0!
0%
#244675000000
1!
1%
#244680000000
0!
0%
#244685000000
1!
1%
#244690000000
0!
0%
#244695000000
1!
1%
#244700000000
0!
0%
#244705000000
1!
1%
#244710000000
0!
0%
#244715000000
1!
1%
#244720000000
0!
0%
#244725000000
1!
1%
#244730000000
0!
0%
#244735000000
1!
1%
#244740000000
0!
0%
#244745000000
1!
1%
#244750000000
0!
0%
#244755000000
1!
1%
#244760000000
0!
0%
#244765000000
1!
1%
#244770000000
0!
0%
#244775000000
1!
1%
#244780000000
0!
0%
#244785000000
1!
1%
#244790000000
0!
0%
#244795000000
1!
1%
#244800000000
0!
0%
#244805000000
1!
1%
#244810000000
0!
0%
#244815000000
1!
1%
#244820000000
0!
0%
#244825000000
1!
1%
#244830000000
0!
0%
#244835000000
1!
1%
#244840000000
0!
0%
#244845000000
1!
1%
#244850000000
0!
0%
#244855000000
1!
1%
#244860000000
0!
0%
#244865000000
1!
1%
#244870000000
0!
0%
#244875000000
1!
1%
#244880000000
0!
0%
#244885000000
1!
1%
#244890000000
0!
0%
#244895000000
1!
1%
#244900000000
0!
0%
#244905000000
1!
1%
#244910000000
0!
0%
#244915000000
1!
1%
#244920000000
0!
0%
#244925000000
1!
1%
#244930000000
0!
0%
#244935000000
1!
1%
#244940000000
0!
0%
#244945000000
1!
1%
#244950000000
0!
0%
#244955000000
1!
1%
#244960000000
0!
0%
#244965000000
1!
1%
#244970000000
0!
0%
#244975000000
1!
1%
#244980000000
0!
0%
#244985000000
1!
1%
#244990000000
0!
0%
#244995000000
1!
1%
#245000000000
0!
0%
#245005000000
1!
1%
#245010000000
0!
0%
#245015000000
1!
1%
#245020000000
0!
0%
#245025000000
1!
1%
#245030000000
0!
0%
#245035000000
1!
1%
#245040000000
0!
0%
#245045000000
1!
1%
#245050000000
0!
0%
#245055000000
1!
1%
#245060000000
0!
0%
#245065000000
1!
1%
#245070000000
0!
0%
#245075000000
1!
1%
#245080000000
0!
0%
#245085000000
1!
1%
#245090000000
0!
0%
#245095000000
1!
1%
#245100000000
0!
0%
#245105000000
1!
1%
#245110000000
0!
0%
#245115000000
1!
1%
#245120000000
0!
0%
#245125000000
1!
1%
#245130000000
0!
0%
#245135000000
1!
1%
#245140000000
0!
0%
#245145000000
1!
1%
#245150000000
0!
0%
#245155000000
1!
1%
#245160000000
0!
0%
#245165000000
1!
1%
#245170000000
0!
0%
#245175000000
1!
1%
#245180000000
0!
0%
#245185000000
1!
1%
#245190000000
0!
0%
#245195000000
1!
1%
#245200000000
0!
0%
#245205000000
1!
1%
#245210000000
0!
0%
#245215000000
1!
1%
#245220000000
0!
0%
#245225000000
1!
1%
#245230000000
0!
0%
#245235000000
1!
1%
#245240000000
0!
0%
#245245000000
1!
1%
#245250000000
0!
0%
#245255000000
1!
1%
#245260000000
0!
0%
#245265000000
1!
1%
#245270000000
0!
0%
#245275000000
1!
1%
#245280000000
0!
0%
#245285000000
1!
1%
#245290000000
0!
0%
#245295000000
1!
1%
#245300000000
0!
0%
#245305000000
1!
1%
#245310000000
0!
0%
#245315000000
1!
1%
#245320000000
0!
0%
#245325000000
1!
1%
#245330000000
0!
0%
#245335000000
1!
1%
#245340000000
0!
0%
#245345000000
1!
1%
#245350000000
0!
0%
#245355000000
1!
1%
#245360000000
0!
0%
#245365000000
1!
1%
#245370000000
0!
0%
#245375000000
1!
1%
#245380000000
0!
0%
#245385000000
1!
1%
#245390000000
0!
0%
#245395000000
1!
1%
#245400000000
0!
0%
#245405000000
1!
1%
#245410000000
0!
0%
#245415000000
1!
1%
#245420000000
0!
0%
#245425000000
1!
1%
#245430000000
0!
0%
#245435000000
1!
1%
#245440000000
0!
0%
#245445000000
1!
1%
#245450000000
0!
0%
#245455000000
1!
1%
#245460000000
0!
0%
#245465000000
1!
1%
#245470000000
0!
0%
#245475000000
1!
1%
#245480000000
0!
0%
#245485000000
1!
1%
#245490000000
0!
0%
#245495000000
1!
1%
#245500000000
0!
0%
#245505000000
1!
1%
#245510000000
0!
0%
#245515000000
1!
1%
#245520000000
0!
0%
#245525000000
1!
1%
#245530000000
0!
0%
#245535000000
1!
1%
#245540000000
0!
0%
#245545000000
1!
1%
#245550000000
0!
0%
#245555000000
1!
1%
#245560000000
0!
0%
#245565000000
1!
1%
#245570000000
0!
0%
#245575000000
1!
1%
#245580000000
0!
0%
#245585000000
1!
1%
#245590000000
0!
0%
#245595000000
1!
1%
#245600000000
0!
0%
#245605000000
1!
1%
#245610000000
0!
0%
#245615000000
1!
1%
#245620000000
0!
0%
#245625000000
1!
1%
#245630000000
0!
0%
#245635000000
1!
1%
#245640000000
0!
0%
#245645000000
1!
1%
#245650000000
0!
0%
#245655000000
1!
1%
#245660000000
0!
0%
#245665000000
1!
1%
#245670000000
0!
0%
#245675000000
1!
1%
#245680000000
0!
0%
#245685000000
1!
1%
#245690000000
0!
0%
#245695000000
1!
1%
#245700000000
0!
0%
#245705000000
1!
1%
#245710000000
0!
0%
#245715000000
1!
1%
#245720000000
0!
0%
#245725000000
1!
1%
#245730000000
0!
0%
#245735000000
1!
1%
#245740000000
0!
0%
#245745000000
1!
1%
#245750000000
0!
0%
#245755000000
1!
1%
#245760000000
0!
0%
#245765000000
1!
1%
#245770000000
0!
0%
#245775000000
1!
1%
#245780000000
0!
0%
#245785000000
1!
1%
#245790000000
0!
0%
#245795000000
1!
1%
#245800000000
0!
0%
#245805000000
1!
1%
#245810000000
0!
0%
#245815000000
1!
1%
#245820000000
0!
0%
#245825000000
1!
1%
#245830000000
0!
0%
#245835000000
1!
1%
#245840000000
0!
0%
#245845000000
1!
1%
#245850000000
0!
0%
#245855000000
1!
1%
#245860000000
0!
0%
#245865000000
1!
1%
#245870000000
0!
0%
#245875000000
1!
1%
#245880000000
0!
0%
#245885000000
1!
1%
#245890000000
0!
0%
#245895000000
1!
1%
#245900000000
0!
0%
#245905000000
1!
1%
#245910000000
0!
0%
#245915000000
1!
1%
#245920000000
0!
0%
#245925000000
1!
1%
#245930000000
0!
0%
#245935000000
1!
1%
#245940000000
0!
0%
#245945000000
1!
1%
#245950000000
0!
0%
#245955000000
1!
1%
#245960000000
0!
0%
#245965000000
1!
1%
#245970000000
0!
0%
#245975000000
1!
1%
#245980000000
0!
0%
#245985000000
1!
1%
#245990000000
0!
0%
#245995000000
1!
1%
#246000000000
0!
0%
#246005000000
1!
1%
#246010000000
0!
0%
#246015000000
1!
1%
#246020000000
0!
0%
#246025000000
1!
1%
#246030000000
0!
0%
#246035000000
1!
1%
#246040000000
0!
0%
#246045000000
1!
1%
#246050000000
0!
0%
#246055000000
1!
1%
#246060000000
0!
0%
#246065000000
1!
1%
#246070000000
0!
0%
#246075000000
1!
1%
#246080000000
0!
0%
#246085000000
1!
1%
#246090000000
0!
0%
#246095000000
1!
1%
#246100000000
0!
0%
#246105000000
1!
1%
#246110000000
0!
0%
#246115000000
1!
1%
#246120000000
0!
0%
#246125000000
1!
1%
#246130000000
0!
0%
#246135000000
1!
1%
#246140000000
0!
0%
#246145000000
1!
1%
#246150000000
0!
0%
#246155000000
1!
1%
#246160000000
0!
0%
#246165000000
1!
1%
#246170000000
0!
0%
#246175000000
1!
1%
#246180000000
0!
0%
#246185000000
1!
1%
#246190000000
0!
0%
#246195000000
1!
1%
#246200000000
0!
0%
#246205000000
1!
1%
#246210000000
0!
0%
#246215000000
1!
1%
#246220000000
0!
0%
#246225000000
1!
1%
#246230000000
0!
0%
#246235000000
1!
1%
#246240000000
0!
0%
#246245000000
1!
1%
#246250000000
0!
0%
#246255000000
1!
1%
#246260000000
0!
0%
#246265000000
1!
1%
#246270000000
0!
0%
#246275000000
1!
1%
#246280000000
0!
0%
#246285000000
1!
1%
#246290000000
0!
0%
#246295000000
1!
1%
#246300000000
0!
0%
#246305000000
1!
1%
#246310000000
0!
0%
#246315000000
1!
1%
#246320000000
0!
0%
#246325000000
1!
1%
#246330000000
0!
0%
#246335000000
1!
1%
#246340000000
0!
0%
#246345000000
1!
1%
#246350000000
0!
0%
#246355000000
1!
1%
#246360000000
0!
0%
#246365000000
1!
1%
#246370000000
0!
0%
#246375000000
1!
1%
#246380000000
0!
0%
#246385000000
1!
1%
#246390000000
0!
0%
#246395000000
1!
1%
#246400000000
0!
0%
#246405000000
1!
1%
#246410000000
0!
0%
#246415000000
1!
1%
#246420000000
0!
0%
#246425000000
1!
1%
#246430000000
0!
0%
#246435000000
1!
1%
#246440000000
0!
0%
#246445000000
1!
1%
#246450000000
0!
0%
#246455000000
1!
1%
#246460000000
0!
0%
#246465000000
1!
1%
#246470000000
0!
0%
#246475000000
1!
1%
#246480000000
0!
0%
#246485000000
1!
1%
#246490000000
0!
0%
#246495000000
1!
1%
#246500000000
0!
0%
#246505000000
1!
1%
#246510000000
0!
0%
#246515000000
1!
1%
#246520000000
0!
0%
#246525000000
1!
1%
#246530000000
0!
0%
#246535000000
1!
1%
#246540000000
0!
0%
#246545000000
1!
1%
#246550000000
0!
0%
#246555000000
1!
1%
#246560000000
0!
0%
#246565000000
1!
1%
#246570000000
0!
0%
#246575000000
1!
1%
#246580000000
0!
0%
#246585000000
1!
1%
#246590000000
0!
0%
#246595000000
1!
1%
#246600000000
0!
0%
#246605000000
1!
1%
#246610000000
0!
0%
#246615000000
1!
1%
#246620000000
0!
0%
#246625000000
1!
1%
#246630000000
0!
0%
#246635000000
1!
1%
#246640000000
0!
0%
#246645000000
1!
1%
#246650000000
0!
0%
#246655000000
1!
1%
#246660000000
0!
0%
#246665000000
1!
1%
#246670000000
0!
0%
#246675000000
1!
1%
#246680000000
0!
0%
#246685000000
1!
1%
#246690000000
0!
0%
#246695000000
1!
1%
#246700000000
0!
0%
#246705000000
1!
1%
#246710000000
0!
0%
#246715000000
1!
1%
#246720000000
0!
0%
#246725000000
1!
1%
#246730000000
0!
0%
#246735000000
1!
1%
#246740000000
0!
0%
#246745000000
1!
1%
#246750000000
0!
0%
#246755000000
1!
1%
#246760000000
0!
0%
#246765000000
1!
1%
#246770000000
0!
0%
#246775000000
1!
1%
#246780000000
0!
0%
#246785000000
1!
1%
#246790000000
0!
0%
#246795000000
1!
1%
#246800000000
0!
0%
#246805000000
1!
1%
#246810000000
0!
0%
#246815000000
1!
1%
#246820000000
0!
0%
#246825000000
1!
1%
#246830000000
0!
0%
#246835000000
1!
1%
#246840000000
0!
0%
#246845000000
1!
1%
#246850000000
0!
0%
#246855000000
1!
1%
#246860000000
0!
0%
#246865000000
1!
1%
#246870000000
0!
0%
#246875000000
1!
1%
#246880000000
0!
0%
#246885000000
1!
1%
#246890000000
0!
0%
#246895000000
1!
1%
#246900000000
0!
0%
#246905000000
1!
1%
#246910000000
0!
0%
#246915000000
1!
1%
#246920000000
0!
0%
#246925000000
1!
1%
#246930000000
0!
0%
#246935000000
1!
1%
#246940000000
0!
0%
#246945000000
1!
1%
#246950000000
0!
0%
#246955000000
1!
1%
#246960000000
0!
0%
#246965000000
1!
1%
#246970000000
0!
0%
#246975000000
1!
1%
#246980000000
0!
0%
#246985000000
1!
1%
#246990000000
0!
0%
#246995000000
1!
1%
#247000000000
0!
0%
#247005000000
1!
1%
#247010000000
0!
0%
#247015000000
1!
1%
#247020000000
0!
0%
#247025000000
1!
1%
#247030000000
0!
0%
#247035000000
1!
1%
#247040000000
0!
0%
#247045000000
1!
1%
#247050000000
0!
0%
#247055000000
1!
1%
#247060000000
0!
0%
#247065000000
1!
1%
#247070000000
0!
0%
#247075000000
1!
1%
#247080000000
0!
0%
#247085000000
1!
1%
#247090000000
0!
0%
#247095000000
1!
1%
#247100000000
0!
0%
#247105000000
1!
1%
#247110000000
0!
0%
#247115000000
1!
1%
#247120000000
0!
0%
#247125000000
1!
1%
#247130000000
0!
0%
#247135000000
1!
1%
#247140000000
0!
0%
#247145000000
1!
1%
#247150000000
0!
0%
#247155000000
1!
1%
#247160000000
0!
0%
#247165000000
1!
1%
#247170000000
0!
0%
#247175000000
1!
1%
#247180000000
0!
0%
#247185000000
1!
1%
#247190000000
0!
0%
#247195000000
1!
1%
#247200000000
0!
0%
#247205000000
1!
1%
#247210000000
0!
0%
#247215000000
1!
1%
#247220000000
0!
0%
#247225000000
1!
1%
#247230000000
0!
0%
#247235000000
1!
1%
#247240000000
0!
0%
#247245000000
1!
1%
#247250000000
0!
0%
#247255000000
1!
1%
#247260000000
0!
0%
#247265000000
1!
1%
#247270000000
0!
0%
#247275000000
1!
1%
#247280000000
0!
0%
#247285000000
1!
1%
#247290000000
0!
0%
#247295000000
1!
1%
#247300000000
0!
0%
#247305000000
1!
1%
#247310000000
0!
0%
#247315000000
1!
1%
#247320000000
0!
0%
#247325000000
1!
1%
#247330000000
0!
0%
#247335000000
1!
1%
#247340000000
0!
0%
#247345000000
1!
1%
#247350000000
0!
0%
#247355000000
1!
1%
#247360000000
0!
0%
#247365000000
1!
1%
#247370000000
0!
0%
#247375000000
1!
1%
#247380000000
0!
0%
#247385000000
1!
1%
#247390000000
0!
0%
#247395000000
1!
1%
#247400000000
0!
0%
#247405000000
1!
1%
#247410000000
0!
0%
#247415000000
1!
1%
#247420000000
0!
0%
#247425000000
1!
1%
#247430000000
0!
0%
#247435000000
1!
1%
#247440000000
0!
0%
#247445000000
1!
1%
#247450000000
0!
0%
#247455000000
1!
1%
#247460000000
0!
0%
#247465000000
1!
1%
#247470000000
0!
0%
#247475000000
1!
1%
#247480000000
0!
0%
#247485000000
1!
1%
#247490000000
0!
0%
#247495000000
1!
1%
#247500000000
0!
0%
#247505000000
1!
1%
#247510000000
0!
0%
#247515000000
1!
1%
#247520000000
0!
0%
#247525000000
1!
1%
#247530000000
0!
0%
#247535000000
1!
1%
#247540000000
0!
0%
#247545000000
1!
1%
#247550000000
0!
0%
#247555000000
1!
1%
#247560000000
0!
0%
#247565000000
1!
1%
#247570000000
0!
0%
#247575000000
1!
1%
#247580000000
0!
0%
#247585000000
1!
1%
#247590000000
0!
0%
#247595000000
1!
1%
#247600000000
0!
0%
#247605000000
1!
1%
#247610000000
0!
0%
#247615000000
1!
1%
#247620000000
0!
0%
#247625000000
1!
1%
#247630000000
0!
0%
#247635000000
1!
1%
#247640000000
0!
0%
#247645000000
1!
1%
#247650000000
0!
0%
#247655000000
1!
1%
#247660000000
0!
0%
#247665000000
1!
1%
#247670000000
0!
0%
#247675000000
1!
1%
#247680000000
0!
0%
#247685000000
1!
1%
#247690000000
0!
0%
#247695000000
1!
1%
#247700000000
0!
0%
#247705000000
1!
1%
#247710000000
0!
0%
#247715000000
1!
1%
#247720000000
0!
0%
#247725000000
1!
1%
#247730000000
0!
0%
#247735000000
1!
1%
#247740000000
0!
0%
#247745000000
1!
1%
#247750000000
0!
0%
#247755000000
1!
1%
#247760000000
0!
0%
#247765000000
1!
1%
#247770000000
0!
0%
#247775000000
1!
1%
#247780000000
0!
0%
#247785000000
1!
1%
#247790000000
0!
0%
#247795000000
1!
1%
#247800000000
0!
0%
#247805000000
1!
1%
#247810000000
0!
0%
#247815000000
1!
1%
#247820000000
0!
0%
#247825000000
1!
1%
#247830000000
0!
0%
#247835000000
1!
1%
#247840000000
0!
0%
#247845000000
1!
1%
#247850000000
0!
0%
#247855000000
1!
1%
#247860000000
0!
0%
#247865000000
1!
1%
#247870000000
0!
0%
#247875000000
1!
1%
#247880000000
0!
0%
#247885000000
1!
1%
#247890000000
0!
0%
#247895000000
1!
1%
#247900000000
0!
0%
#247905000000
1!
1%
#247910000000
0!
0%
#247915000000
1!
1%
#247920000000
0!
0%
#247925000000
1!
1%
#247930000000
0!
0%
#247935000000
1!
1%
#247940000000
0!
0%
#247945000000
1!
1%
#247950000000
0!
0%
#247955000000
1!
1%
#247960000000
0!
0%
#247965000000
1!
1%
#247970000000
0!
0%
#247975000000
1!
1%
#247980000000
0!
0%
#247985000000
1!
1%
#247990000000
0!
0%
#247995000000
1!
1%
#248000000000
0!
0%
#248005000000
1!
1%
#248010000000
0!
0%
#248015000000
1!
1%
#248020000000
0!
0%
#248025000000
1!
1%
#248030000000
0!
0%
#248035000000
1!
1%
#248040000000
0!
0%
#248045000000
1!
1%
#248050000000
0!
0%
#248055000000
1!
1%
#248060000000
0!
0%
#248065000000
1!
1%
#248070000000
0!
0%
#248075000000
1!
1%
#248080000000
0!
0%
#248085000000
1!
1%
#248090000000
0!
0%
#248095000000
1!
1%
#248100000000
0!
0%
#248105000000
1!
1%
#248110000000
0!
0%
#248115000000
1!
1%
#248120000000
0!
0%
#248125000000
1!
1%
#248130000000
0!
0%
#248135000000
1!
1%
#248140000000
0!
0%
#248145000000
1!
1%
#248150000000
0!
0%
#248155000000
1!
1%
#248160000000
0!
0%
#248165000000
1!
1%
#248170000000
0!
0%
#248175000000
1!
1%
#248180000000
0!
0%
#248185000000
1!
1%
#248190000000
0!
0%
#248195000000
1!
1%
#248200000000
0!
0%
#248205000000
1!
1%
#248210000000
0!
0%
#248215000000
1!
1%
#248220000000
0!
0%
#248225000000
1!
1%
#248230000000
0!
0%
#248235000000
1!
1%
#248240000000
0!
0%
#248245000000
1!
1%
#248250000000
0!
0%
#248255000000
1!
1%
#248260000000
0!
0%
#248265000000
1!
1%
#248270000000
0!
0%
#248275000000
1!
1%
#248280000000
0!
0%
#248285000000
1!
1%
#248290000000
0!
0%
#248295000000
1!
1%
#248300000000
0!
0%
#248305000000
1!
1%
#248310000000
0!
0%
#248315000000
1!
1%
#248320000000
0!
0%
#248325000000
1!
1%
#248330000000
0!
0%
#248335000000
1!
1%
#248340000000
0!
0%
#248345000000
1!
1%
#248350000000
0!
0%
#248355000000
1!
1%
#248360000000
0!
0%
#248365000000
1!
1%
#248370000000
0!
0%
#248375000000
1!
1%
#248380000000
0!
0%
#248385000000
1!
1%
#248390000000
0!
0%
#248395000000
1!
1%
#248400000000
0!
0%
#248405000000
1!
1%
#248410000000
0!
0%
#248415000000
1!
1%
#248420000000
0!
0%
#248425000000
1!
1%
#248430000000
0!
0%
#248435000000
1!
1%
#248440000000
0!
0%
#248445000000
1!
1%
#248450000000
0!
0%
#248455000000
1!
1%
#248460000000
0!
0%
#248465000000
1!
1%
#248470000000
0!
0%
#248475000000
1!
1%
#248480000000
0!
0%
#248485000000
1!
1%
#248490000000
0!
0%
#248495000000
1!
1%
#248500000000
0!
0%
#248505000000
1!
1%
#248510000000
0!
0%
#248515000000
1!
1%
#248520000000
0!
0%
#248525000000
1!
1%
#248530000000
0!
0%
#248535000000
1!
1%
#248540000000
0!
0%
#248545000000
1!
1%
#248550000000
0!
0%
#248555000000
1!
1%
#248560000000
0!
0%
#248565000000
1!
1%
#248570000000
0!
0%
#248575000000
1!
1%
#248580000000
0!
0%
#248585000000
1!
1%
#248590000000
0!
0%
#248595000000
1!
1%
#248600000000
0!
0%
#248605000000
1!
1%
#248610000000
0!
0%
#248615000000
1!
1%
#248620000000
0!
0%
#248625000000
1!
1%
#248630000000
0!
0%
#248635000000
1!
1%
#248640000000
0!
0%
#248645000000
1!
1%
#248650000000
0!
0%
#248655000000
1!
1%
#248660000000
0!
0%
#248665000000
1!
1%
#248670000000
0!
0%
#248675000000
1!
1%
#248680000000
0!
0%
#248685000000
1!
1%
#248690000000
0!
0%
#248695000000
1!
1%
#248700000000
0!
0%
#248705000000
1!
1%
#248710000000
0!
0%
#248715000000
1!
1%
#248720000000
0!
0%
#248725000000
1!
1%
#248730000000
0!
0%
#248735000000
1!
1%
#248740000000
0!
0%
#248745000000
1!
1%
#248750000000
0!
0%
#248755000000
1!
1%
#248760000000
0!
0%
#248765000000
1!
1%
#248770000000
0!
0%
#248775000000
1!
1%
#248780000000
0!
0%
#248785000000
1!
1%
#248790000000
0!
0%
#248795000000
1!
1%
#248800000000
0!
0%
#248805000000
1!
1%
#248810000000
0!
0%
#248815000000
1!
1%
#248820000000
0!
0%
#248825000000
1!
1%
#248830000000
0!
0%
#248835000000
1!
1%
#248840000000
0!
0%
#248845000000
1!
1%
#248850000000
0!
0%
#248855000000
1!
1%
#248860000000
0!
0%
#248865000000
1!
1%
#248870000000
0!
0%
#248875000000
1!
1%
#248880000000
0!
0%
#248885000000
1!
1%
#248890000000
0!
0%
#248895000000
1!
1%
#248900000000
0!
0%
#248905000000
1!
1%
#248910000000
0!
0%
#248915000000
1!
1%
#248920000000
0!
0%
#248925000000
1!
1%
#248930000000
0!
0%
#248935000000
1!
1%
#248940000000
0!
0%
#248945000000
1!
1%
#248950000000
0!
0%
#248955000000
1!
1%
#248960000000
0!
0%
#248965000000
1!
1%
#248970000000
0!
0%
#248975000000
1!
1%
#248980000000
0!
0%
#248985000000
1!
1%
#248990000000
0!
0%
#248995000000
1!
1%
#249000000000
0!
0%
#249005000000
1!
1%
#249010000000
0!
0%
#249015000000
1!
1%
#249020000000
0!
0%
#249025000000
1!
1%
#249030000000
0!
0%
#249035000000
1!
1%
#249040000000
0!
0%
#249045000000
1!
1%
#249050000000
0!
0%
#249055000000
1!
1%
#249060000000
0!
0%
#249065000000
1!
1%
#249070000000
0!
0%
#249075000000
1!
1%
#249080000000
0!
0%
#249085000000
1!
1%
#249090000000
0!
0%
#249095000000
1!
1%
#249100000000
0!
0%
#249105000000
1!
1%
#249110000000
0!
0%
#249115000000
1!
1%
#249120000000
0!
0%
#249125000000
1!
1%
#249130000000
0!
0%
#249135000000
1!
1%
#249140000000
0!
0%
#249145000000
1!
1%
#249150000000
0!
0%
#249155000000
1!
1%
#249160000000
0!
0%
#249165000000
1!
1%
#249170000000
0!
0%
#249175000000
1!
1%
#249180000000
0!
0%
#249185000000
1!
1%
#249190000000
0!
0%
#249195000000
1!
1%
#249200000000
0!
0%
#249205000000
1!
1%
#249210000000
0!
0%
#249215000000
1!
1%
#249220000000
0!
0%
#249225000000
1!
1%
#249230000000
0!
0%
#249235000000
1!
1%
#249240000000
0!
0%
#249245000000
1!
1%
#249250000000
0!
0%
#249255000000
1!
1%
#249260000000
0!
0%
#249265000000
1!
1%
#249270000000
0!
0%
#249275000000
1!
1%
#249280000000
0!
0%
#249285000000
1!
1%
#249290000000
0!
0%
#249295000000
1!
1%
#249300000000
0!
0%
#249305000000
1!
1%
#249310000000
0!
0%
#249315000000
1!
1%
#249320000000
0!
0%
#249325000000
1!
1%
#249330000000
0!
0%
#249335000000
1!
1%
#249340000000
0!
0%
#249345000000
1!
1%
#249350000000
0!
0%
#249355000000
1!
1%
#249360000000
0!
0%
#249365000000
1!
1%
#249370000000
0!
0%
#249375000000
1!
1%
#249380000000
0!
0%
#249385000000
1!
1%
#249390000000
0!
0%
#249395000000
1!
1%
#249400000000
0!
0%
#249405000000
1!
1%
#249410000000
0!
0%
#249415000000
1!
1%
#249420000000
0!
0%
#249425000000
1!
1%
#249430000000
0!
0%
#249435000000
1!
1%
#249440000000
0!
0%
#249445000000
1!
1%
#249450000000
0!
0%
#249455000000
1!
1%
#249460000000
0!
0%
#249465000000
1!
1%
#249470000000
0!
0%
#249475000000
1!
1%
#249480000000
0!
0%
#249485000000
1!
1%
#249490000000
0!
0%
#249495000000
1!
1%
#249500000000
0!
0%
#249505000000
1!
1%
#249510000000
0!
0%
#249515000000
1!
1%
#249520000000
0!
0%
#249525000000
1!
1%
#249530000000
0!
0%
#249535000000
1!
1%
#249540000000
0!
0%
#249545000000
1!
1%
#249550000000
0!
0%
#249555000000
1!
1%
#249560000000
0!
0%
#249565000000
1!
1%
#249570000000
0!
0%
#249575000000
1!
1%
#249580000000
0!
0%
#249585000000
1!
1%
#249590000000
0!
0%
#249595000000
1!
1%
#249600000000
0!
0%
#249605000000
1!
1%
#249610000000
0!
0%
#249615000000
1!
1%
#249620000000
0!
0%
#249625000000
1!
1%
#249630000000
0!
0%
#249635000000
1!
1%
#249640000000
0!
0%
#249645000000
1!
1%
#249650000000
0!
0%
#249655000000
1!
1%
#249660000000
0!
0%
#249665000000
1!
1%
#249670000000
0!
0%
#249675000000
1!
1%
#249680000000
0!
0%
#249685000000
1!
1%
#249690000000
0!
0%
#249695000000
1!
1%
#249700000000
0!
0%
#249705000000
1!
1%
#249710000000
0!
0%
#249715000000
1!
1%
#249720000000
0!
0%
#249725000000
1!
1%
#249730000000
0!
0%
#249735000000
1!
1%
#249740000000
0!
0%
#249745000000
1!
1%
#249750000000
0!
0%
#249755000000
1!
1%
#249760000000
0!
0%
#249765000000
1!
1%
#249770000000
0!
0%
#249775000000
1!
1%
#249780000000
0!
0%
#249785000000
1!
1%
#249790000000
0!
0%
#249795000000
1!
1%
#249800000000
0!
0%
#249805000000
1!
1%
#249810000000
0!
0%
#249815000000
1!
1%
#249820000000
0!
0%
#249825000000
1!
1%
#249830000000
0!
0%
#249835000000
1!
1%
#249840000000
0!
0%
#249845000000
1!
1%
#249850000000
0!
0%
#249855000000
1!
1%
#249860000000
0!
0%
#249865000000
1!
1%
#249870000000
0!
0%
#249875000000
1!
1%
#249880000000
0!
0%
#249885000000
1!
1%
#249890000000
0!
0%
#249895000000
1!
1%
#249900000000
0!
0%
#249905000000
1!
1%
#249910000000
0!
0%
#249915000000
1!
1%
#249920000000
0!
0%
#249925000000
1!
1%
#249930000000
0!
0%
#249935000000
1!
1%
#249940000000
0!
0%
#249945000000
1!
1%
#249950000000
0!
0%
#249955000000
1!
1%
#249960000000
0!
0%
#249965000000
1!
1%
#249970000000
0!
0%
#249975000000
1!
1%
#249980000000
0!
0%
#249985000000
1!
1%
#249990000000
0!
0%
#249995000000
1!
1%
#250000000000
0!
0%
#250005000000
1!
1%
#250010000000
0!
0%
#250015000000
1!
1%
#250020000000
0!
0%
#250025000000
1!
1%
#250030000000
0!
0%
#250035000000
1!
1%
#250040000000
0!
0%
#250045000000
1!
1%
#250050000000
0!
0%
#250055000000
1!
1%
#250060000000
0!
0%
#250065000000
1!
1%
#250070000000
0!
0%
#250075000000
1!
1%
#250080000000
0!
0%
#250085000000
1!
1%
#250090000000
0!
0%
#250095000000
1!
1%
#250100000000
0!
0%
#250105000000
1!
1%
#250110000000
0!
0%
#250115000000
1!
1%
#250120000000
0!
0%
#250125000000
1!
1%
#250130000000
0!
0%
#250135000000
1!
1%
#250140000000
0!
0%
#250145000000
1!
1%
#250150000000
0!
0%
#250155000000
1!
1%
#250160000000
0!
0%
#250165000000
1!
1%
#250170000000
0!
0%
#250175000000
1!
1%
#250180000000
0!
0%
#250185000000
1!
1%
#250190000000
0!
0%
#250195000000
1!
1%
#250200000000
0!
0%
#250205000000
1!
1%
#250210000000
0!
0%
#250215000000
1!
1%
#250220000000
0!
0%
#250225000000
1!
1%
#250230000000
0!
0%
#250235000000
1!
1%
#250240000000
0!
0%
#250245000000
1!
1%
#250250000000
0!
0%
#250255000000
1!
1%
#250260000000
0!
0%
#250265000000
1!
1%
#250270000000
0!
0%
#250275000000
1!
1%
#250280000000
0!
0%
#250285000000
1!
1%
#250290000000
0!
0%
#250295000000
1!
1%
#250300000000
0!
0%
#250305000000
1!
1%
#250310000000
0!
0%
#250315000000
1!
1%
#250320000000
0!
0%
#250325000000
1!
1%
#250330000000
0!
0%
#250335000000
1!
1%
#250340000000
0!
0%
#250345000000
1!
1%
#250350000000
0!
0%
#250355000000
1!
1%
#250360000000
0!
0%
#250365000000
1!
1%
#250370000000
0!
0%
#250375000000
1!
1%
#250380000000
0!
0%
#250385000000
1!
1%
#250390000000
0!
0%
#250395000000
1!
1%
#250400000000
0!
0%
#250405000000
1!
1%
#250410000000
0!
0%
#250415000000
1!
1%
#250420000000
0!
0%
#250425000000
1!
1%
#250430000000
0!
0%
#250435000000
1!
1%
#250440000000
0!
0%
#250445000000
1!
1%
#250450000000
0!
0%
#250455000000
1!
1%
#250460000000
0!
0%
#250465000000
1!
1%
#250470000000
0!
0%
#250475000000
1!
1%
#250480000000
0!
0%
#250485000000
1!
1%
#250490000000
0!
0%
#250495000000
1!
1%
#250500000000
0!
0%
#250505000000
1!
1%
#250510000000
0!
0%
#250515000000
1!
1%
#250520000000
0!
0%
#250525000000
1!
1%
#250530000000
0!
0%
#250535000000
1!
1%
#250540000000
0!
0%
#250545000000
1!
1%
#250550000000
0!
0%
#250555000000
1!
1%
#250560000000
0!
0%
#250565000000
1!
1%
#250570000000
0!
0%
#250575000000
1!
1%
#250580000000
0!
0%
#250585000000
1!
1%
#250590000000
0!
0%
#250595000000
1!
1%
#250600000000
0!
0%
#250605000000
1!
1%
#250610000000
0!
0%
#250615000000
1!
1%
#250620000000
0!
0%
#250625000000
1!
1%
#250630000000
0!
0%
#250635000000
1!
1%
#250640000000
0!
0%
#250645000000
1!
1%
#250650000000
0!
0%
#250655000000
1!
1%
#250660000000
0!
0%
#250665000000
1!
1%
#250670000000
0!
0%
#250675000000
1!
1%
#250680000000
0!
0%
#250685000000
1!
1%
#250690000000
0!
0%
#250695000000
1!
1%
#250700000000
0!
0%
#250705000000
1!
1%
#250710000000
0!
0%
#250715000000
1!
1%
#250720000000
0!
0%
#250725000000
1!
1%
#250730000000
0!
0%
#250735000000
1!
1%
#250740000000
0!
0%
#250745000000
1!
1%
#250750000000
0!
0%
#250755000000
1!
1%
#250760000000
0!
0%
#250765000000
1!
1%
#250770000000
0!
0%
#250775000000
1!
1%
#250780000000
0!
0%
#250785000000
1!
1%
#250790000000
0!
0%
#250795000000
1!
1%
#250800000000
0!
0%
#250805000000
1!
1%
#250810000000
0!
0%
#250815000000
1!
1%
#250820000000
0!
0%
#250825000000
1!
1%
#250830000000
0!
0%
#250835000000
1!
1%
#250840000000
0!
0%
#250845000000
1!
1%
#250850000000
0!
0%
#250855000000
1!
1%
#250860000000
0!
0%
#250865000000
1!
1%
#250870000000
0!
0%
#250875000000
1!
1%
#250880000000
0!
0%
#250885000000
1!
1%
#250890000000
0!
0%
#250895000000
1!
1%
#250900000000
0!
0%
#250905000000
1!
1%
#250910000000
0!
0%
#250915000000
1!
1%
#250920000000
0!
0%
#250925000000
1!
1%
#250930000000
0!
0%
#250935000000
1!
1%
#250940000000
0!
0%
#250945000000
1!
1%
#250950000000
0!
0%
#250955000000
1!
1%
#250960000000
0!
0%
#250965000000
1!
1%
#250970000000
0!
0%
#250975000000
1!
1%
#250980000000
0!
0%
#250985000000
1!
1%
#250990000000
0!
0%
#250995000000
1!
1%
#251000000000
0!
0%
#251005000000
1!
1%
#251010000000
0!
0%
#251015000000
1!
1%
#251020000000
0!
0%
#251025000000
1!
1%
#251030000000
0!
0%
#251035000000
1!
1%
#251040000000
0!
0%
#251045000000
1!
1%
#251050000000
0!
0%
#251055000000
1!
1%
#251060000000
0!
0%
#251065000000
1!
1%
#251070000000
0!
0%
#251075000000
1!
1%
#251080000000
0!
0%
#251085000000
1!
1%
#251090000000
0!
0%
#251095000000
1!
1%
#251100000000
0!
0%
#251105000000
1!
1%
#251110000000
0!
0%
#251115000000
1!
1%
#251120000000
0!
0%
#251125000000
1!
1%
#251130000000
0!
0%
#251135000000
1!
1%
#251140000000
0!
0%
#251145000000
1!
1%
#251150000000
0!
0%
#251155000000
1!
1%
#251160000000
0!
0%
#251165000000
1!
1%
#251170000000
0!
0%
#251175000000
1!
1%
#251180000000
0!
0%
#251185000000
1!
1%
#251190000000
0!
0%
#251195000000
1!
1%
#251200000000
0!
0%
#251205000000
1!
1%
#251210000000
0!
0%
#251215000000
1!
1%
#251220000000
0!
0%
#251225000000
1!
1%
#251230000000
0!
0%
#251235000000
1!
1%
#251240000000
0!
0%
#251245000000
1!
1%
#251250000000
0!
0%
#251255000000
1!
1%
#251260000000
0!
0%
#251265000000
1!
1%
#251270000000
0!
0%
#251275000000
1!
1%
#251280000000
0!
0%
#251285000000
1!
1%
#251290000000
0!
0%
#251295000000
1!
1%
#251300000000
0!
0%
#251305000000
1!
1%
#251310000000
0!
0%
#251315000000
1!
1%
#251320000000
0!
0%
#251325000000
1!
1%
#251330000000
0!
0%
#251335000000
1!
1%
#251340000000
0!
0%
#251345000000
1!
1%
#251350000000
0!
0%
#251355000000
1!
1%
#251360000000
0!
0%
#251365000000
1!
1%
#251370000000
0!
0%
#251375000000
1!
1%
#251380000000
0!
0%
#251385000000
1!
1%
#251390000000
0!
0%
#251395000000
1!
1%
#251400000000
0!
0%
#251405000000
1!
1%
#251410000000
0!
0%
#251415000000
1!
1%
#251420000000
0!
0%
#251425000000
1!
1%
#251430000000
0!
0%
#251435000000
1!
1%
#251440000000
0!
0%
#251445000000
1!
1%
#251450000000
0!
0%
#251455000000
1!
1%
#251460000000
0!
0%
#251465000000
1!
1%
#251470000000
0!
0%
#251475000000
1!
1%
#251480000000
0!
0%
#251485000000
1!
1%
#251490000000
0!
0%
#251495000000
1!
1%
#251500000000
0!
0%
#251505000000
1!
1%
#251510000000
0!
0%
#251515000000
1!
1%
#251520000000
0!
0%
#251525000000
1!
1%
#251530000000
0!
0%
#251535000000
1!
1%
#251540000000
0!
0%
#251545000000
1!
1%
#251550000000
0!
0%
#251555000000
1!
1%
#251560000000
0!
0%
#251565000000
1!
1%
#251570000000
0!
0%
#251575000000
1!
1%
#251580000000
0!
0%
#251585000000
1!
1%
#251590000000
0!
0%
#251595000000
1!
1%
#251600000000
0!
0%
#251605000000
1!
1%
#251610000000
0!
0%
#251615000000
1!
1%
#251620000000
0!
0%
#251625000000
1!
1%
#251630000000
0!
0%
#251635000000
1!
1%
#251640000000
0!
0%
#251645000000
1!
1%
#251650000000
0!
0%
#251655000000
1!
1%
#251660000000
0!
0%
#251665000000
1!
1%
#251670000000
0!
0%
#251675000000
1!
1%
#251680000000
0!
0%
#251685000000
1!
1%
#251690000000
0!
0%
#251695000000
1!
1%
#251700000000
0!
0%
#251705000000
1!
1%
#251710000000
0!
0%
#251715000000
1!
1%
#251720000000
0!
0%
#251725000000
1!
1%
#251730000000
0!
0%
#251735000000
1!
1%
#251740000000
0!
0%
#251745000000
1!
1%
#251750000000
0!
0%
#251755000000
1!
1%
#251760000000
0!
0%
#251765000000
1!
1%
#251770000000
0!
0%
#251775000000
1!
1%
#251780000000
0!
0%
#251785000000
1!
1%
#251790000000
0!
0%
#251795000000
1!
1%
#251800000000
0!
0%
#251805000000
1!
1%
#251810000000
0!
0%
#251815000000
1!
1%
#251820000000
0!
0%
#251825000000
1!
1%
#251830000000
0!
0%
#251835000000
1!
1%
#251840000000
0!
0%
#251845000000
1!
1%
#251850000000
0!
0%
#251855000000
1!
1%
#251860000000
0!
0%
#251865000000
1!
1%
#251870000000
0!
0%
#251875000000
1!
1%
#251880000000
0!
0%
#251885000000
1!
1%
#251890000000
0!
0%
#251895000000
1!
1%
#251900000000
0!
0%
#251905000000
1!
1%
#251910000000
0!
0%
#251915000000
1!
1%
#251920000000
0!
0%
#251925000000
1!
1%
#251930000000
0!
0%
#251935000000
1!
1%
#251940000000
0!
0%
#251945000000
1!
1%
#251950000000
0!
0%
#251955000000
1!
1%
#251960000000
0!
0%
#251965000000
1!
1%
#251970000000
0!
0%
#251975000000
1!
1%
#251980000000
0!
0%
#251985000000
1!
1%
#251990000000
0!
0%
#251995000000
1!
1%
#252000000000
0!
0%
#252005000000
1!
1%
#252010000000
0!
0%
#252015000000
1!
1%
#252020000000
0!
0%
#252025000000
1!
1%
#252030000000
0!
0%
#252035000000
1!
1%
#252040000000
0!
0%
#252045000000
1!
1%
#252050000000
0!
0%
#252055000000
1!
1%
#252060000000
0!
0%
#252065000000
1!
1%
#252070000000
0!
0%
#252075000000
1!
1%
#252080000000
0!
0%
#252085000000
1!
1%
#252090000000
0!
0%
#252095000000
1!
1%
#252100000000
0!
0%
#252105000000
1!
1%
#252110000000
0!
0%
#252115000000
1!
1%
#252120000000
0!
0%
#252125000000
1!
1%
#252130000000
0!
0%
#252135000000
1!
1%
#252140000000
0!
0%
#252145000000
1!
1%
#252150000000
0!
0%
#252155000000
1!
1%
#252160000000
0!
0%
#252165000000
1!
1%
#252170000000
0!
0%
#252175000000
1!
1%
#252180000000
0!
0%
#252185000000
1!
1%
#252190000000
0!
0%
#252195000000
1!
1%
#252200000000
0!
0%
#252205000000
1!
1%
#252210000000
0!
0%
#252215000000
1!
1%
#252220000000
0!
0%
#252225000000
1!
1%
#252230000000
0!
0%
#252235000000
1!
1%
#252240000000
0!
0%
#252245000000
1!
1%
#252250000000
0!
0%
#252255000000
1!
1%
#252260000000
0!
0%
#252265000000
1!
1%
#252270000000
0!
0%
#252275000000
1!
1%
#252280000000
0!
0%
#252285000000
1!
1%
#252290000000
0!
0%
#252295000000
1!
1%
#252300000000
0!
0%
#252305000000
1!
1%
#252310000000
0!
0%
#252315000000
1!
1%
#252320000000
0!
0%
#252325000000
1!
1%
#252330000000
0!
0%
#252335000000
1!
1%
#252340000000
0!
0%
#252345000000
1!
1%
#252350000000
0!
0%
#252355000000
1!
1%
#252360000000
0!
0%
#252365000000
1!
1%
#252370000000
0!
0%
#252375000000
1!
1%
#252380000000
0!
0%
#252385000000
1!
1%
#252390000000
0!
0%
#252395000000
1!
1%
#252400000000
0!
0%
#252405000000
1!
1%
#252410000000
0!
0%
#252415000000
1!
1%
#252420000000
0!
0%
#252425000000
1!
1%
#252430000000
0!
0%
#252435000000
1!
1%
#252440000000
0!
0%
#252445000000
1!
1%
#252450000000
0!
0%
#252455000000
1!
1%
#252460000000
0!
0%
#252465000000
1!
1%
#252470000000
0!
0%
#252475000000
1!
1%
#252480000000
0!
0%
#252485000000
1!
1%
#252490000000
0!
0%
#252495000000
1!
1%
#252500000000
0!
0%
#252505000000
1!
1%
#252510000000
0!
0%
#252515000000
1!
1%
#252520000000
0!
0%
#252525000000
1!
1%
#252530000000
0!
0%
#252535000000
1!
1%
#252540000000
0!
0%
#252545000000
1!
1%
#252550000000
0!
0%
#252555000000
1!
1%
#252560000000
0!
0%
#252565000000
1!
1%
#252570000000
0!
0%
#252575000000
1!
1%
#252580000000
0!
0%
#252585000000
1!
1%
#252590000000
0!
0%
#252595000000
1!
1%
#252600000000
0!
0%
#252605000000
1!
1%
#252610000000
0!
0%
#252615000000
1!
1%
#252620000000
0!
0%
#252625000000
1!
1%
#252630000000
0!
0%
#252635000000
1!
1%
#252640000000
0!
0%
#252645000000
1!
1%
#252650000000
0!
0%
#252655000000
1!
1%
#252660000000
0!
0%
#252665000000
1!
1%
#252670000000
0!
0%
#252675000000
1!
1%
#252680000000
0!
0%
#252685000000
1!
1%
#252690000000
0!
0%
#252695000000
1!
1%
#252700000000
0!
0%
#252705000000
1!
1%
#252710000000
0!
0%
#252715000000
1!
1%
#252720000000
0!
0%
#252725000000
1!
1%
#252730000000
0!
0%
#252735000000
1!
1%
#252740000000
0!
0%
#252745000000
1!
1%
#252750000000
0!
0%
#252755000000
1!
1%
#252760000000
0!
0%
#252765000000
1!
1%
#252770000000
0!
0%
#252775000000
1!
1%
#252780000000
0!
0%
#252785000000
1!
1%
#252790000000
0!
0%
#252795000000
1!
1%
#252800000000
0!
0%
#252805000000
1!
1%
#252810000000
0!
0%
#252815000000
1!
1%
#252820000000
0!
0%
#252825000000
1!
1%
#252830000000
0!
0%
#252835000000
1!
1%
#252840000000
0!
0%
#252845000000
1!
1%
#252850000000
0!
0%
#252855000000
1!
1%
#252860000000
0!
0%
#252865000000
1!
1%
#252870000000
0!
0%
#252875000000
1!
1%
#252880000000
0!
0%
#252885000000
1!
1%
#252890000000
0!
0%
#252895000000
1!
1%
#252900000000
0!
0%
#252905000000
1!
1%
#252910000000
0!
0%
#252915000000
1!
1%
#252920000000
0!
0%
#252925000000
1!
1%
#252930000000
0!
0%
#252935000000
1!
1%
#252940000000
0!
0%
#252945000000
1!
1%
#252950000000
0!
0%
#252955000000
1!
1%
#252960000000
0!
0%
#252965000000
1!
1%
#252970000000
0!
0%
#252975000000
1!
1%
#252980000000
0!
0%
#252985000000
1!
1%
#252990000000
0!
0%
#252995000000
1!
1%
#253000000000
0!
0%
#253005000000
1!
1%
#253010000000
0!
0%
#253015000000
1!
1%
#253020000000
0!
0%
#253025000000
1!
1%
#253030000000
0!
0%
#253035000000
1!
1%
#253040000000
0!
0%
#253045000000
1!
1%
#253050000000
0!
0%
#253055000000
1!
1%
#253060000000
0!
0%
#253065000000
1!
1%
#253070000000
0!
0%
#253075000000
1!
1%
#253080000000
0!
0%
#253085000000
1!
1%
#253090000000
0!
0%
#253095000000
1!
1%
#253100000000
0!
0%
#253105000000
1!
1%
#253110000000
0!
0%
#253115000000
1!
1%
#253120000000
0!
0%
#253125000000
1!
1%
#253130000000
0!
0%
#253135000000
1!
1%
#253140000000
0!
0%
#253145000000
1!
1%
#253150000000
0!
0%
#253155000000
1!
1%
#253160000000
0!
0%
#253165000000
1!
1%
#253170000000
0!
0%
#253175000000
1!
1%
#253180000000
0!
0%
#253185000000
1!
1%
#253190000000
0!
0%
#253195000000
1!
1%
#253200000000
0!
0%
#253205000000
1!
1%
#253210000000
0!
0%
#253215000000
1!
1%
#253220000000
0!
0%
#253225000000
1!
1%
#253230000000
0!
0%
#253235000000
1!
1%
#253240000000
0!
0%
#253245000000
1!
1%
#253250000000
0!
0%
#253255000000
1!
1%
#253260000000
0!
0%
#253265000000
1!
1%
#253270000000
0!
0%
#253275000000
1!
1%
#253280000000
0!
0%
#253285000000
1!
1%
#253290000000
0!
0%
#253295000000
1!
1%
#253300000000
0!
0%
#253305000000
1!
1%
#253310000000
0!
0%
#253315000000
1!
1%
#253320000000
0!
0%
#253325000000
1!
1%
#253330000000
0!
0%
#253335000000
1!
1%
#253340000000
0!
0%
#253345000000
1!
1%
#253350000000
0!
0%
#253355000000
1!
1%
#253360000000
0!
0%
#253365000000
1!
1%
#253370000000
0!
0%
#253375000000
1!
1%
#253380000000
0!
0%
#253385000000
1!
1%
#253390000000
0!
0%
#253395000000
1!
1%
#253400000000
0!
0%
#253405000000
1!
1%
#253410000000
0!
0%
#253415000000
1!
1%
#253420000000
0!
0%
#253425000000
1!
1%
#253430000000
0!
0%
#253435000000
1!
1%
#253440000000
0!
0%
#253445000000
1!
1%
#253450000000
0!
0%
#253455000000
1!
1%
#253460000000
0!
0%
#253465000000
1!
1%
#253470000000
0!
0%
#253475000000
1!
1%
#253480000000
0!
0%
#253485000000
1!
1%
#253490000000
0!
0%
#253495000000
1!
1%
#253500000000
0!
0%
#253505000000
1!
1%
#253510000000
0!
0%
#253515000000
1!
1%
#253520000000
0!
0%
#253525000000
1!
1%
#253530000000
0!
0%
#253535000000
1!
1%
#253540000000
0!
0%
#253545000000
1!
1%
#253550000000
0!
0%
#253555000000
1!
1%
#253560000000
0!
0%
#253565000000
1!
1%
#253570000000
0!
0%
#253575000000
1!
1%
#253580000000
0!
0%
#253585000000
1!
1%
#253590000000
0!
0%
#253595000000
1!
1%
#253600000000
0!
0%
#253605000000
1!
1%
#253610000000
0!
0%
#253615000000
1!
1%
#253620000000
0!
0%
#253625000000
1!
1%
#253630000000
0!
0%
#253635000000
1!
1%
#253640000000
0!
0%
#253645000000
1!
1%
#253650000000
0!
0%
#253655000000
1!
1%
#253660000000
0!
0%
#253665000000
1!
1%
#253670000000
0!
0%
#253675000000
1!
1%
#253680000000
0!
0%
#253685000000
1!
1%
#253690000000
0!
0%
#253695000000
1!
1%
#253700000000
0!
0%
#253705000000
1!
1%
#253710000000
0!
0%
#253715000000
1!
1%
#253720000000
0!
0%
#253725000000
1!
1%
#253730000000
0!
0%
#253735000000
1!
1%
#253740000000
0!
0%
#253745000000
1!
1%
#253750000000
0!
0%
#253755000000
1!
1%
#253760000000
0!
0%
#253765000000
1!
1%
#253770000000
0!
0%
#253775000000
1!
1%
#253780000000
0!
0%
#253785000000
1!
1%
#253790000000
0!
0%
#253795000000
1!
1%
#253800000000
0!
0%
#253805000000
1!
1%
#253810000000
0!
0%
#253815000000
1!
1%
#253820000000
0!
0%
#253825000000
1!
1%
#253830000000
0!
0%
#253835000000
1!
1%
#253840000000
0!
0%
#253845000000
1!
1%
#253850000000
0!
0%
#253855000000
1!
1%
#253860000000
0!
0%
#253865000000
1!
1%
#253870000000
0!
0%
#253875000000
1!
1%
#253880000000
0!
0%
#253885000000
1!
1%
#253890000000
0!
0%
#253895000000
1!
1%
#253900000000
0!
0%
#253905000000
1!
1%
#253910000000
0!
0%
#253915000000
1!
1%
#253920000000
0!
0%
#253925000000
1!
1%
#253930000000
0!
0%
#253935000000
1!
1%
#253940000000
0!
0%
#253945000000
1!
1%
#253950000000
0!
0%
#253955000000
1!
1%
#253960000000
0!
0%
#253965000000
1!
1%
#253970000000
0!
0%
#253975000000
1!
1%
#253980000000
0!
0%
#253985000000
1!
1%
#253990000000
0!
0%
#253995000000
1!
1%
#254000000000
0!
0%
#254005000000
1!
1%
#254010000000
0!
0%
#254015000000
1!
1%
#254020000000
0!
0%
#254025000000
1!
1%
#254030000000
0!
0%
#254035000000
1!
1%
#254040000000
0!
0%
#254045000000
1!
1%
#254050000000
0!
0%
#254055000000
1!
1%
#254060000000
0!
0%
#254065000000
1!
1%
#254070000000
0!
0%
#254075000000
1!
1%
#254080000000
0!
0%
#254085000000
1!
1%
#254090000000
0!
0%
#254095000000
1!
1%
#254100000000
0!
0%
#254105000000
1!
1%
#254110000000
0!
0%
#254115000000
1!
1%
#254120000000
0!
0%
#254125000000
1!
1%
#254130000000
0!
0%
#254135000000
1!
1%
#254140000000
0!
0%
#254145000000
1!
1%
#254150000000
0!
0%
#254155000000
1!
1%
#254160000000
0!
0%
#254165000000
1!
1%
#254170000000
0!
0%
#254175000000
1!
1%
#254180000000
0!
0%
#254185000000
1!
1%
#254190000000
0!
0%
#254195000000
1!
1%
#254200000000
0!
0%
#254205000000
1!
1%
#254210000000
0!
0%
#254215000000
1!
1%
#254220000000
0!
0%
#254225000000
1!
1%
#254230000000
0!
0%
#254235000000
1!
1%
#254240000000
0!
0%
#254245000000
1!
1%
#254250000000
0!
0%
#254255000000
1!
1%
#254260000000
0!
0%
#254265000000
1!
1%
#254270000000
0!
0%
#254275000000
1!
1%
#254280000000
0!
0%
#254285000000
1!
1%
#254290000000
0!
0%
#254295000000
1!
1%
#254300000000
0!
0%
#254305000000
1!
1%
#254310000000
0!
0%
#254315000000
1!
1%
#254320000000
0!
0%
#254325000000
1!
1%
#254330000000
0!
0%
#254335000000
1!
1%
#254340000000
0!
0%
#254345000000
1!
1%
#254350000000
0!
0%
#254355000000
1!
1%
#254360000000
0!
0%
#254365000000
1!
1%
#254370000000
0!
0%
#254375000000
1!
1%
#254380000000
0!
0%
#254385000000
1!
1%
#254390000000
0!
0%
#254395000000
1!
1%
#254400000000
0!
0%
#254405000000
1!
1%
#254410000000
0!
0%
#254415000000
1!
1%
#254420000000
0!
0%
#254425000000
1!
1%
#254430000000
0!
0%
#254435000000
1!
1%
#254440000000
0!
0%
#254445000000
1!
1%
#254450000000
0!
0%
#254455000000
1!
1%
#254460000000
0!
0%
#254465000000
1!
1%
#254470000000
0!
0%
#254475000000
1!
1%
#254480000000
0!
0%
#254485000000
1!
1%
#254490000000
0!
0%
#254495000000
1!
1%
#254500000000
0!
0%
#254505000000
1!
1%
#254510000000
0!
0%
#254515000000
1!
1%
#254520000000
0!
0%
#254525000000
1!
1%
#254530000000
0!
0%
#254535000000
1!
1%
#254540000000
0!
0%
#254545000000
1!
1%
#254550000000
0!
0%
#254555000000
1!
1%
#254560000000
0!
0%
#254565000000
1!
1%
#254570000000
0!
0%
#254575000000
1!
1%
#254580000000
0!
0%
#254585000000
1!
1%
#254590000000
0!
0%
#254595000000
1!
1%
#254600000000
0!
0%
#254605000000
1!
1%
#254610000000
0!
0%
#254615000000
1!
1%
#254620000000
0!
0%
#254625000000
1!
1%
#254630000000
0!
0%
#254635000000
1!
1%
#254640000000
0!
0%
#254645000000
1!
1%
#254650000000
0!
0%
#254655000000
1!
1%
#254660000000
0!
0%
#254665000000
1!
1%
#254670000000
0!
0%
#254675000000
1!
1%
#254680000000
0!
0%
#254685000000
1!
1%
#254690000000
0!
0%
#254695000000
1!
1%
#254700000000
0!
0%
#254705000000
1!
1%
#254710000000
0!
0%
#254715000000
1!
1%
#254720000000
0!
0%
#254725000000
1!
1%
#254730000000
0!
0%
#254735000000
1!
1%
#254740000000
0!
0%
#254745000000
1!
1%
#254750000000
0!
0%
#254755000000
1!
1%
#254760000000
0!
0%
#254765000000
1!
1%
#254770000000
0!
0%
#254775000000
1!
1%
#254780000000
0!
0%
#254785000000
1!
1%
#254790000000
0!
0%
#254795000000
1!
1%
#254800000000
0!
0%
#254805000000
1!
1%
#254810000000
0!
0%
#254815000000
1!
1%
#254820000000
0!
0%
#254825000000
1!
1%
#254830000000
0!
0%
#254835000000
1!
1%
#254840000000
0!
0%
#254845000000
1!
1%
#254850000000
0!
0%
#254855000000
1!
1%
#254860000000
0!
0%
#254865000000
1!
1%
#254870000000
0!
0%
#254875000000
1!
1%
#254880000000
0!
0%
#254885000000
1!
1%
#254890000000
0!
0%
#254895000000
1!
1%
#254900000000
0!
0%
#254905000000
1!
1%
#254910000000
0!
0%
#254915000000
1!
1%
#254920000000
0!
0%
#254925000000
1!
1%
#254930000000
0!
0%
#254935000000
1!
1%
#254940000000
0!
0%
#254945000000
1!
1%
#254950000000
0!
0%
#254955000000
1!
1%
#254960000000
0!
0%
#254965000000
1!
1%
#254970000000
0!
0%
#254975000000
1!
1%
#254980000000
0!
0%
#254985000000
1!
1%
#254990000000
0!
0%
#254995000000
1!
1%
#255000000000
0!
0%
#255005000000
1!
1%
#255010000000
0!
0%
#255015000000
1!
1%
#255020000000
0!
0%
#255025000000
1!
1%
#255030000000
0!
0%
#255035000000
1!
1%
#255040000000
0!
0%
#255045000000
1!
1%
#255050000000
0!
0%
#255055000000
1!
1%
#255060000000
0!
0%
#255065000000
1!
1%
#255070000000
0!
0%
#255075000000
1!
1%
#255080000000
0!
0%
#255085000000
1!
1%
#255090000000
0!
0%
#255095000000
1!
1%
#255100000000
0!
0%
#255105000000
1!
1%
#255110000000
0!
0%
#255115000000
1!
1%
#255120000000
0!
0%
#255125000000
1!
1%
#255130000000
0!
0%
#255135000000
1!
1%
#255140000000
0!
0%
#255145000000
1!
1%
#255150000000
0!
0%
#255155000000
1!
1%
#255160000000
0!
0%
#255165000000
1!
1%
#255170000000
0!
0%
#255175000000
1!
1%
#255180000000
0!
0%
#255185000000
1!
1%
#255190000000
0!
0%
#255195000000
1!
1%
#255200000000
0!
0%
#255205000000
1!
1%
#255210000000
0!
0%
#255215000000
1!
1%
#255220000000
0!
0%
#255225000000
1!
1%
#255230000000
0!
0%
#255235000000
1!
1%
#255240000000
0!
0%
#255245000000
1!
1%
#255250000000
0!
0%
#255255000000
1!
1%
#255260000000
0!
0%
#255265000000
1!
1%
#255270000000
0!
0%
#255275000000
1!
1%
#255280000000
0!
0%
#255285000000
1!
1%
#255290000000
0!
0%
#255295000000
1!
1%
#255300000000
0!
0%
#255305000000
1!
1%
#255310000000
0!
0%
#255315000000
1!
1%
#255320000000
0!
0%
#255325000000
1!
1%
#255330000000
0!
0%
#255335000000
1!
1%
#255340000000
0!
0%
#255345000000
1!
1%
#255350000000
0!
0%
#255355000000
1!
1%
#255360000000
0!
0%
#255365000000
1!
1%
#255370000000
0!
0%
#255375000000
1!
1%
#255380000000
0!
0%
#255385000000
1!
1%
#255390000000
0!
0%
#255395000000
1!
1%
#255400000000
0!
0%
#255405000000
1!
1%
#255410000000
0!
0%
#255415000000
1!
1%
#255420000000
0!
0%
#255425000000
1!
1%
#255430000000
0!
0%
#255435000000
1!
1%
#255440000000
0!
0%
#255445000000
1!
1%
#255450000000
0!
0%
#255455000000
1!
1%
#255460000000
0!
0%
#255465000000
1!
1%
#255470000000
0!
0%
#255475000000
1!
1%
#255480000000
0!
0%
#255485000000
1!
1%
#255490000000
0!
0%
#255495000000
1!
1%
#255500000000
0!
0%
#255505000000
1!
1%
#255510000000
0!
0%
#255515000000
1!
1%
#255520000000
0!
0%
#255525000000
1!
1%
#255530000000
0!
0%
#255535000000
1!
1%
#255540000000
0!
0%
#255545000000
1!
1%
#255550000000
0!
0%
#255555000000
1!
1%
#255560000000
0!
0%
#255565000000
1!
1%
#255570000000
0!
0%
#255575000000
1!
1%
#255580000000
0!
0%
#255585000000
1!
1%
#255590000000
0!
0%
#255595000000
1!
1%
#255600000000
0!
0%
#255605000000
1!
1%
#255610000000
0!
0%
#255615000000
1!
1%
#255620000000
0!
0%
#255625000000
1!
1%
#255630000000
0!
0%
#255635000000
1!
1%
#255640000000
0!
0%
#255645000000
1!
1%
#255650000000
0!
0%
#255655000000
1!
1%
#255660000000
0!
0%
#255665000000
1!
1%
#255670000000
0!
0%
#255675000000
1!
1%
#255680000000
0!
0%
#255685000000
1!
1%
#255690000000
0!
0%
#255695000000
1!
1%
#255700000000
0!
0%
#255705000000
1!
1%
#255710000000
0!
0%
#255715000000
1!
1%
#255720000000
0!
0%
#255725000000
1!
1%
#255730000000
0!
0%
#255735000000
1!
1%
#255740000000
0!
0%
#255745000000
1!
1%
#255750000000
0!
0%
#255755000000
1!
1%
#255760000000
0!
0%
#255765000000
1!
1%
#255770000000
0!
0%
#255775000000
1!
1%
#255780000000
0!
0%
#255785000000
1!
1%
#255790000000
0!
0%
#255795000000
1!
1%
#255800000000
0!
0%
#255805000000
1!
1%
#255810000000
0!
0%
#255815000000
1!
1%
#255820000000
0!
0%
#255825000000
1!
1%
#255830000000
0!
0%
#255835000000
1!
1%
#255840000000
0!
0%
#255845000000
1!
1%
#255850000000
0!
0%
#255855000000
1!
1%
#255860000000
0!
0%
#255865000000
1!
1%
#255870000000
0!
0%
#255875000000
1!
1%
#255880000000
0!
0%
#255885000000
1!
1%
#255890000000
0!
0%
#255895000000
1!
1%
#255900000000
0!
0%
#255905000000
1!
1%
#255910000000
0!
0%
#255915000000
1!
1%
#255920000000
0!
0%
#255925000000
1!
1%
#255930000000
0!
0%
#255935000000
1!
1%
#255940000000
0!
0%
#255945000000
1!
1%
#255950000000
0!
0%
#255955000000
1!
1%
#255960000000
0!
0%
#255965000000
1!
1%
#255970000000
0!
0%
#255975000000
1!
1%
#255980000000
0!
0%
#255985000000
1!
1%
#255990000000
0!
0%
#255995000000
1!
1%
#256000000000
0!
0%
#256005000000
1!
1%
#256010000000
0!
0%
#256015000000
1!
1%
#256020000000
0!
0%
#256025000000
1!
1%
#256030000000
0!
0%
#256035000000
1!
1%
#256040000000
0!
0%
#256045000000
1!
1%
#256050000000
0!
0%
#256055000000
1!
1%
#256060000000
0!
0%
#256065000000
1!
1%
#256070000000
0!
0%
#256075000000
1!
1%
#256080000000
0!
0%
#256085000000
1!
1%
#256090000000
0!
0%
#256095000000
1!
1%
#256100000000
0!
0%
#256105000000
1!
1%
#256110000000
0!
0%
#256115000000
1!
1%
#256120000000
0!
0%
#256125000000
1!
1%
#256130000000
0!
0%
#256135000000
1!
1%
#256140000000
0!
0%
#256145000000
1!
1%
#256150000000
0!
0%
#256155000000
1!
1%
#256160000000
0!
0%
#256165000000
1!
1%
#256170000000
0!
0%
#256175000000
1!
1%
#256180000000
0!
0%
#256185000000
1!
1%
#256190000000
0!
0%
#256195000000
1!
1%
#256200000000
0!
0%
#256205000000
1!
1%
#256210000000
0!
0%
#256215000000
1!
1%
#256220000000
0!
0%
#256225000000
1!
1%
#256230000000
0!
0%
#256235000000
1!
1%
#256240000000
0!
0%
#256245000000
1!
1%
#256250000000
0!
0%
#256255000000
1!
1%
#256260000000
0!
0%
#256265000000
1!
1%
#256270000000
0!
0%
#256275000000
1!
1%
#256280000000
0!
0%
#256285000000
1!
1%
#256290000000
0!
0%
#256295000000
1!
1%
#256300000000
0!
0%
#256305000000
1!
1%
#256310000000
0!
0%
#256315000000
1!
1%
#256320000000
0!
0%
#256325000000
1!
1%
#256330000000
0!
0%
#256335000000
1!
1%
#256340000000
0!
0%
#256345000000
1!
1%
#256350000000
0!
0%
#256355000000
1!
1%
#256360000000
0!
0%
#256365000000
1!
1%
#256370000000
0!
0%
#256375000000
1!
1%
#256380000000
0!
0%
#256385000000
1!
1%
#256390000000
0!
0%
#256395000000
1!
1%
#256400000000
0!
0%
#256405000000
1!
1%
#256410000000
0!
0%
#256415000000
1!
1%
#256420000000
0!
0%
#256425000000
1!
1%
#256430000000
0!
0%
#256435000000
1!
1%
#256440000000
0!
0%
#256445000000
1!
1%
#256450000000
0!
0%
#256455000000
1!
1%
#256460000000
0!
0%
#256465000000
1!
1%
#256470000000
0!
0%
#256475000000
1!
1%
#256480000000
0!
0%
#256485000000
1!
1%
#256490000000
0!
0%
#256495000000
1!
1%
#256500000000
0!
0%
#256505000000
1!
1%
#256510000000
0!
0%
#256515000000
1!
1%
#256520000000
0!
0%
#256525000000
1!
1%
#256530000000
0!
0%
#256535000000
1!
1%
#256540000000
0!
0%
#256545000000
1!
1%
#256550000000
0!
0%
#256555000000
1!
1%
#256560000000
0!
0%
#256565000000
1!
1%
#256570000000
0!
0%
#256575000000
1!
1%
#256580000000
0!
0%
#256585000000
1!
1%
#256590000000
0!
0%
#256595000000
1!
1%
#256600000000
0!
0%
#256605000000
1!
1%
#256610000000
0!
0%
#256615000000
1!
1%
#256620000000
0!
0%
#256625000000
1!
1%
#256630000000
0!
0%
#256635000000
1!
1%
#256640000000
0!
0%
#256645000000
1!
1%
#256650000000
0!
0%
#256655000000
1!
1%
#256660000000
0!
0%
#256665000000
1!
1%
#256670000000
0!
0%
#256675000000
1!
1%
#256680000000
0!
0%
#256685000000
1!
1%
#256690000000
0!
0%
#256695000000
1!
1%
#256700000000
0!
0%
#256705000000
1!
1%
#256710000000
0!
0%
#256715000000
1!
1%
#256720000000
0!
0%
#256725000000
1!
1%
#256730000000
0!
0%
#256735000000
1!
1%
#256740000000
0!
0%
#256745000000
1!
1%
#256750000000
0!
0%
#256755000000
1!
1%
#256760000000
0!
0%
#256765000000
1!
1%
#256770000000
0!
0%
#256775000000
1!
1%
#256780000000
0!
0%
#256785000000
1!
1%
#256790000000
0!
0%
#256795000000
1!
1%
#256800000000
0!
0%
#256805000000
1!
1%
#256810000000
0!
0%
#256815000000
1!
1%
#256820000000
0!
0%
#256825000000
1!
1%
#256830000000
0!
0%
#256835000000
1!
1%
#256840000000
0!
0%
#256845000000
1!
1%
#256850000000
0!
0%
#256855000000
1!
1%
#256860000000
0!
0%
#256865000000
1!
1%
#256870000000
0!
0%
#256875000000
1!
1%
#256880000000
0!
0%
#256885000000
1!
1%
#256890000000
0!
0%
#256895000000
1!
1%
#256900000000
0!
0%
#256905000000
1!
1%
#256910000000
0!
0%
#256915000000
1!
1%
#256920000000
0!
0%
#256925000000
1!
1%
#256930000000
0!
0%
#256935000000
1!
1%
#256940000000
0!
0%
#256945000000
1!
1%
#256950000000
0!
0%
#256955000000
1!
1%
#256960000000
0!
0%
#256965000000
1!
1%
#256970000000
0!
0%
#256975000000
1!
1%
#256980000000
0!
0%
#256985000000
1!
1%
#256990000000
0!
0%
#256995000000
1!
1%
#257000000000
0!
0%
#257005000000
1!
1%
#257010000000
0!
0%
#257015000000
1!
1%
#257020000000
0!
0%
#257025000000
1!
1%
#257030000000
0!
0%
#257035000000
1!
1%
#257040000000
0!
0%
#257045000000
1!
1%
#257050000000
0!
0%
#257055000000
1!
1%
#257060000000
0!
0%
#257065000000
1!
1%
#257070000000
0!
0%
#257075000000
1!
1%
#257080000000
0!
0%
#257085000000
1!
1%
#257090000000
0!
0%
#257095000000
1!
1%
#257100000000
0!
0%
#257105000000
1!
1%
#257110000000
0!
0%
#257115000000
1!
1%
#257120000000
0!
0%
#257125000000
1!
1%
#257130000000
0!
0%
#257135000000
1!
1%
#257140000000
0!
0%
#257145000000
1!
1%
#257150000000
0!
0%
#257155000000
1!
1%
#257160000000
0!
0%
#257165000000
1!
1%
#257170000000
0!
0%
#257175000000
1!
1%
#257180000000
0!
0%
#257185000000
1!
1%
#257190000000
0!
0%
#257195000000
1!
1%
#257200000000
0!
0%
#257205000000
1!
1%
#257210000000
0!
0%
#257215000000
1!
1%
#257220000000
0!
0%
#257225000000
1!
1%
#257230000000
0!
0%
#257235000000
1!
1%
#257240000000
0!
0%
#257245000000
1!
1%
#257250000000
0!
0%
#257255000000
1!
1%
#257260000000
0!
0%
#257265000000
1!
1%
#257270000000
0!
0%
#257275000000
1!
1%
#257280000000
0!
0%
#257285000000
1!
1%
#257290000000
0!
0%
#257295000000
1!
1%
#257300000000
0!
0%
#257305000000
1!
1%
#257310000000
0!
0%
#257315000000
1!
1%
#257320000000
0!
0%
#257325000000
1!
1%
#257330000000
0!
0%
#257335000000
1!
1%
#257340000000
0!
0%
#257345000000
1!
1%
#257350000000
0!
0%
#257355000000
1!
1%
#257360000000
0!
0%
#257365000000
1!
1%
#257370000000
0!
0%
#257375000000
1!
1%
#257380000000
0!
0%
#257385000000
1!
1%
#257390000000
0!
0%
#257395000000
1!
1%
#257400000000
0!
0%
#257405000000
1!
1%
#257410000000
0!
0%
#257415000000
1!
1%
#257420000000
0!
0%
#257425000000
1!
1%
#257430000000
0!
0%
#257435000000
1!
1%
#257440000000
0!
0%
#257445000000
1!
1%
#257450000000
0!
0%
#257455000000
1!
1%
#257460000000
0!
0%
#257465000000
1!
1%
#257470000000
0!
0%
#257475000000
1!
1%
#257480000000
0!
0%
#257485000000
1!
1%
#257490000000
0!
0%
#257495000000
1!
1%
#257500000000
0!
0%
#257505000000
1!
1%
#257510000000
0!
0%
#257515000000
1!
1%
#257520000000
0!
0%
#257525000000
1!
1%
#257530000000
0!
0%
#257535000000
1!
1%
#257540000000
0!
0%
#257545000000
1!
1%
#257550000000
0!
0%
#257555000000
1!
1%
#257560000000
0!
0%
#257565000000
1!
1%
#257570000000
0!
0%
#257575000000
1!
1%
#257580000000
0!
0%
#257585000000
1!
1%
#257590000000
0!
0%
#257595000000
1!
1%
#257600000000
0!
0%
#257605000000
1!
1%
#257610000000
0!
0%
#257615000000
1!
1%
#257620000000
0!
0%
#257625000000
1!
1%
#257630000000
0!
0%
#257635000000
1!
1%
#257640000000
0!
0%
#257645000000
1!
1%
#257650000000
0!
0%
#257655000000
1!
1%
#257660000000
0!
0%
#257665000000
1!
1%
#257670000000
0!
0%
#257675000000
1!
1%
#257680000000
0!
0%
#257685000000
1!
1%
#257690000000
0!
0%
#257695000000
1!
1%
#257700000000
0!
0%
#257705000000
1!
1%
#257710000000
0!
0%
#257715000000
1!
1%
#257720000000
0!
0%
#257725000000
1!
1%
#257730000000
0!
0%
#257735000000
1!
1%
#257740000000
0!
0%
#257745000000
1!
1%
#257750000000
0!
0%
#257755000000
1!
1%
#257760000000
0!
0%
#257765000000
1!
1%
#257770000000
0!
0%
#257775000000
1!
1%
#257780000000
0!
0%
#257785000000
1!
1%
#257790000000
0!
0%
#257795000000
1!
1%
#257800000000
0!
0%
#257805000000
1!
1%
#257810000000
0!
0%
#257815000000
1!
1%
#257820000000
0!
0%
#257825000000
1!
1%
#257830000000
0!
0%
#257835000000
1!
1%
#257840000000
0!
0%
#257845000000
1!
1%
#257850000000
0!
0%
#257855000000
1!
1%
#257860000000
0!
0%
#257865000000
1!
1%
#257870000000
0!
0%
#257875000000
1!
1%
#257880000000
0!
0%
#257885000000
1!
1%
#257890000000
0!
0%
#257895000000
1!
1%
#257900000000
0!
0%
#257905000000
1!
1%
#257910000000
0!
0%
#257915000000
1!
1%
#257920000000
0!
0%
#257925000000
1!
1%
#257930000000
0!
0%
#257935000000
1!
1%
#257940000000
0!
0%
#257945000000
1!
1%
#257950000000
0!
0%
#257955000000
1!
1%
#257960000000
0!
0%
#257965000000
1!
1%
#257970000000
0!
0%
#257975000000
1!
1%
#257980000000
0!
0%
#257985000000
1!
1%
#257990000000
0!
0%
#257995000000
1!
1%
#258000000000
0!
0%
#258005000000
1!
1%
#258010000000
0!
0%
#258015000000
1!
1%
#258020000000
0!
0%
#258025000000
1!
1%
#258030000000
0!
0%
#258035000000
1!
1%
#258040000000
0!
0%
#258045000000
1!
1%
#258050000000
0!
0%
#258055000000
1!
1%
#258060000000
0!
0%
#258065000000
1!
1%
#258070000000
0!
0%
#258075000000
1!
1%
#258080000000
0!
0%
#258085000000
1!
1%
#258090000000
0!
0%
#258095000000
1!
1%
#258100000000
0!
0%
#258105000000
1!
1%
#258110000000
0!
0%
#258115000000
1!
1%
#258120000000
0!
0%
#258125000000
1!
1%
#258130000000
0!
0%
#258135000000
1!
1%
#258140000000
0!
0%
#258145000000
1!
1%
#258150000000
0!
0%
#258155000000
1!
1%
#258160000000
0!
0%
#258165000000
1!
1%
#258170000000
0!
0%
#258175000000
1!
1%
#258180000000
0!
0%
#258185000000
1!
1%
#258190000000
0!
0%
#258195000000
1!
1%
#258200000000
0!
0%
#258205000000
1!
1%
#258210000000
0!
0%
#258215000000
1!
1%
#258220000000
0!
0%
#258225000000
1!
1%
#258230000000
0!
0%
#258235000000
1!
1%
#258240000000
0!
0%
#258245000000
1!
1%
#258250000000
0!
0%
#258255000000
1!
1%
#258260000000
0!
0%
#258265000000
1!
1%
#258270000000
0!
0%
#258275000000
1!
1%
#258280000000
0!
0%
#258285000000
1!
1%
#258290000000
0!
0%
#258295000000
1!
1%
#258300000000
0!
0%
#258305000000
1!
1%
#258310000000
0!
0%
#258315000000
1!
1%
#258320000000
0!
0%
#258325000000
1!
1%
#258330000000
0!
0%
#258335000000
1!
1%
#258340000000
0!
0%
#258345000000
1!
1%
#258350000000
0!
0%
#258355000000
1!
1%
#258360000000
0!
0%
#258365000000
1!
1%
#258370000000
0!
0%
#258375000000
1!
1%
#258380000000
0!
0%
#258385000000
1!
1%
#258390000000
0!
0%
#258395000000
1!
1%
#258400000000
0!
0%
#258405000000
1!
1%
#258410000000
0!
0%
#258415000000
1!
1%
#258420000000
0!
0%
#258425000000
1!
1%
#258430000000
0!
0%
#258435000000
1!
1%
#258440000000
0!
0%
#258445000000
1!
1%
#258450000000
0!
0%
#258455000000
1!
1%
#258460000000
0!
0%
#258465000000
1!
1%
#258470000000
0!
0%
#258475000000
1!
1%
#258480000000
0!
0%
#258485000000
1!
1%
#258490000000
0!
0%
#258495000000
1!
1%
#258500000000
0!
0%
#258505000000
1!
1%
#258510000000
0!
0%
#258515000000
1!
1%
#258520000000
0!
0%
#258525000000
1!
1%
#258530000000
0!
0%
#258535000000
1!
1%
#258540000000
0!
0%
#258545000000
1!
1%
#258550000000
0!
0%
#258555000000
1!
1%
#258560000000
0!
0%
#258565000000
1!
1%
#258570000000
0!
0%
#258575000000
1!
1%
#258580000000
0!
0%
#258585000000
1!
1%
#258590000000
0!
0%
#258595000000
1!
1%
#258600000000
0!
0%
#258605000000
1!
1%
#258610000000
0!
0%
#258615000000
1!
1%
#258620000000
0!
0%
#258625000000
1!
1%
#258630000000
0!
0%
#258635000000
1!
1%
#258640000000
0!
0%
#258645000000
1!
1%
#258650000000
0!
0%
#258655000000
1!
1%
#258660000000
0!
0%
#258665000000
1!
1%
#258670000000
0!
0%
#258675000000
1!
1%
#258680000000
0!
0%
#258685000000
1!
1%
#258690000000
0!
0%
#258695000000
1!
1%
#258700000000
0!
0%
#258705000000
1!
1%
#258710000000
0!
0%
#258715000000
1!
1%
#258720000000
0!
0%
#258725000000
1!
1%
#258730000000
0!
0%
#258735000000
1!
1%
#258740000000
0!
0%
#258745000000
1!
1%
#258750000000
0!
0%
#258755000000
1!
1%
#258760000000
0!
0%
#258765000000
1!
1%
#258770000000
0!
0%
#258775000000
1!
1%
#258780000000
0!
0%
#258785000000
1!
1%
#258790000000
0!
0%
#258795000000
1!
1%
#258800000000
0!
0%
#258805000000
1!
1%
#258810000000
0!
0%
#258815000000
1!
1%
#258820000000
0!
0%
#258825000000
1!
1%
#258830000000
0!
0%
#258835000000
1!
1%
#258840000000
0!
0%
#258845000000
1!
1%
#258850000000
0!
0%
#258855000000
1!
1%
#258860000000
0!
0%
#258865000000
1!
1%
#258870000000
0!
0%
#258875000000
1!
1%
#258880000000
0!
0%
#258885000000
1!
1%
#258890000000
0!
0%
#258895000000
1!
1%
#258900000000
0!
0%
#258905000000
1!
1%
#258910000000
0!
0%
#258915000000
1!
1%
#258920000000
0!
0%
#258925000000
1!
1%
#258930000000
0!
0%
#258935000000
1!
1%
#258940000000
0!
0%
#258945000000
1!
1%
#258950000000
0!
0%
#258955000000
1!
1%
#258960000000
0!
0%
#258965000000
1!
1%
#258970000000
0!
0%
#258975000000
1!
1%
#258980000000
0!
0%
#258985000000
1!
1%
#258990000000
0!
0%
#258995000000
1!
1%
#259000000000
0!
0%
#259005000000
1!
1%
#259010000000
0!
0%
#259015000000
1!
1%
#259020000000
0!
0%
#259025000000
1!
1%
#259030000000
0!
0%
#259035000000
1!
1%
#259040000000
0!
0%
#259045000000
1!
1%
#259050000000
0!
0%
#259055000000
1!
1%
#259060000000
0!
0%
#259065000000
1!
1%
#259070000000
0!
0%
#259075000000
1!
1%
#259080000000
0!
0%
#259085000000
1!
1%
#259090000000
0!
0%
#259095000000
1!
1%
#259100000000
0!
0%
#259105000000
1!
1%
#259110000000
0!
0%
#259115000000
1!
1%
#259120000000
0!
0%
#259125000000
1!
1%
#259130000000
0!
0%
#259135000000
1!
1%
#259140000000
0!
0%
#259145000000
1!
1%
#259150000000
0!
0%
#259155000000
1!
1%
#259160000000
0!
0%
#259165000000
1!
1%
#259170000000
0!
0%
#259175000000
1!
1%
#259180000000
0!
0%
#259185000000
1!
1%
#259190000000
0!
0%
#259195000000
1!
1%
#259200000000
0!
0%
#259205000000
1!
1%
#259210000000
0!
0%
#259215000000
1!
1%
#259220000000
0!
0%
#259225000000
1!
1%
#259230000000
0!
0%
#259235000000
1!
1%
#259240000000
0!
0%
#259245000000
1!
1%
#259250000000
0!
0%
#259255000000
1!
1%
#259260000000
0!
0%
#259265000000
1!
1%
#259270000000
0!
0%
#259275000000
1!
1%
#259280000000
0!
0%
#259285000000
1!
1%
#259290000000
0!
0%
#259295000000
1!
1%
#259300000000
0!
0%
#259305000000
1!
1%
#259310000000
0!
0%
#259315000000
1!
1%
#259320000000
0!
0%
#259325000000
1!
1%
#259330000000
0!
0%
#259335000000
1!
1%
#259340000000
0!
0%
#259345000000
1!
1%
#259350000000
0!
0%
#259355000000
1!
1%
#259360000000
0!
0%
#259365000000
1!
1%
#259370000000
0!
0%
#259375000000
1!
1%
#259380000000
0!
0%
#259385000000
1!
1%
#259390000000
0!
0%
#259395000000
1!
1%
#259400000000
0!
0%
#259405000000
1!
1%
#259410000000
0!
0%
#259415000000
1!
1%
#259420000000
0!
0%
#259425000000
1!
1%
#259430000000
0!
0%
#259435000000
1!
1%
#259440000000
0!
0%
#259445000000
1!
1%
#259450000000
0!
0%
#259455000000
1!
1%
#259460000000
0!
0%
#259465000000
1!
1%
#259470000000
0!
0%
#259475000000
1!
1%
#259480000000
0!
0%
#259485000000
1!
1%
#259490000000
0!
0%
#259495000000
1!
1%
#259500000000
0!
0%
#259505000000
1!
1%
#259510000000
0!
0%
#259515000000
1!
1%
#259520000000
0!
0%
#259525000000
1!
1%
#259530000000
0!
0%
#259535000000
1!
1%
#259540000000
0!
0%
#259545000000
1!
1%
#259550000000
0!
0%
#259555000000
1!
1%
#259560000000
0!
0%
#259565000000
1!
1%
#259570000000
0!
0%
#259575000000
1!
1%
#259580000000
0!
0%
#259585000000
1!
1%
#259590000000
0!
0%
#259595000000
1!
1%
#259600000000
0!
0%
#259605000000
1!
1%
#259610000000
0!
0%
#259615000000
1!
1%
#259620000000
0!
0%
#259625000000
1!
1%
#259630000000
0!
0%
#259635000000
1!
1%
#259640000000
0!
0%
#259645000000
1!
1%
#259650000000
0!
0%
#259655000000
1!
1%
#259660000000
0!
0%
#259665000000
1!
1%
#259670000000
0!
0%
#259675000000
1!
1%
#259680000000
0!
0%
#259685000000
1!
1%
#259690000000
0!
0%
#259695000000
1!
1%
#259700000000
0!
0%
#259705000000
1!
1%
#259710000000
0!
0%
#259715000000
1!
1%
#259720000000
0!
0%
#259725000000
1!
1%
#259730000000
0!
0%
#259735000000
1!
1%
#259740000000
0!
0%
#259745000000
1!
1%
#259750000000
0!
0%
#259755000000
1!
1%
#259760000000
0!
0%
#259765000000
1!
1%
#259770000000
0!
0%
#259775000000
1!
1%
#259780000000
0!
0%
#259785000000
1!
1%
#259790000000
0!
0%
#259795000000
1!
1%
#259800000000
0!
0%
#259805000000
1!
1%
#259810000000
0!
0%
#259815000000
1!
1%
#259820000000
0!
0%
#259825000000
1!
1%
#259830000000
0!
0%
#259835000000
1!
1%
#259840000000
0!
0%
#259845000000
1!
1%
#259850000000
0!
0%
#259855000000
1!
1%
#259860000000
0!
0%
#259865000000
1!
1%
#259870000000
0!
0%
#259875000000
1!
1%
#259880000000
0!
0%
#259885000000
1!
1%
#259890000000
0!
0%
#259895000000
1!
1%
#259900000000
0!
0%
#259905000000
1!
1%
#259910000000
0!
0%
#259915000000
1!
1%
#259920000000
0!
0%
#259925000000
1!
1%
#259930000000
0!
0%
#259935000000
1!
1%
#259940000000
0!
0%
#259945000000
1!
1%
#259950000000
0!
0%
#259955000000
1!
1%
#259960000000
0!
0%
#259965000000
1!
1%
#259970000000
0!
0%
#259975000000
1!
1%
#259980000000
0!
0%
#259985000000
1!
1%
#259990000000
0!
0%
#259995000000
1!
1%
#260000000000
0!
0%
#260005000000
1!
1%
#260010000000
0!
0%
#260015000000
1!
1%
#260020000000
0!
0%
#260025000000
1!
1%
#260030000000
0!
0%
#260035000000
1!
1%
#260040000000
0!
0%
#260045000000
1!
1%
#260050000000
0!
0%
#260055000000
1!
1%
#260060000000
0!
0%
#260065000000
1!
1%
#260070000000
0!
0%
#260075000000
1!
1%
#260080000000
0!
0%
#260085000000
1!
1%
#260090000000
0!
0%
#260095000000
1!
1%
#260100000000
0!
0%
#260105000000
1!
1%
#260110000000
0!
0%
#260115000000
1!
1%
#260120000000
0!
0%
#260125000000
1!
1%
#260130000000
0!
0%
#260135000000
1!
1%
#260140000000
0!
0%
#260145000000
1!
1%
#260150000000
0!
0%
#260155000000
1!
1%
#260160000000
0!
0%
#260165000000
1!
1%
#260170000000
0!
0%
#260175000000
1!
1%
#260180000000
0!
0%
#260185000000
1!
1%
#260190000000
0!
0%
#260195000000
1!
1%
#260200000000
0!
0%
#260205000000
1!
1%
#260210000000
0!
0%
#260215000000
1!
1%
#260220000000
0!
0%
#260225000000
1!
1%
#260230000000
0!
0%
#260235000000
1!
1%
#260240000000
0!
0%
#260245000000
1!
1%
#260250000000
0!
0%
#260255000000
1!
1%
#260260000000
0!
0%
#260265000000
1!
1%
#260270000000
0!
0%
#260275000000
1!
1%
#260280000000
0!
0%
#260285000000
1!
1%
#260290000000
0!
0%
#260295000000
1!
1%
#260300000000
0!
0%
#260305000000
1!
1%
#260310000000
0!
0%
#260315000000
1!
1%
#260320000000
0!
0%
#260325000000
1!
1%
#260330000000
0!
0%
#260335000000
1!
1%
#260340000000
0!
0%
#260345000000
1!
1%
#260350000000
0!
0%
#260355000000
1!
1%
#260360000000
0!
0%
#260365000000
1!
1%
#260370000000
0!
0%
#260375000000
1!
1%
#260380000000
0!
0%
#260385000000
1!
1%
#260390000000
0!
0%
#260395000000
1!
1%
#260400000000
0!
0%
#260405000000
1!
1%
#260410000000
0!
0%
#260415000000
1!
1%
#260420000000
0!
0%
#260425000000
1!
1%
#260430000000
0!
0%
#260435000000
1!
1%
#260440000000
0!
0%
#260445000000
1!
1%
#260450000000
0!
0%
#260455000000
1!
1%
#260460000000
0!
0%
#260465000000
1!
1%
#260470000000
0!
0%
#260475000000
1!
1%
#260480000000
0!
0%
#260485000000
1!
1%
#260490000000
0!
0%
#260495000000
1!
1%
#260500000000
0!
0%
#260505000000
1!
1%
#260510000000
0!
0%
#260515000000
1!
1%
#260520000000
0!
0%
#260525000000
1!
1%
#260530000000
0!
0%
#260535000000
1!
1%
#260540000000
0!
0%
#260545000000
1!
1%
#260550000000
0!
0%
#260555000000
1!
1%
#260560000000
0!
0%
#260565000000
1!
1%
#260570000000
0!
0%
#260575000000
1!
1%
#260580000000
0!
0%
#260585000000
1!
1%
#260590000000
0!
0%
#260595000000
1!
1%
#260600000000
0!
0%
#260605000000
1!
1%
#260610000000
0!
0%
#260615000000
1!
1%
#260620000000
0!
0%
#260625000000
1!
1%
#260630000000
0!
0%
#260635000000
1!
1%
#260640000000
0!
0%
#260645000000
1!
1%
#260650000000
0!
0%
#260655000000
1!
1%
#260660000000
0!
0%
#260665000000
1!
1%
#260670000000
0!
0%
#260675000000
1!
1%
#260680000000
0!
0%
#260685000000
1!
1%
#260690000000
0!
0%
#260695000000
1!
1%
#260700000000
0!
0%
#260705000000
1!
1%
#260710000000
0!
0%
#260715000000
1!
1%
#260720000000
0!
0%
#260725000000
1!
1%
#260730000000
0!
0%
#260735000000
1!
1%
#260740000000
0!
0%
#260745000000
1!
1%
#260750000000
0!
0%
#260755000000
1!
1%
#260760000000
0!
0%
#260765000000
1!
1%
#260770000000
0!
0%
#260775000000
1!
1%
#260780000000
0!
0%
#260785000000
1!
1%
#260790000000
0!
0%
#260795000000
1!
1%
#260800000000
0!
0%
#260805000000
1!
1%
#260810000000
0!
0%
#260815000000
1!
1%
#260820000000
0!
0%
#260825000000
1!
1%
#260830000000
0!
0%
#260835000000
1!
1%
#260840000000
0!
0%
#260845000000
1!
1%
#260850000000
0!
0%
#260855000000
1!
1%
#260860000000
0!
0%
#260865000000
1!
1%
#260870000000
0!
0%
#260875000000
1!
1%
#260880000000
0!
0%
#260885000000
1!
1%
#260890000000
0!
0%
#260895000000
1!
1%
#260900000000
0!
0%
#260905000000
1!
1%
#260910000000
0!
0%
#260915000000
1!
1%
#260920000000
0!
0%
#260925000000
1!
1%
#260930000000
0!
0%
#260935000000
1!
1%
#260940000000
0!
0%
#260945000000
1!
1%
#260950000000
0!
0%
#260955000000
1!
1%
#260960000000
0!
0%
#260965000000
1!
1%
#260970000000
0!
0%
#260975000000
1!
1%
#260980000000
0!
0%
#260985000000
1!
1%
#260990000000
0!
0%
#260995000000
1!
1%
#261000000000
0!
0%
#261005000000
1!
1%
#261010000000
0!
0%
#261015000000
1!
1%
#261020000000
0!
0%
#261025000000
1!
1%
#261030000000
0!
0%
#261035000000
1!
1%
#261040000000
0!
0%
#261045000000
1!
1%
#261050000000
0!
0%
#261055000000
1!
1%
#261060000000
0!
0%
#261065000000
1!
1%
#261070000000
0!
0%
#261075000000
1!
1%
#261080000000
0!
0%
#261085000000
1!
1%
#261090000000
0!
0%
#261095000000
1!
1%
#261100000000
0!
0%
#261105000000
1!
1%
#261110000000
0!
0%
#261115000000
1!
1%
#261120000000
0!
0%
#261125000000
1!
1%
#261130000000
0!
0%
#261135000000
1!
1%
#261140000000
0!
0%
#261145000000
1!
1%
#261150000000
0!
0%
#261155000000
1!
1%
#261160000000
0!
0%
#261165000000
1!
1%
#261170000000
0!
0%
#261175000000
1!
1%
#261180000000
0!
0%
#261185000000
1!
1%
#261190000000
0!
0%
#261195000000
1!
1%
#261200000000
0!
0%
#261205000000
1!
1%
#261210000000
0!
0%
#261215000000
1!
1%
#261220000000
0!
0%
#261225000000
1!
1%
#261230000000
0!
0%
#261235000000
1!
1%
#261240000000
0!
0%
#261245000000
1!
1%
#261250000000
0!
0%
#261255000000
1!
1%
#261260000000
0!
0%
#261265000000
1!
1%
#261270000000
0!
0%
#261275000000
1!
1%
#261280000000
0!
0%
#261285000000
1!
1%
#261290000000
0!
0%
#261295000000
1!
1%
#261300000000
0!
0%
#261305000000
1!
1%
#261310000000
0!
0%
#261315000000
1!
1%
#261320000000
0!
0%
#261325000000
1!
1%
#261330000000
0!
0%
#261335000000
1!
1%
#261340000000
0!
0%
#261345000000
1!
1%
#261350000000
0!
0%
#261355000000
1!
1%
#261360000000
0!
0%
#261365000000
1!
1%
#261370000000
0!
0%
#261375000000
1!
1%
#261380000000
0!
0%
#261385000000
1!
1%
#261390000000
0!
0%
#261395000000
1!
1%
#261400000000
0!
0%
#261405000000
1!
1%
#261410000000
0!
0%
#261415000000
1!
1%
#261420000000
0!
0%
#261425000000
1!
1%
#261430000000
0!
0%
#261435000000
1!
1%
#261440000000
0!
0%
#261445000000
1!
1%
#261450000000
0!
0%
#261455000000
1!
1%
#261460000000
0!
0%
#261465000000
1!
1%
#261470000000
0!
0%
#261475000000
1!
1%
#261480000000
0!
0%
#261485000000
1!
1%
#261490000000
0!
0%
#261495000000
1!
1%
#261500000000
0!
0%
#261505000000
1!
1%
#261510000000
0!
0%
#261515000000
1!
1%
#261520000000
0!
0%
#261525000000
1!
1%
#261530000000
0!
0%
#261535000000
1!
1%
#261540000000
0!
0%
#261545000000
1!
1%
#261550000000
0!
0%
#261555000000
1!
1%
#261560000000
0!
0%
#261565000000
1!
1%
#261570000000
0!
0%
#261575000000
1!
1%
#261580000000
0!
0%
#261585000000
1!
1%
#261590000000
0!
0%
#261595000000
1!
1%
#261600000000
0!
0%
#261605000000
1!
1%
#261610000000
0!
0%
#261615000000
1!
1%
#261620000000
0!
0%
#261625000000
1!
1%
#261630000000
0!
0%
#261635000000
1!
1%
#261640000000
0!
0%
#261645000000
1!
1%
#261650000000
0!
0%
#261655000000
1!
1%
#261660000000
0!
0%
#261665000000
1!
1%
#261670000000
0!
0%
#261675000000
1!
1%
#261680000000
0!
0%
#261685000000
1!
1%
#261690000000
0!
0%
#261695000000
1!
1%
#261700000000
0!
0%
#261705000000
1!
1%
#261710000000
0!
0%
#261715000000
1!
1%
#261720000000
0!
0%
#261725000000
1!
1%
#261730000000
0!
0%
#261735000000
1!
1%
#261740000000
0!
0%
#261745000000
1!
1%
#261750000000
0!
0%
#261755000000
1!
1%
#261760000000
0!
0%
#261765000000
1!
1%
#261770000000
0!
0%
#261775000000
1!
1%
#261780000000
0!
0%
#261785000000
1!
1%
#261790000000
0!
0%
#261795000000
1!
1%
#261800000000
0!
0%
#261805000000
1!
1%
#261810000000
0!
0%
#261815000000
1!
1%
#261820000000
0!
0%
#261825000000
1!
1%
#261830000000
0!
0%
#261835000000
1!
1%
#261840000000
0!
0%
#261845000000
1!
1%
#261850000000
0!
0%
#261855000000
1!
1%
#261860000000
0!
0%
#261865000000
1!
1%
#261870000000
0!
0%
#261875000000
1!
1%
#261880000000
0!
0%
#261885000000
1!
1%
#261890000000
0!
0%
#261895000000
1!
1%
#261900000000
0!
0%
#261905000000
1!
1%
#261910000000
0!
0%
#261915000000
1!
1%
#261920000000
0!
0%
#261925000000
1!
1%
#261930000000
0!
0%
#261935000000
1!
1%
#261940000000
0!
0%
#261945000000
1!
1%
#261950000000
0!
0%
#261955000000
1!
1%
#261960000000
0!
0%
#261965000000
1!
1%
#261970000000
0!
0%
#261975000000
1!
1%
#261980000000
0!
0%
#261985000000
1!
1%
#261990000000
0!
0%
#261995000000
1!
1%
#262000000000
0!
0%
#262005000000
1!
1%
#262010000000
0!
0%
#262015000000
1!
1%
#262020000000
0!
0%
#262025000000
1!
1%
#262030000000
0!
0%
#262035000000
1!
1%
#262040000000
0!
0%
#262045000000
1!
1%
#262050000000
0!
0%
#262055000000
1!
1%
#262060000000
0!
0%
#262065000000
1!
1%
#262070000000
0!
0%
#262075000000
1!
1%
#262080000000
0!
0%
#262085000000
1!
1%
#262090000000
0!
0%
#262095000000
1!
1%
#262100000000
0!
0%
#262105000000
1!
1%
#262110000000
0!
0%
#262115000000
1!
1%
#262120000000
0!
0%
#262125000000
1!
1%
#262130000000
0!
0%
#262135000000
1!
1%
#262140000000
0!
0%
#262145000000
1!
1%
#262150000000
0!
0%
#262155000000
1!
1%
#262160000000
0!
0%
#262165000000
1!
1%
#262170000000
0!
0%
#262175000000
1!
1%
#262180000000
0!
0%
#262185000000
1!
1%
#262190000000
0!
0%
#262195000000
1!
1%
#262200000000
0!
0%
#262205000000
1!
1%
#262210000000
0!
0%
#262215000000
1!
1%
#262220000000
0!
0%
#262225000000
1!
1%
#262230000000
0!
0%
#262235000000
1!
1%
#262240000000
0!
0%
#262245000000
1!
1%
#262250000000
0!
0%
#262255000000
1!
1%
#262260000000
0!
0%
#262265000000
1!
1%
#262270000000
0!
0%
#262275000000
1!
1%
#262280000000
0!
0%
#262285000000
1!
1%
#262290000000
0!
0%
#262295000000
1!
1%
#262300000000
0!
0%
#262305000000
1!
1%
#262310000000
0!
0%
#262315000000
1!
1%
#262320000000
0!
0%
#262325000000
1!
1%
#262330000000
0!
0%
#262335000000
1!
1%
#262340000000
0!
0%
#262345000000
1!
1%
#262350000000
0!
0%
#262355000000
1!
1%
#262360000000
0!
0%
#262365000000
1!
1%
#262370000000
0!
0%
#262375000000
1!
1%
#262380000000
0!
0%
#262385000000
1!
1%
#262390000000
0!
0%
#262395000000
1!
1%
#262400000000
0!
0%
#262405000000
1!
1%
#262410000000
0!
0%
#262415000000
1!
1%
#262420000000
0!
0%
#262425000000
1!
1%
#262430000000
0!
0%
#262435000000
1!
1%
#262440000000
0!
0%
#262445000000
1!
1%
#262450000000
0!
0%
#262455000000
1!
1%
#262460000000
0!
0%
#262465000000
1!
1%
#262470000000
0!
0%
#262475000000
1!
1%
#262480000000
0!
0%
#262485000000
1!
1%
#262490000000
0!
0%
#262495000000
1!
1%
#262500000000
0!
0%
#262505000000
1!
1%
#262510000000
0!
0%
#262515000000
1!
1%
#262520000000
0!
0%
#262525000000
1!
1%
#262530000000
0!
0%
#262535000000
1!
1%
#262540000000
0!
0%
#262545000000
1!
1%
#262550000000
0!
0%
#262555000000
1!
1%
#262560000000
0!
0%
#262565000000
1!
1%
#262570000000
0!
0%
#262575000000
1!
1%
#262580000000
0!
0%
#262585000000
1!
1%
#262590000000
0!
0%
#262595000000
1!
1%
#262600000000
0!
0%
#262605000000
1!
1%
#262610000000
0!
0%
#262615000000
1!
1%
#262620000000
0!
0%
#262625000000
1!
1%
#262630000000
0!
0%
#262635000000
1!
1%
#262640000000
0!
0%
#262645000000
1!
1%
#262650000000
0!
0%
#262655000000
1!
1%
#262660000000
0!
0%
#262665000000
1!
1%
#262670000000
0!
0%
#262675000000
1!
1%
#262680000000
0!
0%
#262685000000
1!
1%
#262690000000
0!
0%
#262695000000
1!
1%
#262700000000
0!
0%
#262705000000
1!
1%
#262710000000
0!
0%
#262715000000
1!
1%
#262720000000
0!
0%
#262725000000
1!
1%
#262730000000
0!
0%
#262735000000
1!
1%
#262740000000
0!
0%
#262745000000
1!
1%
#262750000000
0!
0%
#262755000000
1!
1%
#262760000000
0!
0%
#262765000000
1!
1%
#262770000000
0!
0%
#262775000000
1!
1%
#262780000000
0!
0%
#262785000000
1!
1%
#262790000000
0!
0%
#262795000000
1!
1%
#262800000000
0!
0%
#262805000000
1!
1%
#262810000000
0!
0%
#262815000000
1!
1%
#262820000000
0!
0%
#262825000000
1!
1%
#262830000000
0!
0%
#262835000000
1!
1%
#262840000000
0!
0%
#262845000000
1!
1%
#262850000000
0!
0%
#262855000000
1!
1%
#262860000000
0!
0%
#262865000000
1!
1%
#262870000000
0!
0%
#262875000000
1!
1%
#262880000000
0!
0%
#262885000000
1!
1%
#262890000000
0!
0%
#262895000000
1!
1%
#262900000000
0!
0%
#262905000000
1!
1%
#262910000000
0!
0%
#262915000000
1!
1%
#262920000000
0!
0%
#262925000000
1!
1%
#262930000000
0!
0%
#262935000000
1!
1%
#262940000000
0!
0%
#262945000000
1!
1%
#262950000000
0!
0%
#262955000000
1!
1%
#262960000000
0!
0%
#262965000000
1!
1%
#262970000000
0!
0%
#262975000000
1!
1%
#262980000000
0!
0%
#262985000000
1!
1%
#262990000000
0!
0%
#262995000000
1!
1%
#263000000000
0!
0%
#263005000000
1!
1%
#263010000000
0!
0%
#263015000000
1!
1%
#263020000000
0!
0%
#263025000000
1!
1%
#263030000000
0!
0%
#263035000000
1!
1%
#263040000000
0!
0%
#263045000000
1!
1%
#263050000000
0!
0%
#263055000000
1!
1%
#263060000000
0!
0%
#263065000000
1!
1%
#263070000000
0!
0%
#263075000000
1!
1%
#263080000000
0!
0%
#263085000000
1!
1%
#263090000000
0!
0%
#263095000000
1!
1%
#263100000000
0!
0%
#263105000000
1!
1%
#263110000000
0!
0%
#263115000000
1!
1%
#263120000000
0!
0%
#263125000000
1!
1%
#263130000000
0!
0%
#263135000000
1!
1%
#263140000000
0!
0%
#263145000000
1!
1%
#263150000000
0!
0%
#263155000000
1!
1%
#263160000000
0!
0%
#263165000000
1!
1%
#263170000000
0!
0%
#263175000000
1!
1%
#263180000000
0!
0%
#263185000000
1!
1%
#263190000000
0!
0%
#263195000000
1!
1%
#263200000000
0!
0%
#263205000000
1!
1%
#263210000000
0!
0%
#263215000000
1!
1%
#263220000000
0!
0%
#263225000000
1!
1%
#263230000000
0!
0%
#263235000000
1!
1%
#263240000000
0!
0%
#263245000000
1!
1%
#263250000000
0!
0%
#263255000000
1!
1%
#263260000000
0!
0%
#263265000000
1!
1%
#263270000000
0!
0%
#263275000000
1!
1%
#263280000000
0!
0%
#263285000000
1!
1%
#263290000000
0!
0%
#263295000000
1!
1%
#263300000000
0!
0%
#263305000000
1!
1%
#263310000000
0!
0%
#263315000000
1!
1%
#263320000000
0!
0%
#263325000000
1!
1%
#263330000000
0!
0%
#263335000000
1!
1%
#263340000000
0!
0%
#263345000000
1!
1%
#263350000000
0!
0%
#263355000000
1!
1%
#263360000000
0!
0%
#263365000000
1!
1%
#263370000000
0!
0%
#263375000000
1!
1%
#263380000000
0!
0%
#263385000000
1!
1%
#263390000000
0!
0%
#263395000000
1!
1%
#263400000000
0!
0%
#263405000000
1!
1%
#263410000000
0!
0%
#263415000000
1!
1%
#263420000000
0!
0%
#263425000000
1!
1%
#263430000000
0!
0%
#263435000000
1!
1%
#263440000000
0!
0%
#263445000000
1!
1%
#263450000000
0!
0%
#263455000000
1!
1%
#263460000000
0!
0%
#263465000000
1!
1%
#263470000000
0!
0%
#263475000000
1!
1%
#263480000000
0!
0%
#263485000000
1!
1%
#263490000000
0!
0%
#263495000000
1!
1%
#263500000000
0!
0%
#263505000000
1!
1%
#263510000000
0!
0%
#263515000000
1!
1%
#263520000000
0!
0%
#263525000000
1!
1%
#263530000000
0!
0%
#263535000000
1!
1%
#263540000000
0!
0%
#263545000000
1!
1%
#263550000000
0!
0%
#263555000000
1!
1%
#263560000000
0!
0%
#263565000000
1!
1%
#263570000000
0!
0%
#263575000000
1!
1%
#263580000000
0!
0%
#263585000000
1!
1%
#263590000000
0!
0%
#263595000000
1!
1%
#263600000000
0!
0%
#263605000000
1!
1%
#263610000000
0!
0%
#263615000000
1!
1%
#263620000000
0!
0%
#263625000000
1!
1%
#263630000000
0!
0%
#263635000000
1!
1%
#263640000000
0!
0%
#263645000000
1!
1%
#263650000000
0!
0%
#263655000000
1!
1%
#263660000000
0!
0%
#263665000000
1!
1%
#263670000000
0!
0%
#263675000000
1!
1%
#263680000000
0!
0%
#263685000000
1!
1%
#263690000000
0!
0%
#263695000000
1!
1%
#263700000000
0!
0%
#263705000000
1!
1%
#263710000000
0!
0%
#263715000000
1!
1%
#263720000000
0!
0%
#263725000000
1!
1%
#263730000000
0!
0%
#263735000000
1!
1%
#263740000000
0!
0%
#263745000000
1!
1%
#263750000000
0!
0%
#263755000000
1!
1%
#263760000000
0!
0%
#263765000000
1!
1%
#263770000000
0!
0%
#263775000000
1!
1%
#263780000000
0!
0%
#263785000000
1!
1%
#263790000000
0!
0%
#263795000000
1!
1%
#263800000000
0!
0%
#263805000000
1!
1%
#263810000000
0!
0%
#263815000000
1!
1%
#263820000000
0!
0%
#263825000000
1!
1%
#263830000000
0!
0%
#263835000000
1!
1%
#263840000000
0!
0%
#263845000000
1!
1%
#263850000000
0!
0%
#263855000000
1!
1%
#263860000000
0!
0%
#263865000000
1!
1%
#263870000000
0!
0%
#263875000000
1!
1%
#263880000000
0!
0%
#263885000000
1!
1%
#263890000000
0!
0%
#263895000000
1!
1%
#263900000000
0!
0%
#263905000000
1!
1%
#263910000000
0!
0%
#263915000000
1!
1%
#263920000000
0!
0%
#263925000000
1!
1%
#263930000000
0!
0%
#263935000000
1!
1%
#263940000000
0!
0%
#263945000000
1!
1%
#263950000000
0!
0%
#263955000000
1!
1%
#263960000000
0!
0%
#263965000000
1!
1%
#263970000000
0!
0%
#263975000000
1!
1%
#263980000000
0!
0%
#263985000000
1!
1%
#263990000000
0!
0%
#263995000000
1!
1%
#264000000000
0!
0%
#264005000000
1!
1%
#264010000000
0!
0%
#264015000000
1!
1%
#264020000000
0!
0%
#264025000000
1!
1%
#264030000000
0!
0%
#264035000000
1!
1%
#264040000000
0!
0%
#264045000000
1!
1%
#264050000000
0!
0%
#264055000000
1!
1%
#264060000000
0!
0%
#264065000000
1!
1%
#264070000000
0!
0%
#264075000000
1!
1%
#264080000000
0!
0%
#264085000000
1!
1%
#264090000000
0!
0%
#264095000000
1!
1%
#264100000000
0!
0%
#264105000000
1!
1%
#264110000000
0!
0%
#264115000000
1!
1%
#264120000000
0!
0%
#264125000000
1!
1%
#264130000000
0!
0%
#264135000000
1!
1%
#264140000000
0!
0%
#264145000000
1!
1%
#264150000000
0!
0%
#264155000000
1!
1%
#264160000000
0!
0%
#264165000000
1!
1%
#264170000000
0!
0%
#264175000000
1!
1%
#264180000000
0!
0%
#264185000000
1!
1%
#264190000000
0!
0%
#264195000000
1!
1%
#264200000000
0!
0%
#264205000000
1!
1%
#264210000000
0!
0%
#264215000000
1!
1%
#264220000000
0!
0%
#264225000000
1!
1%
#264230000000
0!
0%
#264235000000
1!
1%
#264240000000
0!
0%
#264245000000
1!
1%
#264250000000
0!
0%
#264255000000
1!
1%
#264260000000
0!
0%
#264265000000
1!
1%
#264270000000
0!
0%
#264275000000
1!
1%
#264280000000
0!
0%
#264285000000
1!
1%
#264290000000
0!
0%
#264295000000
1!
1%
#264300000000
0!
0%
#264305000000
1!
1%
#264310000000
0!
0%
#264315000000
1!
1%
#264320000000
0!
0%
#264325000000
1!
1%
#264330000000
0!
0%
#264335000000
1!
1%
#264340000000
0!
0%
#264345000000
1!
1%
#264350000000
0!
0%
#264355000000
1!
1%
#264360000000
0!
0%
#264365000000
1!
1%
#264370000000
0!
0%
#264375000000
1!
1%
#264380000000
0!
0%
#264385000000
1!
1%
#264390000000
0!
0%
#264395000000
1!
1%
#264400000000
0!
0%
#264405000000
1!
1%
#264410000000
0!
0%
#264415000000
1!
1%
#264420000000
0!
0%
#264425000000
1!
1%
#264430000000
0!
0%
#264435000000
1!
1%
#264440000000
0!
0%
#264445000000
1!
1%
#264450000000
0!
0%
#264455000000
1!
1%
#264460000000
0!
0%
#264465000000
1!
1%
#264470000000
0!
0%
#264475000000
1!
1%
#264480000000
0!
0%
#264485000000
1!
1%
#264490000000
0!
0%
#264495000000
1!
1%
#264500000000
0!
0%
#264505000000
1!
1%
#264510000000
0!
0%
#264515000000
1!
1%
#264520000000
0!
0%
#264525000000
1!
1%
#264530000000
0!
0%
#264535000000
1!
1%
#264540000000
0!
0%
#264545000000
1!
1%
#264550000000
0!
0%
#264555000000
1!
1%
#264560000000
0!
0%
#264565000000
1!
1%
#264570000000
0!
0%
#264575000000
1!
1%
#264580000000
0!
0%
#264585000000
1!
1%
#264590000000
0!
0%
#264595000000
1!
1%
#264600000000
0!
0%
#264605000000
1!
1%
#264610000000
0!
0%
#264615000000
1!
1%
#264620000000
0!
0%
#264625000000
1!
1%
#264630000000
0!
0%
#264635000000
1!
1%
#264640000000
0!
0%
#264645000000
1!
1%
#264650000000
0!
0%
#264655000000
1!
1%
#264660000000
0!
0%
#264665000000
1!
1%
#264670000000
0!
0%
#264675000000
1!
1%
#264680000000
0!
0%
#264685000000
1!
1%
#264690000000
0!
0%
#264695000000
1!
1%
#264700000000
0!
0%
#264705000000
1!
1%
#264710000000
0!
0%
#264715000000
1!
1%
#264720000000
0!
0%
#264725000000
1!
1%
#264730000000
0!
0%
#264735000000
1!
1%
#264740000000
0!
0%
#264745000000
1!
1%
#264750000000
0!
0%
#264755000000
1!
1%
#264760000000
0!
0%
#264765000000
1!
1%
#264770000000
0!
0%
#264775000000
1!
1%
#264780000000
0!
0%
#264785000000
1!
1%
#264790000000
0!
0%
#264795000000
1!
1%
#264800000000
0!
0%
#264805000000
1!
1%
#264810000000
0!
0%
#264815000000
1!
1%
#264820000000
0!
0%
#264825000000
1!
1%
#264830000000
0!
0%
#264835000000
1!
1%
#264840000000
0!
0%
#264845000000
1!
1%
#264850000000
0!
0%
#264855000000
1!
1%
#264860000000
0!
0%
#264865000000
1!
1%
#264870000000
0!
0%
#264875000000
1!
1%
#264880000000
0!
0%
#264885000000
1!
1%
#264890000000
0!
0%
#264895000000
1!
1%
#264900000000
0!
0%
#264905000000
1!
1%
#264910000000
0!
0%
#264915000000
1!
1%
#264920000000
0!
0%
#264925000000
1!
1%
#264930000000
0!
0%
#264935000000
1!
1%
#264940000000
0!
0%
#264945000000
1!
1%
#264950000000
0!
0%
#264955000000
1!
1%
#264960000000
0!
0%
#264965000000
1!
1%
#264970000000
0!
0%
#264975000000
1!
1%
#264980000000
0!
0%
#264985000000
1!
1%
#264990000000
0!
0%
#264995000000
1!
1%
#265000000000
0!
0%
#265005000000
1!
1%
#265010000000
0!
0%
#265015000000
1!
1%
#265020000000
0!
0%
#265025000000
1!
1%
#265030000000
0!
0%
#265035000000
1!
1%
#265040000000
0!
0%
#265045000000
1!
1%
#265050000000
0!
0%
#265055000000
1!
1%
#265060000000
0!
0%
#265065000000
1!
1%
#265070000000
0!
0%
#265075000000
1!
1%
#265080000000
0!
0%
#265085000000
1!
1%
#265090000000
0!
0%
#265095000000
1!
1%
#265100000000
0!
0%
#265105000000
1!
1%
#265110000000
0!
0%
#265115000000
1!
1%
#265120000000
0!
0%
#265125000000
1!
1%
#265130000000
0!
0%
#265135000000
1!
1%
#265140000000
0!
0%
#265145000000
1!
1%
#265150000000
0!
0%
#265155000000
1!
1%
#265160000000
0!
0%
#265165000000
1!
1%
#265170000000
0!
0%
#265175000000
1!
1%
#265180000000
0!
0%
#265185000000
1!
1%
#265190000000
0!
0%
#265195000000
1!
1%
#265200000000
0!
0%
#265205000000
1!
1%
#265210000000
0!
0%
#265215000000
1!
1%
#265220000000
0!
0%
#265225000000
1!
1%
#265230000000
0!
0%
#265235000000
1!
1%
#265240000000
0!
0%
#265245000000
1!
1%
#265250000000
0!
0%
#265255000000
1!
1%
#265260000000
0!
0%
#265265000000
1!
1%
#265270000000
0!
0%
#265275000000
1!
1%
#265280000000
0!
0%
#265285000000
1!
1%
#265290000000
0!
0%
#265295000000
1!
1%
#265300000000
0!
0%
#265305000000
1!
1%
#265310000000
0!
0%
#265315000000
1!
1%
#265320000000
0!
0%
#265325000000
1!
1%
#265330000000
0!
0%
#265335000000
1!
1%
#265340000000
0!
0%
#265345000000
1!
1%
#265350000000
0!
0%
#265355000000
1!
1%
#265360000000
0!
0%
#265365000000
1!
1%
#265370000000
0!
0%
#265375000000
1!
1%
#265380000000
0!
0%
#265385000000
1!
1%
#265390000000
0!
0%
#265395000000
1!
1%
#265400000000
0!
0%
#265405000000
1!
1%
#265410000000
0!
0%
#265415000000
1!
1%
#265420000000
0!
0%
#265425000000
1!
1%
#265430000000
0!
0%
#265435000000
1!
1%
#265440000000
0!
0%
#265445000000
1!
1%
#265450000000
0!
0%
#265455000000
1!
1%
#265460000000
0!
0%
#265465000000
1!
1%
#265470000000
0!
0%
#265475000000
1!
1%
#265480000000
0!
0%
#265485000000
1!
1%
#265490000000
0!
0%
#265495000000
1!
1%
#265500000000
0!
0%
#265505000000
1!
1%
#265510000000
0!
0%
#265515000000
1!
1%
#265520000000
0!
0%
#265525000000
1!
1%
#265530000000
0!
0%
#265535000000
1!
1%
#265540000000
0!
0%
#265545000000
1!
1%
#265550000000
0!
0%
#265555000000
1!
1%
#265560000000
0!
0%
#265565000000
1!
1%
#265570000000
0!
0%
#265575000000
1!
1%
#265580000000
0!
0%
#265585000000
1!
1%
#265590000000
0!
0%
#265595000000
1!
1%
#265600000000
0!
0%
#265605000000
1!
1%
#265610000000
0!
0%
#265615000000
1!
1%
#265620000000
0!
0%
#265625000000
1!
1%
#265630000000
0!
0%
#265635000000
1!
1%
#265640000000
0!
0%
#265645000000
1!
1%
#265650000000
0!
0%
#265655000000
1!
1%
#265660000000
0!
0%
#265665000000
1!
1%
#265670000000
0!
0%
#265675000000
1!
1%
#265680000000
0!
0%
#265685000000
1!
1%
#265690000000
0!
0%
#265695000000
1!
1%
#265700000000
0!
0%
#265705000000
1!
1%
#265710000000
0!
0%
#265715000000
1!
1%
#265720000000
0!
0%
#265725000000
1!
1%
#265730000000
0!
0%
#265735000000
1!
1%
#265740000000
0!
0%
#265745000000
1!
1%
#265750000000
0!
0%
#265755000000
1!
1%
#265760000000
0!
0%
#265765000000
1!
1%
#265770000000
0!
0%
#265775000000
1!
1%
#265780000000
0!
0%
#265785000000
1!
1%
#265790000000
0!
0%
#265795000000
1!
1%
#265800000000
0!
0%
#265805000000
1!
1%
#265810000000
0!
0%
#265815000000
1!
1%
#265820000000
0!
0%
#265825000000
1!
1%
#265830000000
0!
0%
#265835000000
1!
1%
#265840000000
0!
0%
#265845000000
1!
1%
#265850000000
0!
0%
#265855000000
1!
1%
#265860000000
0!
0%
#265865000000
1!
1%
#265870000000
0!
0%
#265875000000
1!
1%
#265880000000
0!
0%
#265885000000
1!
1%
#265890000000
0!
0%
#265895000000
1!
1%
#265900000000
0!
0%
#265905000000
1!
1%
#265910000000
0!
0%
#265915000000
1!
1%
#265920000000
0!
0%
#265925000000
1!
1%
#265930000000
0!
0%
#265935000000
1!
1%
#265940000000
0!
0%
#265945000000
1!
1%
#265950000000
0!
0%
#265955000000
1!
1%
#265960000000
0!
0%
#265965000000
1!
1%
#265970000000
0!
0%
#265975000000
1!
1%
#265980000000
0!
0%
#265985000000
1!
1%
#265990000000
0!
0%
#265995000000
1!
1%
#266000000000
0!
0%
#266005000000
1!
1%
#266010000000
0!
0%
#266015000000
1!
1%
#266020000000
0!
0%
#266025000000
1!
1%
#266030000000
0!
0%
#266035000000
1!
1%
#266040000000
0!
0%
#266045000000
1!
1%
#266050000000
0!
0%
#266055000000
1!
1%
#266060000000
0!
0%
#266065000000
1!
1%
#266070000000
0!
0%
#266075000000
1!
1%
#266080000000
0!
0%
#266085000000
1!
1%
#266090000000
0!
0%
#266095000000
1!
1%
#266100000000
0!
0%
#266105000000
1!
1%
#266110000000
0!
0%
#266115000000
1!
1%
#266120000000
0!
0%
#266125000000
1!
1%
#266130000000
0!
0%
#266135000000
1!
1%
#266140000000
0!
0%
#266145000000
1!
1%
#266150000000
0!
0%
#266155000000
1!
1%
#266160000000
0!
0%
#266165000000
1!
1%
#266170000000
0!
0%
#266175000000
1!
1%
#266180000000
0!
0%
#266185000000
1!
1%
#266190000000
0!
0%
#266195000000
1!
1%
#266200000000
0!
0%
#266205000000
1!
1%
#266210000000
0!
0%
#266215000000
1!
1%
#266220000000
0!
0%
#266225000000
1!
1%
#266230000000
0!
0%
#266235000000
1!
1%
#266240000000
0!
0%
#266245000000
1!
1%
#266250000000
0!
0%
#266255000000
1!
1%
#266260000000
0!
0%
#266265000000
1!
1%
#266270000000
0!
0%
#266275000000
1!
1%
#266280000000
0!
0%
#266285000000
1!
1%
#266290000000
0!
0%
#266295000000
1!
1%
#266300000000
0!
0%
#266305000000
1!
1%
#266310000000
0!
0%
#266315000000
1!
1%
#266320000000
0!
0%
#266325000000
1!
1%
#266330000000
0!
0%
#266335000000
1!
1%
#266340000000
0!
0%
#266345000000
1!
1%
#266350000000
0!
0%
#266355000000
1!
1%
#266360000000
0!
0%
#266365000000
1!
1%
#266370000000
0!
0%
#266375000000
1!
1%
#266380000000
0!
0%
#266385000000
1!
1%
#266390000000
0!
0%
#266395000000
1!
1%
#266400000000
0!
0%
#266405000000
1!
1%
#266410000000
0!
0%
#266415000000
1!
1%
#266420000000
0!
0%
#266425000000
1!
1%
#266430000000
0!
0%
#266435000000
1!
1%
#266440000000
0!
0%
#266445000000
1!
1%
#266450000000
0!
0%
#266455000000
1!
1%
#266460000000
0!
0%
#266465000000
1!
1%
#266470000000
0!
0%
#266475000000
1!
1%
#266480000000
0!
0%
#266485000000
1!
1%
#266490000000
0!
0%
#266495000000
1!
1%
#266500000000
0!
0%
#266505000000
1!
1%
#266510000000
0!
0%
#266515000000
1!
1%
#266520000000
0!
0%
#266525000000
1!
1%
#266530000000
0!
0%
#266535000000
1!
1%
#266540000000
0!
0%
#266545000000
1!
1%
#266550000000
0!
0%
#266555000000
1!
1%
#266560000000
0!
0%
#266565000000
1!
1%
#266570000000
0!
0%
#266575000000
1!
1%
#266580000000
0!
0%
#266585000000
1!
1%
#266590000000
0!
0%
#266595000000
1!
1%
#266600000000
0!
0%
#266605000000
1!
1%
#266610000000
0!
0%
#266615000000
1!
1%
#266620000000
0!
0%
#266625000000
1!
1%
#266630000000
0!
0%
#266635000000
1!
1%
#266640000000
0!
0%
#266645000000
1!
1%
#266650000000
0!
0%
#266655000000
1!
1%
#266660000000
0!
0%
#266665000000
1!
1%
#266670000000
0!
0%
#266675000000
1!
1%
#266680000000
0!
0%
#266685000000
1!
1%
#266690000000
0!
0%
#266695000000
1!
1%
#266700000000
0!
0%
#266705000000
1!
1%
#266710000000
0!
0%
#266715000000
1!
1%
#266720000000
0!
0%
#266725000000
1!
1%
#266730000000
0!
0%
#266735000000
1!
1%
#266740000000
0!
0%
#266745000000
1!
1%
#266750000000
0!
0%
#266755000000
1!
1%
#266760000000
0!
0%
#266765000000
1!
1%
#266770000000
0!
0%
#266775000000
1!
1%
#266780000000
0!
0%
#266785000000
1!
1%
#266790000000
0!
0%
#266795000000
1!
1%
#266800000000
0!
0%
#266805000000
1!
1%
#266810000000
0!
0%
#266815000000
1!
1%
#266820000000
0!
0%
#266825000000
1!
1%
#266830000000
0!
0%
#266835000000
1!
1%
#266840000000
0!
0%
#266845000000
1!
1%
#266850000000
0!
0%
#266855000000
1!
1%
#266860000000
0!
0%
#266865000000
1!
1%
#266870000000
0!
0%
#266875000000
1!
1%
#266880000000
0!
0%
#266885000000
1!
1%
#266890000000
0!
0%
#266895000000
1!
1%
#266900000000
0!
0%
#266905000000
1!
1%
#266910000000
0!
0%
#266915000000
1!
1%
#266920000000
0!
0%
#266925000000
1!
1%
#266930000000
0!
0%
#266935000000
1!
1%
#266940000000
0!
0%
#266945000000
1!
1%
#266950000000
0!
0%
#266955000000
1!
1%
#266960000000
0!
0%
#266965000000
1!
1%
#266970000000
0!
0%
#266975000000
1!
1%
#266980000000
0!
0%
#266985000000
1!
1%
#266990000000
0!
0%
#266995000000
1!
1%
#267000000000
0!
0%
#267005000000
1!
1%
#267010000000
0!
0%
#267015000000
1!
1%
#267020000000
0!
0%
#267025000000
1!
1%
#267030000000
0!
0%
#267035000000
1!
1%
#267040000000
0!
0%
#267045000000
1!
1%
#267050000000
0!
0%
#267055000000
1!
1%
#267060000000
0!
0%
#267065000000
1!
1%
#267070000000
0!
0%
#267075000000
1!
1%
#267080000000
0!
0%
#267085000000
1!
1%
#267090000000
0!
0%
#267095000000
1!
1%
#267100000000
0!
0%
#267105000000
1!
1%
#267110000000
0!
0%
#267115000000
1!
1%
#267120000000
0!
0%
#267125000000
1!
1%
#267130000000
0!
0%
#267135000000
1!
1%
#267140000000
0!
0%
#267145000000
1!
1%
#267150000000
0!
0%
#267155000000
1!
1%
#267160000000
0!
0%
#267165000000
1!
1%
#267170000000
0!
0%
#267175000000
1!
1%
#267180000000
0!
0%
#267185000000
1!
1%
#267190000000
0!
0%
#267195000000
1!
1%
#267200000000
0!
0%
#267205000000
1!
1%
#267210000000
0!
0%
#267215000000
1!
1%
#267220000000
0!
0%
#267225000000
1!
1%
#267230000000
0!
0%
#267235000000
1!
1%
#267240000000
0!
0%
#267245000000
1!
1%
#267250000000
0!
0%
#267255000000
1!
1%
#267260000000
0!
0%
#267265000000
1!
1%
#267270000000
0!
0%
#267275000000
1!
1%
#267280000000
0!
0%
#267285000000
1!
1%
#267290000000
0!
0%
#267295000000
1!
1%
#267300000000
0!
0%
#267305000000
1!
1%
#267310000000
0!
0%
#267315000000
1!
1%
#267320000000
0!
0%
#267325000000
1!
1%
#267330000000
0!
0%
#267335000000
1!
1%
#267340000000
0!
0%
#267345000000
1!
1%
#267350000000
0!
0%
#267355000000
1!
1%
#267360000000
0!
0%
#267365000000
1!
1%
#267370000000
0!
0%
#267375000000
1!
1%
#267380000000
0!
0%
#267385000000
1!
1%
#267390000000
0!
0%
#267395000000
1!
1%
#267400000000
0!
0%
#267405000000
1!
1%
#267410000000
0!
0%
#267415000000
1!
1%
#267420000000
0!
0%
#267425000000
1!
1%
#267430000000
0!
0%
#267435000000
1!
1%
#267440000000
0!
0%
#267445000000
1!
1%
#267450000000
0!
0%
#267455000000
1!
1%
#267460000000
0!
0%
#267465000000
1!
1%
#267470000000
0!
0%
#267475000000
1!
1%
#267480000000
0!
0%
#267485000000
1!
1%
#267490000000
0!
0%
#267495000000
1!
1%
#267500000000
0!
0%
#267505000000
1!
1%
#267510000000
0!
0%
#267515000000
1!
1%
#267520000000
0!
0%
#267525000000
1!
1%
#267530000000
0!
0%
#267535000000
1!
1%
#267540000000
0!
0%
#267545000000
1!
1%
#267550000000
0!
0%
#267555000000
1!
1%
#267560000000
0!
0%
#267565000000
1!
1%
#267570000000
0!
0%
#267575000000
1!
1%
#267580000000
0!
0%
#267585000000
1!
1%
#267590000000
0!
0%
#267595000000
1!
1%
#267600000000
0!
0%
#267605000000
1!
1%
#267610000000
0!
0%
#267615000000
1!
1%
#267620000000
0!
0%
#267625000000
1!
1%
#267630000000
0!
0%
#267635000000
1!
1%
#267640000000
0!
0%
#267645000000
1!
1%
#267650000000
0!
0%
#267655000000
1!
1%
#267660000000
0!
0%
#267665000000
1!
1%
#267670000000
0!
0%
#267675000000
1!
1%
#267680000000
0!
0%
#267685000000
1!
1%
#267690000000
0!
0%
#267695000000
1!
1%
#267700000000
0!
0%
#267705000000
1!
1%
#267710000000
0!
0%
#267715000000
1!
1%
#267720000000
0!
0%
#267725000000
1!
1%
#267730000000
0!
0%
#267735000000
1!
1%
#267740000000
0!
0%
#267745000000
1!
1%
#267750000000
0!
0%
#267755000000
1!
1%
#267760000000
0!
0%
#267765000000
1!
1%
#267770000000
0!
0%
#267775000000
1!
1%
#267780000000
0!
0%
#267785000000
1!
1%
#267790000000
0!
0%
#267795000000
1!
1%
#267800000000
0!
0%
#267805000000
1!
1%
#267810000000
0!
0%
#267815000000
1!
1%
#267820000000
0!
0%
#267825000000
1!
1%
#267830000000
0!
0%
#267835000000
1!
1%
#267840000000
0!
0%
#267845000000
1!
1%
#267850000000
0!
0%
#267855000000
1!
1%
#267860000000
0!
0%
#267865000000
1!
1%
#267870000000
0!
0%
#267875000000
1!
1%
#267880000000
0!
0%
#267885000000
1!
1%
#267890000000
0!
0%
#267895000000
1!
1%
#267900000000
0!
0%
#267905000000
1!
1%
#267910000000
0!
0%
#267915000000
1!
1%
#267920000000
0!
0%
#267925000000
1!
1%
#267930000000
0!
0%
#267935000000
1!
1%
#267940000000
0!
0%
#267945000000
1!
1%
#267950000000
0!
0%
#267955000000
1!
1%
#267960000000
0!
0%
#267965000000
1!
1%
#267970000000
0!
0%
#267975000000
1!
1%
#267980000000
0!
0%
#267985000000
1!
1%
#267990000000
0!
0%
#267995000000
1!
1%
#268000000000
0!
0%
#268005000000
1!
1%
#268010000000
0!
0%
#268015000000
1!
1%
#268020000000
0!
0%
#268025000000
1!
1%
#268030000000
0!
0%
#268035000000
1!
1%
#268040000000
0!
0%
#268045000000
1!
1%
#268050000000
0!
0%
#268055000000
1!
1%
#268060000000
0!
0%
#268065000000
1!
1%
#268070000000
0!
0%
#268075000000
1!
1%
#268080000000
0!
0%
#268085000000
1!
1%
#268090000000
0!
0%
#268095000000
1!
1%
#268100000000
0!
0%
#268105000000
1!
1%
#268110000000
0!
0%
#268115000000
1!
1%
#268120000000
0!
0%
#268125000000
1!
1%
#268130000000
0!
0%
#268135000000
1!
1%
#268140000000
0!
0%
#268145000000
1!
1%
#268150000000
0!
0%
#268155000000
1!
1%
#268160000000
0!
0%
#268165000000
1!
1%
#268170000000
0!
0%
#268175000000
1!
1%
#268180000000
0!
0%
#268185000000
1!
1%
#268190000000
0!
0%
#268195000000
1!
1%
#268200000000
0!
0%
#268205000000
1!
1%
#268210000000
0!
0%
#268215000000
1!
1%
#268220000000
0!
0%
#268225000000
1!
1%
#268230000000
0!
0%
#268235000000
1!
1%
#268240000000
0!
0%
#268245000000
1!
1%
#268250000000
0!
0%
#268255000000
1!
1%
#268260000000
0!
0%
#268265000000
1!
1%
#268270000000
0!
0%
#268275000000
1!
1%
#268280000000
0!
0%
#268285000000
1!
1%
#268290000000
0!
0%
#268295000000
1!
1%
#268300000000
0!
0%
#268305000000
1!
1%
#268310000000
0!
0%
#268315000000
1!
1%
#268320000000
0!
0%
#268325000000
1!
1%
#268330000000
0!
0%
#268335000000
1!
1%
#268340000000
0!
0%
#268345000000
1!
1%
#268350000000
0!
0%
#268355000000
1!
1%
#268360000000
0!
0%
#268365000000
1!
1%
#268370000000
0!
0%
#268375000000
1!
1%
#268380000000
0!
0%
#268385000000
1!
1%
#268390000000
0!
0%
#268395000000
1!
1%
#268400000000
0!
0%
#268405000000
1!
1%
#268410000000
0!
0%
#268415000000
1!
1%
#268420000000
0!
0%
#268425000000
1!
1%
#268430000000
0!
0%
#268435000000
1!
1%
#268440000000
0!
0%
#268445000000
1!
1%
#268450000000
0!
0%
#268455000000
1!
1%
#268460000000
0!
0%
#268465000000
1!
1%
#268470000000
0!
0%
#268475000000
1!
1%
#268480000000
0!
0%
#268485000000
1!
1%
#268490000000
0!
0%
#268495000000
1!
1%
#268500000000
0!
0%
#268505000000
1!
1%
#268510000000
0!
0%
#268515000000
1!
1%
#268520000000
0!
0%
#268525000000
1!
1%
#268530000000
0!
0%
#268535000000
1!
1%
#268540000000
0!
0%
#268545000000
1!
1%
#268550000000
0!
0%
#268555000000
1!
1%
#268560000000
0!
0%
#268565000000
1!
1%
#268570000000
0!
0%
#268575000000
1!
1%
#268580000000
0!
0%
#268585000000
1!
1%
#268590000000
0!
0%
#268595000000
1!
1%
#268600000000
0!
0%
#268605000000
1!
1%
#268610000000
0!
0%
#268615000000
1!
1%
#268620000000
0!
0%
#268625000000
1!
1%
#268630000000
0!
0%
#268635000000
1!
1%
#268640000000
0!
0%
#268645000000
1!
1%
#268650000000
0!
0%
#268655000000
1!
1%
#268660000000
0!
0%
#268665000000
1!
1%
#268670000000
0!
0%
#268675000000
1!
1%
#268680000000
0!
0%
#268685000000
1!
1%
#268690000000
0!
0%
#268695000000
1!
1%
#268700000000
0!
0%
#268705000000
1!
1%
#268710000000
0!
0%
#268715000000
1!
1%
#268720000000
0!
0%
#268725000000
1!
1%
#268730000000
0!
0%
#268735000000
1!
1%
#268740000000
0!
0%
#268745000000
1!
1%
#268750000000
0!
0%
#268755000000
1!
1%
#268760000000
0!
0%
#268765000000
1!
1%
#268770000000
0!
0%
#268775000000
1!
1%
#268780000000
0!
0%
#268785000000
1!
1%
#268790000000
0!
0%
#268795000000
1!
1%
#268800000000
0!
0%
#268805000000
1!
1%
#268810000000
0!
0%
#268815000000
1!
1%
#268820000000
0!
0%
#268825000000
1!
1%
#268830000000
0!
0%
#268835000000
1!
1%
#268840000000
0!
0%
#268845000000
1!
1%
#268850000000
0!
0%
#268855000000
1!
1%
#268860000000
0!
0%
#268865000000
1!
1%
#268870000000
0!
0%
#268875000000
1!
1%
#268880000000
0!
0%
#268885000000
1!
1%
#268890000000
0!
0%
#268895000000
1!
1%
#268900000000
0!
0%
#268905000000
1!
1%
#268910000000
0!
0%
#268915000000
1!
1%
#268920000000
0!
0%
#268925000000
1!
1%
#268930000000
0!
0%
#268935000000
1!
1%
#268940000000
0!
0%
#268945000000
1!
1%
#268950000000
0!
0%
#268955000000
1!
1%
#268960000000
0!
0%
#268965000000
1!
1%
#268970000000
0!
0%
#268975000000
1!
1%
#268980000000
0!
0%
#268985000000
1!
1%
#268990000000
0!
0%
#268995000000
1!
1%
#269000000000
0!
0%
#269005000000
1!
1%
#269010000000
0!
0%
#269015000000
1!
1%
#269020000000
0!
0%
#269025000000
1!
1%
#269030000000
0!
0%
#269035000000
1!
1%
#269040000000
0!
0%
#269045000000
1!
1%
#269050000000
0!
0%
#269055000000
1!
1%
#269060000000
0!
0%
#269065000000
1!
1%
#269070000000
0!
0%
#269075000000
1!
1%
#269080000000
0!
0%
#269085000000
1!
1%
#269090000000
0!
0%
#269095000000
1!
1%
#269100000000
0!
0%
#269105000000
1!
1%
#269110000000
0!
0%
#269115000000
1!
1%
#269120000000
0!
0%
#269125000000
1!
1%
#269130000000
0!
0%
#269135000000
1!
1%
#269140000000
0!
0%
#269145000000
1!
1%
#269150000000
0!
0%
#269155000000
1!
1%
#269160000000
0!
0%
#269165000000
1!
1%
#269170000000
0!
0%
#269175000000
1!
1%
#269180000000
0!
0%
#269185000000
1!
1%
#269190000000
0!
0%
#269195000000
1!
1%
#269200000000
0!
0%
#269205000000
1!
1%
#269210000000
0!
0%
#269215000000
1!
1%
#269220000000
0!
0%
#269225000000
1!
1%
#269230000000
0!
0%
#269235000000
1!
1%
#269240000000
0!
0%
#269245000000
1!
1%
#269250000000
0!
0%
#269255000000
1!
1%
#269260000000
0!
0%
#269265000000
1!
1%
#269270000000
0!
0%
#269275000000
1!
1%
#269280000000
0!
0%
#269285000000
1!
1%
#269290000000
0!
0%
#269295000000
1!
1%
#269300000000
0!
0%
#269305000000
1!
1%
#269310000000
0!
0%
#269315000000
1!
1%
#269320000000
0!
0%
#269325000000
1!
1%
#269330000000
0!
0%
#269335000000
1!
1%
#269340000000
0!
0%
#269345000000
1!
1%
#269350000000
0!
0%
#269355000000
1!
1%
#269360000000
0!
0%
#269365000000
1!
1%
#269370000000
0!
0%
#269375000000
1!
1%
#269380000000
0!
0%
#269385000000
1!
1%
#269390000000
0!
0%
#269395000000
1!
1%
#269400000000
0!
0%
#269405000000
1!
1%
#269410000000
0!
0%
#269415000000
1!
1%
#269420000000
0!
0%
#269425000000
1!
1%
#269430000000
0!
0%
#269435000000
1!
1%
#269440000000
0!
0%
#269445000000
1!
1%
#269450000000
0!
0%
#269455000000
1!
1%
#269460000000
0!
0%
#269465000000
1!
1%
#269470000000
0!
0%
#269475000000
1!
1%
#269480000000
0!
0%
#269485000000
1!
1%
#269490000000
0!
0%
#269495000000
1!
1%
#269500000000
0!
0%
#269505000000
1!
1%
#269510000000
0!
0%
#269515000000
1!
1%
#269520000000
0!
0%
#269525000000
1!
1%
#269530000000
0!
0%
#269535000000
1!
1%
#269540000000
0!
0%
#269545000000
1!
1%
#269550000000
0!
0%
#269555000000
1!
1%
#269560000000
0!
0%
#269565000000
1!
1%
#269570000000
0!
0%
#269575000000
1!
1%
#269580000000
0!
0%
#269585000000
1!
1%
#269590000000
0!
0%
#269595000000
1!
1%
#269600000000
0!
0%
#269605000000
1!
1%
#269610000000
0!
0%
#269615000000
1!
1%
#269620000000
0!
0%
#269625000000
1!
1%
#269630000000
0!
0%
#269635000000
1!
1%
#269640000000
0!
0%
#269645000000
1!
1%
#269650000000
0!
0%
#269655000000
1!
1%
#269660000000
0!
0%
#269665000000
1!
1%
#269670000000
0!
0%
#269675000000
1!
1%
#269680000000
0!
0%
#269685000000
1!
1%
#269690000000
0!
0%
#269695000000
1!
1%
#269700000000
0!
0%
#269705000000
1!
1%
#269710000000
0!
0%
#269715000000
1!
1%
#269720000000
0!
0%
#269725000000
1!
1%
#269730000000
0!
0%
#269735000000
1!
1%
#269740000000
0!
0%
#269745000000
1!
1%
#269750000000
0!
0%
#269755000000
1!
1%
#269760000000
0!
0%
#269765000000
1!
1%
#269770000000
0!
0%
#269775000000
1!
1%
#269780000000
0!
0%
#269785000000
1!
1%
#269790000000
0!
0%
#269795000000
1!
1%
#269800000000
0!
0%
#269805000000
1!
1%
#269810000000
0!
0%
#269815000000
1!
1%
#269820000000
0!
0%
#269825000000
1!
1%
#269830000000
0!
0%
#269835000000
1!
1%
#269840000000
0!
0%
#269845000000
1!
1%
#269850000000
0!
0%
#269855000000
1!
1%
#269860000000
0!
0%
#269865000000
1!
1%
#269870000000
0!
0%
#269875000000
1!
1%
#269880000000
0!
0%
#269885000000
1!
1%
#269890000000
0!
0%
#269895000000
1!
1%
#269900000000
0!
0%
#269905000000
1!
1%
#269910000000
0!
0%
#269915000000
1!
1%
#269920000000
0!
0%
#269925000000
1!
1%
#269930000000
0!
0%
#269935000000
1!
1%
#269940000000
0!
0%
#269945000000
1!
1%
#269950000000
0!
0%
#269955000000
1!
1%
#269960000000
0!
0%
#269965000000
1!
1%
#269970000000
0!
0%
#269975000000
1!
1%
#269980000000
0!
0%
#269985000000
1!
1%
#269990000000
0!
0%
#269995000000
1!
1%
#270000000000
0!
0%
#270005000000
1!
1%
#270010000000
0!
0%
#270015000000
1!
1%
#270020000000
0!
0%
#270025000000
1!
1%
#270030000000
0!
0%
#270035000000
1!
1%
#270040000000
0!
0%
#270045000000
1!
1%
#270050000000
0!
0%
#270055000000
1!
1%
#270060000000
0!
0%
#270065000000
1!
1%
#270070000000
0!
0%
#270075000000
1!
1%
#270080000000
0!
0%
#270085000000
1!
1%
#270090000000
0!
0%
#270095000000
1!
1%
#270100000000
0!
0%
#270105000000
1!
1%
#270110000000
0!
0%
#270115000000
1!
1%
#270120000000
0!
0%
#270125000000
1!
1%
#270130000000
0!
0%
#270135000000
1!
1%
#270140000000
0!
0%
#270145000000
1!
1%
#270150000000
0!
0%
#270155000000
1!
1%
#270160000000
0!
0%
#270165000000
1!
1%
#270170000000
0!
0%
#270175000000
1!
1%
#270180000000
0!
0%
#270185000000
1!
1%
#270190000000
0!
0%
#270195000000
1!
1%
#270200000000
0!
0%
#270205000000
1!
1%
#270210000000
0!
0%
#270215000000
1!
1%
#270220000000
0!
0%
#270225000000
1!
1%
#270230000000
0!
0%
#270235000000
1!
1%
#270240000000
0!
0%
#270245000000
1!
1%
#270250000000
0!
0%
#270255000000
1!
1%
#270260000000
0!
0%
#270265000000
1!
1%
#270270000000
0!
0%
#270275000000
1!
1%
#270280000000
0!
0%
#270285000000
1!
1%
#270290000000
0!
0%
#270295000000
1!
1%
#270300000000
0!
0%
#270305000000
1!
1%
#270310000000
0!
0%
#270315000000
1!
1%
#270320000000
0!
0%
#270325000000
1!
1%
#270330000000
0!
0%
#270335000000
1!
1%
#270340000000
0!
0%
#270345000000
1!
1%
#270350000000
0!
0%
#270355000000
1!
1%
#270360000000
0!
0%
#270365000000
1!
1%
#270370000000
0!
0%
#270375000000
1!
1%
#270380000000
0!
0%
#270385000000
1!
1%
#270390000000
0!
0%
#270395000000
1!
1%
#270400000000
0!
0%
#270405000000
1!
1%
#270410000000
0!
0%
#270415000000
1!
1%
#270420000000
0!
0%
#270425000000
1!
1%
#270430000000
0!
0%
#270435000000
1!
1%
#270440000000
0!
0%
#270445000000
1!
1%
#270450000000
0!
0%
#270455000000
1!
1%
#270460000000
0!
0%
#270465000000
1!
1%
#270470000000
0!
0%
#270475000000
1!
1%
#270480000000
0!
0%
#270485000000
1!
1%
#270490000000
0!
0%
#270495000000
1!
1%
#270500000000
0!
0%
#270505000000
1!
1%
#270510000000
0!
0%
#270515000000
1!
1%
#270520000000
0!
0%
#270525000000
1!
1%
#270530000000
0!
0%
#270535000000
1!
1%
#270540000000
0!
0%
#270545000000
1!
1%
#270550000000
0!
0%
#270555000000
1!
1%
#270560000000
0!
0%
#270565000000
1!
1%
#270570000000
0!
0%
#270575000000
1!
1%
#270580000000
0!
0%
#270585000000
1!
1%
#270590000000
0!
0%
#270595000000
1!
1%
#270600000000
0!
0%
#270605000000
1!
1%
#270610000000
0!
0%
#270615000000
1!
1%
#270620000000
0!
0%
#270625000000
1!
1%
#270630000000
0!
0%
#270635000000
1!
1%
#270640000000
0!
0%
#270645000000
1!
1%
#270650000000
0!
0%
#270655000000
1!
1%
#270660000000
0!
0%
#270665000000
1!
1%
#270670000000
0!
0%
#270675000000
1!
1%
#270680000000
0!
0%
#270685000000
1!
1%
#270690000000
0!
0%
#270695000000
1!
1%
#270700000000
0!
0%
#270705000000
1!
1%
#270710000000
0!
0%
#270715000000
1!
1%
#270720000000
0!
0%
#270725000000
1!
1%
#270730000000
0!
0%
#270735000000
1!
1%
#270740000000
0!
0%
#270745000000
1!
1%
#270750000000
0!
0%
#270755000000
1!
1%
#270760000000
0!
0%
#270765000000
1!
1%
#270770000000
0!
0%
#270775000000
1!
1%
#270780000000
0!
0%
#270785000000
1!
1%
#270790000000
0!
0%
#270795000000
1!
1%
#270800000000
0!
0%
#270805000000
1!
1%
#270810000000
0!
0%
#270815000000
1!
1%
#270820000000
0!
0%
#270825000000
1!
1%
#270830000000
0!
0%
#270835000000
1!
1%
#270840000000
0!
0%
#270845000000
1!
1%
#270850000000
0!
0%
#270855000000
1!
1%
#270860000000
0!
0%
#270865000000
1!
1%
#270870000000
0!
0%
#270875000000
1!
1%
#270880000000
0!
0%
#270885000000
1!
1%
#270890000000
0!
0%
#270895000000
1!
1%
#270900000000
0!
0%
#270905000000
1!
1%
#270910000000
0!
0%
#270915000000
1!
1%
#270920000000
0!
0%
#270925000000
1!
1%
#270930000000
0!
0%
#270935000000
1!
1%
#270940000000
0!
0%
#270945000000
1!
1%
#270950000000
0!
0%
#270955000000
1!
1%
#270960000000
0!
0%
#270965000000
1!
1%
#270970000000
0!
0%
#270975000000
1!
1%
#270980000000
0!
0%
#270985000000
1!
1%
#270990000000
0!
0%
#270995000000
1!
1%
#271000000000
0!
0%
#271005000000
1!
1%
#271010000000
0!
0%
#271015000000
1!
1%
#271020000000
0!
0%
#271025000000
1!
1%
#271030000000
0!
0%
#271035000000
1!
1%
#271040000000
0!
0%
#271045000000
1!
1%
#271050000000
0!
0%
#271055000000
1!
1%
#271060000000
0!
0%
#271065000000
1!
1%
#271070000000
0!
0%
#271075000000
1!
1%
#271080000000
0!
0%
#271085000000
1!
1%
#271090000000
0!
0%
#271095000000
1!
1%
#271100000000
0!
0%
#271105000000
1!
1%
#271110000000
0!
0%
#271115000000
1!
1%
#271120000000
0!
0%
#271125000000
1!
1%
#271130000000
0!
0%
#271135000000
1!
1%
#271140000000
0!
0%
#271145000000
1!
1%
#271150000000
0!
0%
#271155000000
1!
1%
#271160000000
0!
0%
#271165000000
1!
1%
#271170000000
0!
0%
#271175000000
1!
1%
#271180000000
0!
0%
#271185000000
1!
1%
#271190000000
0!
0%
#271195000000
1!
1%
#271200000000
0!
0%
#271205000000
1!
1%
#271210000000
0!
0%
#271215000000
1!
1%
#271220000000
0!
0%
#271225000000
1!
1%
#271230000000
0!
0%
#271235000000
1!
1%
#271240000000
0!
0%
#271245000000
1!
1%
#271250000000
0!
0%
#271255000000
1!
1%
#271260000000
0!
0%
#271265000000
1!
1%
#271270000000
0!
0%
#271275000000
1!
1%
#271280000000
0!
0%
#271285000000
1!
1%
#271290000000
0!
0%
#271295000000
1!
1%
#271300000000
0!
0%
#271305000000
1!
1%
#271310000000
0!
0%
#271315000000
1!
1%
#271320000000
0!
0%
#271325000000
1!
1%
#271330000000
0!
0%
#271335000000
1!
1%
#271340000000
0!
0%
#271345000000
1!
1%
#271350000000
0!
0%
#271355000000
1!
1%
#271360000000
0!
0%
#271365000000
1!
1%
#271370000000
0!
0%
#271375000000
1!
1%
#271380000000
0!
0%
#271385000000
1!
1%
#271390000000
0!
0%
#271395000000
1!
1%
#271400000000
0!
0%
#271405000000
1!
1%
#271410000000
0!
0%
#271415000000
1!
1%
#271420000000
0!
0%
#271425000000
1!
1%
#271430000000
0!
0%
#271435000000
1!
1%
#271440000000
0!
0%
#271445000000
1!
1%
#271450000000
0!
0%
#271455000000
1!
1%
#271460000000
0!
0%
#271465000000
1!
1%
#271470000000
0!
0%
#271475000000
1!
1%
#271480000000
0!
0%
#271485000000
1!
1%
#271490000000
0!
0%
#271495000000
1!
1%
#271500000000
0!
0%
#271505000000
1!
1%
#271510000000
0!
0%
#271515000000
1!
1%
#271520000000
0!
0%
#271525000000
1!
1%
#271530000000
0!
0%
#271535000000
1!
1%
#271540000000
0!
0%
#271545000000
1!
1%
#271550000000
0!
0%
#271555000000
1!
1%
#271560000000
0!
0%
#271565000000
1!
1%
#271570000000
0!
0%
#271575000000
1!
1%
#271580000000
0!
0%
#271585000000
1!
1%
#271590000000
0!
0%
#271595000000
1!
1%
#271600000000
0!
0%
#271605000000
1!
1%
#271610000000
0!
0%
#271615000000
1!
1%
#271620000000
0!
0%
#271625000000
1!
1%
#271630000000
0!
0%
#271635000000
1!
1%
#271640000000
0!
0%
#271645000000
1!
1%
#271650000000
0!
0%
#271655000000
1!
1%
#271660000000
0!
0%
#271665000000
1!
1%
#271670000000
0!
0%
#271675000000
1!
1%
#271680000000
0!
0%
#271685000000
1!
1%
#271690000000
0!
0%
#271695000000
1!
1%
#271700000000
0!
0%
#271705000000
1!
1%
#271710000000
0!
0%
#271715000000
1!
1%
#271720000000
0!
0%
#271725000000
1!
1%
#271730000000
0!
0%
#271735000000
1!
1%
#271740000000
0!
0%
#271745000000
1!
1%
#271750000000
0!
0%
#271755000000
1!
1%
#271760000000
0!
0%
#271765000000
1!
1%
#271770000000
0!
0%
#271775000000
1!
1%
#271780000000
0!
0%
#271785000000
1!
1%
#271790000000
0!
0%
#271795000000
1!
1%
#271800000000
0!
0%
#271805000000
1!
1%
#271810000000
0!
0%
#271815000000
1!
1%
#271820000000
0!
0%
#271825000000
1!
1%
#271830000000
0!
0%
#271835000000
1!
1%
#271840000000
0!
0%
#271845000000
1!
1%
#271850000000
0!
0%
#271855000000
1!
1%
#271860000000
0!
0%
#271865000000
1!
1%
#271870000000
0!
0%
#271875000000
1!
1%
#271880000000
0!
0%
#271885000000
1!
1%
#271890000000
0!
0%
#271895000000
1!
1%
#271900000000
0!
0%
#271905000000
1!
1%
#271910000000
0!
0%
#271915000000
1!
1%
#271920000000
0!
0%
#271925000000
1!
1%
#271930000000
0!
0%
#271935000000
1!
1%
#271940000000
0!
0%
#271945000000
1!
1%
#271950000000
0!
0%
#271955000000
1!
1%
#271960000000
0!
0%
#271965000000
1!
1%
#271970000000
0!
0%
#271975000000
1!
1%
#271980000000
0!
0%
#271985000000
1!
1%
#271990000000
0!
0%
#271995000000
1!
1%
#272000000000
0!
0%
#272005000000
1!
1%
#272010000000
0!
0%
#272015000000
1!
1%
#272020000000
0!
0%
#272025000000
1!
1%
#272030000000
0!
0%
#272035000000
1!
1%
#272040000000
0!
0%
#272045000000
1!
1%
#272050000000
0!
0%
#272055000000
1!
1%
#272060000000
0!
0%
#272065000000
1!
1%
#272070000000
0!
0%
#272075000000
1!
1%
#272080000000
0!
0%
#272085000000
1!
1%
#272090000000
0!
0%
#272095000000
1!
1%
#272100000000
0!
0%
#272105000000
1!
1%
#272110000000
0!
0%
#272115000000
1!
1%
#272120000000
0!
0%
#272125000000
1!
1%
#272130000000
0!
0%
#272135000000
1!
1%
#272140000000
0!
0%
#272145000000
1!
1%
#272150000000
0!
0%
#272155000000
1!
1%
#272160000000
0!
0%
#272165000000
1!
1%
#272170000000
0!
0%
#272175000000
1!
1%
#272180000000
0!
0%
#272185000000
1!
1%
#272190000000
0!
0%
#272195000000
1!
1%
#272200000000
0!
0%
#272205000000
1!
1%
#272210000000
0!
0%
#272215000000
1!
1%
#272220000000
0!
0%
#272225000000
1!
1%
#272230000000
0!
0%
#272235000000
1!
1%
#272240000000
0!
0%
#272245000000
1!
1%
#272250000000
0!
0%
#272255000000
1!
1%
#272260000000
0!
0%
#272265000000
1!
1%
#272270000000
0!
0%
#272275000000
1!
1%
#272280000000
0!
0%
#272285000000
1!
1%
#272290000000
0!
0%
#272295000000
1!
1%
#272300000000
0!
0%
#272305000000
1!
1%
#272310000000
0!
0%
#272315000000
1!
1%
#272320000000
0!
0%
#272325000000
1!
1%
#272330000000
0!
0%
#272335000000
1!
1%
#272340000000
0!
0%
#272345000000
1!
1%
#272350000000
0!
0%
#272355000000
1!
1%
#272360000000
0!
0%
#272365000000
1!
1%
#272370000000
0!
0%
#272375000000
1!
1%
#272380000000
0!
0%
#272385000000
1!
1%
#272390000000
0!
0%
#272395000000
1!
1%
#272400000000
0!
0%
#272405000000
1!
1%
#272410000000
0!
0%
#272415000000
1!
1%
#272420000000
0!
0%
#272425000000
1!
1%
#272430000000
0!
0%
#272435000000
1!
1%
#272440000000
0!
0%
#272445000000
1!
1%
#272450000000
0!
0%
#272455000000
1!
1%
#272460000000
0!
0%
#272465000000
1!
1%
#272470000000
0!
0%
#272475000000
1!
1%
#272480000000
0!
0%
#272485000000
1!
1%
#272490000000
0!
0%
#272495000000
1!
1%
#272500000000
0!
0%
#272505000000
1!
1%
#272510000000
0!
0%
#272515000000
1!
1%
#272520000000
0!
0%
#272525000000
1!
1%
#272530000000
0!
0%
#272535000000
1!
1%
#272540000000
0!
0%
#272545000000
1!
1%
#272550000000
0!
0%
#272555000000
1!
1%
#272560000000
0!
0%
#272565000000
1!
1%
#272570000000
0!
0%
#272575000000
1!
1%
#272580000000
0!
0%
#272585000000
1!
1%
#272590000000
0!
0%
#272595000000
1!
1%
#272600000000
0!
0%
#272605000000
1!
1%
#272610000000
0!
0%
#272615000000
1!
1%
#272620000000
0!
0%
#272625000000
1!
1%
#272630000000
0!
0%
#272635000000
1!
1%
#272640000000
0!
0%
#272645000000
1!
1%
#272650000000
0!
0%
#272655000000
1!
1%
#272660000000
0!
0%
#272665000000
1!
1%
#272670000000
0!
0%
#272675000000
1!
1%
#272680000000
0!
0%
#272685000000
1!
1%
#272690000000
0!
0%
#272695000000
1!
1%
#272700000000
0!
0%
#272705000000
1!
1%
#272710000000
0!
0%
#272715000000
1!
1%
#272720000000
0!
0%
#272725000000
1!
1%
#272730000000
0!
0%
#272735000000
1!
1%
#272740000000
0!
0%
#272745000000
1!
1%
#272750000000
0!
0%
#272755000000
1!
1%
#272760000000
0!
0%
#272765000000
1!
1%
#272770000000
0!
0%
#272775000000
1!
1%
#272780000000
0!
0%
#272785000000
1!
1%
#272790000000
0!
0%
#272795000000
1!
1%
#272800000000
0!
0%
#272805000000
1!
1%
#272810000000
0!
0%
#272815000000
1!
1%
#272820000000
0!
0%
#272825000000
1!
1%
#272830000000
0!
0%
#272835000000
1!
1%
#272840000000
0!
0%
#272845000000
1!
1%
#272850000000
0!
0%
#272855000000
1!
1%
#272860000000
0!
0%
#272865000000
1!
1%
#272870000000
0!
0%
#272875000000
1!
1%
#272880000000
0!
0%
#272885000000
1!
1%
#272890000000
0!
0%
#272895000000
1!
1%
#272900000000
0!
0%
#272905000000
1!
1%
#272910000000
0!
0%
#272915000000
1!
1%
#272920000000
0!
0%
#272925000000
1!
1%
#272930000000
0!
0%
#272935000000
1!
1%
#272940000000
0!
0%
#272945000000
1!
1%
#272950000000
0!
0%
#272955000000
1!
1%
#272960000000
0!
0%
#272965000000
1!
1%
#272970000000
0!
0%
#272975000000
1!
1%
#272980000000
0!
0%
#272985000000
1!
1%
#272990000000
0!
0%
#272995000000
1!
1%
#273000000000
0!
0%
#273005000000
1!
1%
#273010000000
0!
0%
#273015000000
1!
1%
#273020000000
0!
0%
#273025000000
1!
1%
#273030000000
0!
0%
#273035000000
1!
1%
#273040000000
0!
0%
#273045000000
1!
1%
#273050000000
0!
0%
#273055000000
1!
1%
#273060000000
0!
0%
#273065000000
1!
1%
#273070000000
0!
0%
#273075000000
1!
1%
#273080000000
0!
0%
#273085000000
1!
1%
#273090000000
0!
0%
#273095000000
1!
1%
#273100000000
0!
0%
#273105000000
1!
1%
#273110000000
0!
0%
#273115000000
1!
1%
#273120000000
0!
0%
#273125000000
1!
1%
#273130000000
0!
0%
#273135000000
1!
1%
#273140000000
0!
0%
#273145000000
1!
1%
#273150000000
0!
0%
#273155000000
1!
1%
#273160000000
0!
0%
#273165000000
1!
1%
#273170000000
0!
0%
#273175000000
1!
1%
#273180000000
0!
0%
#273185000000
1!
1%
#273190000000
0!
0%
#273195000000
1!
1%
#273200000000
0!
0%
#273205000000
1!
1%
#273210000000
0!
0%
#273215000000
1!
1%
#273220000000
0!
0%
#273225000000
1!
1%
#273230000000
0!
0%
#273235000000
1!
1%
#273240000000
0!
0%
#273245000000
1!
1%
#273250000000
0!
0%
#273255000000
1!
1%
#273260000000
0!
0%
#273265000000
1!
1%
#273270000000
0!
0%
#273275000000
1!
1%
#273280000000
0!
0%
#273285000000
1!
1%
#273290000000
0!
0%
#273295000000
1!
1%
#273300000000
0!
0%
#273305000000
1!
1%
#273310000000
0!
0%
#273315000000
1!
1%
#273320000000
0!
0%
#273325000000
1!
1%
#273330000000
0!
0%
#273335000000
1!
1%
#273340000000
0!
0%
#273345000000
1!
1%
#273350000000
0!
0%
#273355000000
1!
1%
#273360000000
0!
0%
#273365000000
1!
1%
#273370000000
0!
0%
#273375000000
1!
1%
#273380000000
0!
0%
#273385000000
1!
1%
#273390000000
0!
0%
#273395000000
1!
1%
#273400000000
0!
0%
#273405000000
1!
1%
#273410000000
0!
0%
#273415000000
1!
1%
#273420000000
0!
0%
#273425000000
1!
1%
#273430000000
0!
0%
#273435000000
1!
1%
#273440000000
0!
0%
#273445000000
1!
1%
#273450000000
0!
0%
#273455000000
1!
1%
#273460000000
0!
0%
#273465000000
1!
1%
#273470000000
0!
0%
#273475000000
1!
1%
#273480000000
0!
0%
#273485000000
1!
1%
#273490000000
0!
0%
#273495000000
1!
1%
#273500000000
0!
0%
#273505000000
1!
1%
#273510000000
0!
0%
#273515000000
1!
1%
#273520000000
0!
0%
#273525000000
1!
1%
#273530000000
0!
0%
#273535000000
1!
1%
#273540000000
0!
0%
#273545000000
1!
1%
#273550000000
0!
0%
#273555000000
1!
1%
#273560000000
0!
0%
#273565000000
1!
1%
#273570000000
0!
0%
#273575000000
1!
1%
#273580000000
0!
0%
#273585000000
1!
1%
#273590000000
0!
0%
#273595000000
1!
1%
#273600000000
0!
0%
#273605000000
1!
1%
#273610000000
0!
0%
#273615000000
1!
1%
#273620000000
0!
0%
#273625000000
1!
1%
#273630000000
0!
0%
#273635000000
1!
1%
#273640000000
0!
0%
#273645000000
1!
1%
#273650000000
0!
0%
#273655000000
1!
1%
#273660000000
0!
0%
#273665000000
1!
1%
#273670000000
0!
0%
#273675000000
1!
1%
#273680000000
0!
0%
#273685000000
1!
1%
#273690000000
0!
0%
#273695000000
1!
1%
#273700000000
0!
0%
#273705000000
1!
1%
#273710000000
0!
0%
#273715000000
1!
1%
#273720000000
0!
0%
#273725000000
1!
1%
#273730000000
0!
0%
#273735000000
1!
1%
#273740000000
0!
0%
#273745000000
1!
1%
#273750000000
0!
0%
#273755000000
1!
1%
#273760000000
0!
0%
#273765000000
1!
1%
#273770000000
0!
0%
#273775000000
1!
1%
#273780000000
0!
0%
#273785000000
1!
1%
#273790000000
0!
0%
#273795000000
1!
1%
#273800000000
0!
0%
#273805000000
1!
1%
#273810000000
0!
0%
#273815000000
1!
1%
#273820000000
0!
0%
#273825000000
1!
1%
#273830000000
0!
0%
#273835000000
1!
1%
#273840000000
0!
0%
#273845000000
1!
1%
#273850000000
0!
0%
#273855000000
1!
1%
#273860000000
0!
0%
#273865000000
1!
1%
#273870000000
0!
0%
#273875000000
1!
1%
#273880000000
0!
0%
#273885000000
1!
1%
#273890000000
0!
0%
#273895000000
1!
1%
#273900000000
0!
0%
#273905000000
1!
1%
#273910000000
0!
0%
#273915000000
1!
1%
#273920000000
0!
0%
#273925000000
1!
1%
#273930000000
0!
0%
#273935000000
1!
1%
#273940000000
0!
0%
#273945000000
1!
1%
#273950000000
0!
0%
#273955000000
1!
1%
#273960000000
0!
0%
#273965000000
1!
1%
#273970000000
0!
0%
#273975000000
1!
1%
#273980000000
0!
0%
#273985000000
1!
1%
#273990000000
0!
0%
#273995000000
1!
1%
#274000000000
0!
0%
#274005000000
1!
1%
#274010000000
0!
0%
#274015000000
1!
1%
#274020000000
0!
0%
#274025000000
1!
1%
#274030000000
0!
0%
#274035000000
1!
1%
#274040000000
0!
0%
#274045000000
1!
1%
#274050000000
0!
0%
#274055000000
1!
1%
#274060000000
0!
0%
#274065000000
1!
1%
#274070000000
0!
0%
#274075000000
1!
1%
#274080000000
0!
0%
#274085000000
1!
1%
#274090000000
0!
0%
#274095000000
1!
1%
#274100000000
0!
0%
#274105000000
1!
1%
#274110000000
0!
0%
#274115000000
1!
1%
#274120000000
0!
0%
#274125000000
1!
1%
#274130000000
0!
0%
#274135000000
1!
1%
#274140000000
0!
0%
#274145000000
1!
1%
#274150000000
0!
0%
#274155000000
1!
1%
#274160000000
0!
0%
#274165000000
1!
1%
#274170000000
0!
0%
#274175000000
1!
1%
#274180000000
0!
0%
#274185000000
1!
1%
#274190000000
0!
0%
#274195000000
1!
1%
#274200000000
0!
0%
#274205000000
1!
1%
#274210000000
0!
0%
#274215000000
1!
1%
#274220000000
0!
0%
#274225000000
1!
1%
#274230000000
0!
0%
#274235000000
1!
1%
#274240000000
0!
0%
#274245000000
1!
1%
#274250000000
0!
0%
#274255000000
1!
1%
#274260000000
0!
0%
#274265000000
1!
1%
#274270000000
0!
0%
#274275000000
1!
1%
#274280000000
0!
0%
#274285000000
1!
1%
#274290000000
0!
0%
#274295000000
1!
1%
#274300000000
0!
0%
#274305000000
1!
1%
#274310000000
0!
0%
#274315000000
1!
1%
#274320000000
0!
0%
#274325000000
1!
1%
#274330000000
0!
0%
#274335000000
1!
1%
#274340000000
0!
0%
#274345000000
1!
1%
#274350000000
0!
0%
#274355000000
1!
1%
#274360000000
0!
0%
#274365000000
1!
1%
#274370000000
0!
0%
#274375000000
1!
1%
#274380000000
0!
0%
#274385000000
1!
1%
#274390000000
0!
0%
#274395000000
1!
1%
#274400000000
0!
0%
#274405000000
1!
1%
#274410000000
0!
0%
#274415000000
1!
1%
#274420000000
0!
0%
#274425000000
1!
1%
#274430000000
0!
0%
#274435000000
1!
1%
#274440000000
0!
0%
#274445000000
1!
1%
#274450000000
0!
0%
#274455000000
1!
1%
#274460000000
0!
0%
#274465000000
1!
1%
#274470000000
0!
0%
#274475000000
1!
1%
#274480000000
0!
0%
#274485000000
1!
1%
#274490000000
0!
0%
#274495000000
1!
1%
#274500000000
0!
0%
#274505000000
1!
1%
#274510000000
0!
0%
#274515000000
1!
1%
#274520000000
0!
0%
#274525000000
1!
1%
#274530000000
0!
0%
#274535000000
1!
1%
#274540000000
0!
0%
#274545000000
1!
1%
#274550000000
0!
0%
#274555000000
1!
1%
#274560000000
0!
0%
#274565000000
1!
1%
#274570000000
0!
0%
#274575000000
1!
1%
#274580000000
0!
0%
#274585000000
1!
1%
#274590000000
0!
0%
#274595000000
1!
1%
#274600000000
0!
0%
#274605000000
1!
1%
#274610000000
0!
0%
#274615000000
1!
1%
#274620000000
0!
0%
#274625000000
1!
1%
#274630000000
0!
0%
#274635000000
1!
1%
#274640000000
0!
0%
#274645000000
1!
1%
#274650000000
0!
0%
#274655000000
1!
1%
#274660000000
0!
0%
#274665000000
1!
1%
#274670000000
0!
0%
#274675000000
1!
1%
#274680000000
0!
0%
#274685000000
1!
1%
#274690000000
0!
0%
#274695000000
1!
1%
#274700000000
0!
0%
#274705000000
1!
1%
#274710000000
0!
0%
#274715000000
1!
1%
#274720000000
0!
0%
#274725000000
1!
1%
#274730000000
0!
0%
#274735000000
1!
1%
#274740000000
0!
0%
#274745000000
1!
1%
#274750000000
0!
0%
#274755000000
1!
1%
#274760000000
0!
0%
#274765000000
1!
1%
#274770000000
0!
0%
#274775000000
1!
1%
#274780000000
0!
0%
#274785000000
1!
1%
#274790000000
0!
0%
#274795000000
1!
1%
#274800000000
0!
0%
#274805000000
1!
1%
#274810000000
0!
0%
#274815000000
1!
1%
#274820000000
0!
0%
#274825000000
1!
1%
#274830000000
0!
0%
#274835000000
1!
1%
#274840000000
0!
0%
#274845000000
1!
1%
#274850000000
0!
0%
#274855000000
1!
1%
#274860000000
0!
0%
#274865000000
1!
1%
#274870000000
0!
0%
#274875000000
1!
1%
#274880000000
0!
0%
#274885000000
1!
1%
#274890000000
0!
0%
#274895000000
1!
1%
#274900000000
0!
0%
#274905000000
1!
1%
#274910000000
0!
0%
#274915000000
1!
1%
#274920000000
0!
0%
#274925000000
1!
1%
#274930000000
0!
0%
#274935000000
1!
1%
#274940000000
0!
0%
#274945000000
1!
1%
#274950000000
0!
0%
#274955000000
1!
1%
#274960000000
0!
0%
#274965000000
1!
1%
#274970000000
0!
0%
#274975000000
1!
1%
#274980000000
0!
0%
#274985000000
1!
1%
#274990000000
0!
0%
#274995000000
1!
1%
#275000000000
0!
0%
#275005000000
1!
1%
#275010000000
0!
0%
#275015000000
1!
1%
#275020000000
0!
0%
#275025000000
1!
1%
#275030000000
0!
0%
#275035000000
1!
1%
#275040000000
0!
0%
#275045000000
1!
1%
#275050000000
0!
0%
#275055000000
1!
1%
#275060000000
0!
0%
#275065000000
1!
1%
#275070000000
0!
0%
#275075000000
1!
1%
#275080000000
0!
0%
#275085000000
1!
1%
#275090000000
0!
0%
#275095000000
1!
1%
#275100000000
0!
0%
#275105000000
1!
1%
#275110000000
0!
0%
#275115000000
1!
1%
#275120000000
0!
0%
#275125000000
1!
1%
#275130000000
0!
0%
#275135000000
1!
1%
#275140000000
0!
0%
#275145000000
1!
1%
#275150000000
0!
0%
#275155000000
1!
1%
#275160000000
0!
0%
#275165000000
1!
1%
#275170000000
0!
0%
#275175000000
1!
1%
#275180000000
0!
0%
#275185000000
1!
1%
#275190000000
0!
0%
#275195000000
1!
1%
#275200000000
0!
0%
#275205000000
1!
1%
#275210000000
0!
0%
#275215000000
1!
1%
#275220000000
0!
0%
#275225000000
1!
1%
#275230000000
0!
0%
#275235000000
1!
1%
#275240000000
0!
0%
#275245000000
1!
1%
#275250000000
0!
0%
#275255000000
1!
1%
#275260000000
0!
0%
#275265000000
1!
1%
#275270000000
0!
0%
#275275000000
1!
1%
#275280000000
0!
0%
#275285000000
1!
1%
#275290000000
0!
0%
#275295000000
1!
1%
#275300000000
0!
0%
#275305000000
1!
1%
#275310000000
0!
0%
#275315000000
1!
1%
#275320000000
0!
0%
#275325000000
1!
1%
#275330000000
0!
0%
#275335000000
1!
1%
#275340000000
0!
0%
#275345000000
1!
1%
#275350000000
0!
0%
#275355000000
1!
1%
#275360000000
0!
0%
#275365000000
1!
1%
#275370000000
0!
0%
#275375000000
1!
1%
#275380000000
0!
0%
#275385000000
1!
1%
#275390000000
0!
0%
#275395000000
1!
1%
#275400000000
0!
0%
#275405000000
1!
1%
#275410000000
0!
0%
#275415000000
1!
1%
#275420000000
0!
0%
#275425000000
1!
1%
#275430000000
0!
0%
#275435000000
1!
1%
#275440000000
0!
0%
#275445000000
1!
1%
#275450000000
0!
0%
#275455000000
1!
1%
#275460000000
0!
0%
#275465000000
1!
1%
#275470000000
0!
0%
#275475000000
1!
1%
#275480000000
0!
0%
#275485000000
1!
1%
#275490000000
0!
0%
#275495000000
1!
1%
#275500000000
0!
0%
#275505000000
1!
1%
#275510000000
0!
0%
#275515000000
1!
1%
#275520000000
0!
0%
#275525000000
1!
1%
#275530000000
0!
0%
#275535000000
1!
1%
#275540000000
0!
0%
#275545000000
1!
1%
#275550000000
0!
0%
#275555000000
1!
1%
#275560000000
0!
0%
#275565000000
1!
1%
#275570000000
0!
0%
#275575000000
1!
1%
#275580000000
0!
0%
#275585000000
1!
1%
#275590000000
0!
0%
#275595000000
1!
1%
#275600000000
0!
0%
#275605000000
1!
1%
#275610000000
0!
0%
#275615000000
1!
1%
#275620000000
0!
0%
#275625000000
1!
1%
#275630000000
0!
0%
#275635000000
1!
1%
#275640000000
0!
0%
#275645000000
1!
1%
#275650000000
0!
0%
#275655000000
1!
1%
#275660000000
0!
0%
#275665000000
1!
1%
#275670000000
0!
0%
#275675000000
1!
1%
#275680000000
0!
0%
#275685000000
1!
1%
#275690000000
0!
0%
#275695000000
1!
1%
#275700000000
0!
0%
#275705000000
1!
1%
#275710000000
0!
0%
#275715000000
1!
1%
#275720000000
0!
0%
#275725000000
1!
1%
#275730000000
0!
0%
#275735000000
1!
1%
#275740000000
0!
0%
#275745000000
1!
1%
#275750000000
0!
0%
#275755000000
1!
1%
#275760000000
0!
0%
#275765000000
1!
1%
#275770000000
0!
0%
#275775000000
1!
1%
#275780000000
0!
0%
#275785000000
1!
1%
#275790000000
0!
0%
#275795000000
1!
1%
#275800000000
0!
0%
#275805000000
1!
1%
#275810000000
0!
0%
#275815000000
1!
1%
#275820000000
0!
0%
#275825000000
1!
1%
#275830000000
0!
0%
#275835000000
1!
1%
#275840000000
0!
0%
#275845000000
1!
1%
#275850000000
0!
0%
#275855000000
1!
1%
#275860000000
0!
0%
#275865000000
1!
1%
#275870000000
0!
0%
#275875000000
1!
1%
#275880000000
0!
0%
#275885000000
1!
1%
#275890000000
0!
0%
#275895000000
1!
1%
#275900000000
0!
0%
#275905000000
1!
1%
#275910000000
0!
0%
#275915000000
1!
1%
#275920000000
0!
0%
#275925000000
1!
1%
#275930000000
0!
0%
#275935000000
1!
1%
#275940000000
0!
0%
#275945000000
1!
1%
#275950000000
0!
0%
#275955000000
1!
1%
#275960000000
0!
0%
#275965000000
1!
1%
#275970000000
0!
0%
#275975000000
1!
1%
#275980000000
0!
0%
#275985000000
1!
1%
#275990000000
0!
0%
#275995000000
1!
1%
#276000000000
0!
0%
#276005000000
1!
1%
#276010000000
0!
0%
#276015000000
1!
1%
#276020000000
0!
0%
#276025000000
1!
1%
#276030000000
0!
0%
#276035000000
1!
1%
#276040000000
0!
0%
#276045000000
1!
1%
#276050000000
0!
0%
#276055000000
1!
1%
#276060000000
0!
0%
#276065000000
1!
1%
#276070000000
0!
0%
#276075000000
1!
1%
#276080000000
0!
0%
#276085000000
1!
1%
#276090000000
0!
0%
#276095000000
1!
1%
#276100000000
0!
0%
#276105000000
1!
1%
#276110000000
0!
0%
#276115000000
1!
1%
#276120000000
0!
0%
#276125000000
1!
1%
#276130000000
0!
0%
#276135000000
1!
1%
#276140000000
0!
0%
#276145000000
1!
1%
#276150000000
0!
0%
#276155000000
1!
1%
#276160000000
0!
0%
#276165000000
1!
1%
#276170000000
0!
0%
#276175000000
1!
1%
#276180000000
0!
0%
#276185000000
1!
1%
#276190000000
0!
0%
#276195000000
1!
1%
#276200000000
0!
0%
#276205000000
1!
1%
#276210000000
0!
0%
#276215000000
1!
1%
#276220000000
0!
0%
#276225000000
1!
1%
#276230000000
0!
0%
#276235000000
1!
1%
#276240000000
0!
0%
#276245000000
1!
1%
#276250000000
0!
0%
#276255000000
1!
1%
#276260000000
0!
0%
#276265000000
1!
1%
#276270000000
0!
0%
#276275000000
1!
1%
#276280000000
0!
0%
#276285000000
1!
1%
#276290000000
0!
0%
#276295000000
1!
1%
#276300000000
0!
0%
#276305000000
1!
1%
#276310000000
0!
0%
#276315000000
1!
1%
#276320000000
0!
0%
#276325000000
1!
1%
#276330000000
0!
0%
#276335000000
1!
1%
#276340000000
0!
0%
#276345000000
1!
1%
#276350000000
0!
0%
#276355000000
1!
1%
#276360000000
0!
0%
#276365000000
1!
1%
#276370000000
0!
0%
#276375000000
1!
1%
#276380000000
0!
0%
#276385000000
1!
1%
#276390000000
0!
0%
#276395000000
1!
1%
#276400000000
0!
0%
#276405000000
1!
1%
#276410000000
0!
0%
#276415000000
1!
1%
#276420000000
0!
0%
#276425000000
1!
1%
#276430000000
0!
0%
#276435000000
1!
1%
#276440000000
0!
0%
#276445000000
1!
1%
#276450000000
0!
0%
#276455000000
1!
1%
#276460000000
0!
0%
#276465000000
1!
1%
#276470000000
0!
0%
#276475000000
1!
1%
#276480000000
0!
0%
#276485000000
1!
1%
#276490000000
0!
0%
#276495000000
1!
1%
#276500000000
0!
0%
#276505000000
1!
1%
#276510000000
0!
0%
#276515000000
1!
1%
#276520000000
0!
0%
#276525000000
1!
1%
#276530000000
0!
0%
#276535000000
1!
1%
#276540000000
0!
0%
#276545000000
1!
1%
#276550000000
0!
0%
#276555000000
1!
1%
#276560000000
0!
0%
#276565000000
1!
1%
#276570000000
0!
0%
#276575000000
1!
1%
#276580000000
0!
0%
#276585000000
1!
1%
#276590000000
0!
0%
#276595000000
1!
1%
#276600000000
0!
0%
#276605000000
1!
1%
#276610000000
0!
0%
#276615000000
1!
1%
#276620000000
0!
0%
#276625000000
1!
1%
#276630000000
0!
0%
#276635000000
1!
1%
#276640000000
0!
0%
#276645000000
1!
1%
#276650000000
0!
0%
#276655000000
1!
1%
#276660000000
0!
0%
#276665000000
1!
1%
#276670000000
0!
0%
#276675000000
1!
1%
#276680000000
0!
0%
#276685000000
1!
1%
#276690000000
0!
0%
#276695000000
1!
1%
#276700000000
0!
0%
#276705000000
1!
1%
#276710000000
0!
0%
#276715000000
1!
1%
#276720000000
0!
0%
#276725000000
1!
1%
#276730000000
0!
0%
#276735000000
1!
1%
#276740000000
0!
0%
#276745000000
1!
1%
#276750000000
0!
0%
#276755000000
1!
1%
#276760000000
0!
0%
#276765000000
1!
1%
#276770000000
0!
0%
#276775000000
1!
1%
#276780000000
0!
0%
#276785000000
1!
1%
#276790000000
0!
0%
#276795000000
1!
1%
#276800000000
0!
0%
#276805000000
1!
1%
#276810000000
0!
0%
#276815000000
1!
1%
#276820000000
0!
0%
#276825000000
1!
1%
#276830000000
0!
0%
#276835000000
1!
1%
#276840000000
0!
0%
#276845000000
1!
1%
#276850000000
0!
0%
#276855000000
1!
1%
#276860000000
0!
0%
#276865000000
1!
1%
#276870000000
0!
0%
#276875000000
1!
1%
#276880000000
0!
0%
#276885000000
1!
1%
#276890000000
0!
0%
#276895000000
1!
1%
#276900000000
0!
0%
#276905000000
1!
1%
#276910000000
0!
0%
#276915000000
1!
1%
#276920000000
0!
0%
#276925000000
1!
1%
#276930000000
0!
0%
#276935000000
1!
1%
#276940000000
0!
0%
#276945000000
1!
1%
#276950000000
0!
0%
#276955000000
1!
1%
#276960000000
0!
0%
#276965000000
1!
1%
#276970000000
0!
0%
#276975000000
1!
1%
#276980000000
0!
0%
#276985000000
1!
1%
#276990000000
0!
0%
#276995000000
1!
1%
#277000000000
0!
0%
#277005000000
1!
1%
#277010000000
0!
0%
#277015000000
1!
1%
#277020000000
0!
0%
#277025000000
1!
1%
#277030000000
0!
0%
#277035000000
1!
1%
#277040000000
0!
0%
#277045000000
1!
1%
#277050000000
0!
0%
#277055000000
1!
1%
#277060000000
0!
0%
#277065000000
1!
1%
#277070000000
0!
0%
#277075000000
1!
1%
#277080000000
0!
0%
#277085000000
1!
1%
#277090000000
0!
0%
#277095000000
1!
1%
#277100000000
0!
0%
#277105000000
1!
1%
#277110000000
0!
0%
#277115000000
1!
1%
#277120000000
0!
0%
#277125000000
1!
1%
#277130000000
0!
0%
#277135000000
1!
1%
#277140000000
0!
0%
#277145000000
1!
1%
#277150000000
0!
0%
#277155000000
1!
1%
#277160000000
0!
0%
#277165000000
1!
1%
#277170000000
0!
0%
#277175000000
1!
1%
#277180000000
0!
0%
#277185000000
1!
1%
#277190000000
0!
0%
#277195000000
1!
1%
#277200000000
0!
0%
#277205000000
1!
1%
#277210000000
0!
0%
#277215000000
1!
1%
#277220000000
0!
0%
#277225000000
1!
1%
#277230000000
0!
0%
#277235000000
1!
1%
#277240000000
0!
0%
#277245000000
1!
1%
#277250000000
0!
0%
#277255000000
1!
1%
#277260000000
0!
0%
#277265000000
1!
1%
#277270000000
0!
0%
#277275000000
1!
1%
#277280000000
0!
0%
#277285000000
1!
1%
#277290000000
0!
0%
#277295000000
1!
1%
#277300000000
0!
0%
#277305000000
1!
1%
#277310000000
0!
0%
#277315000000
1!
1%
#277320000000
0!
0%
#277325000000
1!
1%
#277330000000
0!
0%
#277335000000
1!
1%
#277340000000
0!
0%
#277345000000
1!
1%
#277350000000
0!
0%
#277355000000
1!
1%
#277360000000
0!
0%
#277365000000
1!
1%
#277370000000
0!
0%
#277375000000
1!
1%
#277380000000
0!
0%
#277385000000
1!
1%
#277390000000
0!
0%
#277395000000
1!
1%
#277400000000
0!
0%
#277405000000
1!
1%
#277410000000
0!
0%
#277415000000
1!
1%
#277420000000
0!
0%
#277425000000
1!
1%
#277430000000
0!
0%
#277435000000
1!
1%
#277440000000
0!
0%
#277445000000
1!
1%
#277450000000
0!
0%
#277455000000
1!
1%
#277460000000
0!
0%
#277465000000
1!
1%
#277470000000
0!
0%
#277475000000
1!
1%
#277480000000
0!
0%
#277485000000
1!
1%
#277490000000
0!
0%
#277495000000
1!
1%
#277500000000
0!
0%
#277505000000
1!
1%
#277510000000
0!
0%
#277515000000
1!
1%
#277520000000
0!
0%
#277525000000
1!
1%
#277530000000
0!
0%
#277535000000
1!
1%
#277540000000
0!
0%
#277545000000
1!
1%
#277550000000
0!
0%
#277555000000
1!
1%
#277560000000
0!
0%
#277565000000
1!
1%
#277570000000
0!
0%
#277575000000
1!
1%
#277580000000
0!
0%
#277585000000
1!
1%
#277590000000
0!
0%
#277595000000
1!
1%
#277600000000
0!
0%
#277605000000
1!
1%
#277610000000
0!
0%
#277615000000
1!
1%
#277620000000
0!
0%
#277625000000
1!
1%
#277630000000
0!
0%
#277635000000
1!
1%
#277640000000
0!
0%
#277645000000
1!
1%
#277650000000
0!
0%
#277655000000
1!
1%
#277660000000
0!
0%
#277665000000
1!
1%
#277670000000
0!
0%
#277675000000
1!
1%
#277680000000
0!
0%
#277685000000
1!
1%
#277690000000
0!
0%
#277695000000
1!
1%
#277700000000
0!
0%
#277705000000
1!
1%
#277710000000
0!
0%
#277715000000
1!
1%
#277720000000
0!
0%
#277725000000
1!
1%
#277730000000
0!
0%
#277735000000
1!
1%
#277740000000
0!
0%
#277745000000
1!
1%
#277750000000
0!
0%
#277755000000
1!
1%
#277760000000
0!
0%
#277765000000
1!
1%
#277770000000
0!
0%
#277775000000
1!
1%
#277780000000
0!
0%
#277785000000
1!
1%
#277790000000
0!
0%
#277795000000
1!
1%
#277800000000
0!
0%
#277805000000
1!
1%
#277810000000
0!
0%
#277815000000
1!
1%
#277820000000
0!
0%
#277825000000
1!
1%
#277830000000
0!
0%
#277835000000
1!
1%
#277840000000
0!
0%
#277845000000
1!
1%
#277850000000
0!
0%
#277855000000
1!
1%
#277860000000
0!
0%
#277865000000
1!
1%
#277870000000
0!
0%
#277875000000
1!
1%
#277880000000
0!
0%
#277885000000
1!
1%
#277890000000
0!
0%
#277895000000
1!
1%
#277900000000
0!
0%
#277905000000
1!
1%
#277910000000
0!
0%
#277915000000
1!
1%
#277920000000
0!
0%
#277925000000
1!
1%
#277930000000
0!
0%
#277935000000
1!
1%
#277940000000
0!
0%
#277945000000
1!
1%
#277950000000
0!
0%
#277955000000
1!
1%
#277960000000
0!
0%
#277965000000
1!
1%
#277970000000
0!
0%
#277975000000
1!
1%
#277980000000
0!
0%
#277985000000
1!
1%
#277990000000
0!
0%
#277995000000
1!
1%
#278000000000
0!
0%
#278005000000
1!
1%
#278010000000
0!
0%
#278015000000
1!
1%
#278020000000
0!
0%
#278025000000
1!
1%
#278030000000
0!
0%
#278035000000
1!
1%
#278040000000
0!
0%
#278045000000
1!
1%
#278050000000
0!
0%
#278055000000
1!
1%
#278060000000
0!
0%
#278065000000
1!
1%
#278070000000
0!
0%
#278075000000
1!
1%
#278080000000
0!
0%
#278085000000
1!
1%
#278090000000
0!
0%
#278095000000
1!
1%
#278100000000
0!
0%
#278105000000
1!
1%
#278110000000
0!
0%
#278115000000
1!
1%
#278120000000
0!
0%
#278125000000
1!
1%
#278130000000
0!
0%
#278135000000
1!
1%
#278140000000
0!
0%
#278145000000
1!
1%
#278150000000
0!
0%
#278155000000
1!
1%
#278160000000
0!
0%
#278165000000
1!
1%
#278170000000
0!
0%
#278175000000
1!
1%
#278180000000
0!
0%
#278185000000
1!
1%
#278190000000
0!
0%
#278195000000
1!
1%
#278200000000
0!
0%
#278205000000
1!
1%
#278210000000
0!
0%
#278215000000
1!
1%
#278220000000
0!
0%
#278225000000
1!
1%
#278230000000
0!
0%
#278235000000
1!
1%
#278240000000
0!
0%
#278245000000
1!
1%
#278250000000
0!
0%
#278255000000
1!
1%
#278260000000
0!
0%
#278265000000
1!
1%
#278270000000
0!
0%
#278275000000
1!
1%
#278280000000
0!
0%
#278285000000
1!
1%
#278290000000
0!
0%
#278295000000
1!
1%
#278300000000
0!
0%
#278305000000
1!
1%
#278310000000
0!
0%
#278315000000
1!
1%
#278320000000
0!
0%
#278325000000
1!
1%
#278330000000
0!
0%
#278335000000
1!
1%
#278340000000
0!
0%
#278345000000
1!
1%
#278350000000
0!
0%
#278355000000
1!
1%
#278360000000
0!
0%
#278365000000
1!
1%
#278370000000
0!
0%
#278375000000
1!
1%
#278380000000
0!
0%
#278385000000
1!
1%
#278390000000
0!
0%
#278395000000
1!
1%
#278400000000
0!
0%
#278405000000
1!
1%
#278410000000
0!
0%
#278415000000
1!
1%
#278420000000
0!
0%
#278425000000
1!
1%
#278430000000
0!
0%
#278435000000
1!
1%
#278440000000
0!
0%
#278445000000
1!
1%
#278450000000
0!
0%
#278455000000
1!
1%
#278460000000
0!
0%
#278465000000
1!
1%
#278470000000
0!
0%
#278475000000
1!
1%
#278480000000
0!
0%
#278485000000
1!
1%
#278490000000
0!
0%
#278495000000
1!
1%
#278500000000
0!
0%
#278505000000
1!
1%
#278510000000
0!
0%
#278515000000
1!
1%
#278520000000
0!
0%
#278525000000
1!
1%
#278530000000
0!
0%
#278535000000
1!
1%
#278540000000
0!
0%
#278545000000
1!
1%
#278550000000
0!
0%
#278555000000
1!
1%
#278560000000
0!
0%
#278565000000
1!
1%
#278570000000
0!
0%
#278575000000
1!
1%
#278580000000
0!
0%
#278585000000
1!
1%
#278590000000
0!
0%
#278595000000
1!
1%
#278600000000
0!
0%
#278605000000
1!
1%
#278610000000
0!
0%
#278615000000
1!
1%
#278620000000
0!
0%
#278625000000
1!
1%
#278630000000
0!
0%
#278635000000
1!
1%
#278640000000
0!
0%
#278645000000
1!
1%
#278650000000
0!
0%
#278655000000
1!
1%
#278660000000
0!
0%
#278665000000
1!
1%
#278670000000
0!
0%
#278675000000
1!
1%
#278680000000
0!
0%
#278685000000
1!
1%
#278690000000
0!
0%
#278695000000
1!
1%
#278700000000
0!
0%
#278705000000
1!
1%
#278710000000
0!
0%
#278715000000
1!
1%
#278720000000
0!
0%
#278725000000
1!
1%
#278730000000
0!
0%
#278735000000
1!
1%
#278740000000
0!
0%
#278745000000
1!
1%
#278750000000
0!
0%
#278755000000
1!
1%
#278760000000
0!
0%
#278765000000
1!
1%
#278770000000
0!
0%
#278775000000
1!
1%
#278780000000
0!
0%
#278785000000
1!
1%
#278790000000
0!
0%
#278795000000
1!
1%
#278800000000
0!
0%
#278805000000
1!
1%
#278810000000
0!
0%
#278815000000
1!
1%
#278820000000
0!
0%
#278825000000
1!
1%
#278830000000
0!
0%
#278835000000
1!
1%
#278840000000
0!
0%
#278845000000
1!
1%
#278850000000
0!
0%
#278855000000
1!
1%
#278860000000
0!
0%
#278865000000
1!
1%
#278870000000
0!
0%
#278875000000
1!
1%
#278880000000
0!
0%
#278885000000
1!
1%
#278890000000
0!
0%
#278895000000
1!
1%
#278900000000
0!
0%
#278905000000
1!
1%
#278910000000
0!
0%
#278915000000
1!
1%
#278920000000
0!
0%
#278925000000
1!
1%
#278930000000
0!
0%
#278935000000
1!
1%
#278940000000
0!
0%
#278945000000
1!
1%
#278950000000
0!
0%
#278955000000
1!
1%
#278960000000
0!
0%
#278965000000
1!
1%
#278970000000
0!
0%
#278975000000
1!
1%
#278980000000
0!
0%
#278985000000
1!
1%
#278990000000
0!
0%
#278995000000
1!
1%
#279000000000
0!
0%
#279005000000
1!
1%
#279010000000
0!
0%
#279015000000
1!
1%
#279020000000
0!
0%
#279025000000
1!
1%
#279030000000
0!
0%
#279035000000
1!
1%
#279040000000
0!
0%
#279045000000
1!
1%
#279050000000
0!
0%
#279055000000
1!
1%
#279060000000
0!
0%
#279065000000
1!
1%
#279070000000
0!
0%
#279075000000
1!
1%
#279080000000
0!
0%
#279085000000
1!
1%
#279090000000
0!
0%
#279095000000
1!
1%
#279100000000
0!
0%
#279105000000
1!
1%
#279110000000
0!
0%
#279115000000
1!
1%
#279120000000
0!
0%
#279125000000
1!
1%
#279130000000
0!
0%
#279135000000
1!
1%
#279140000000
0!
0%
#279145000000
1!
1%
#279150000000
0!
0%
#279155000000
1!
1%
#279160000000
0!
0%
#279165000000
1!
1%
#279170000000
0!
0%
#279175000000
1!
1%
#279180000000
0!
0%
#279185000000
1!
1%
#279190000000
0!
0%
#279195000000
1!
1%
#279200000000
0!
0%
#279205000000
1!
1%
#279210000000
0!
0%
#279215000000
1!
1%
#279220000000
0!
0%
#279225000000
1!
1%
#279230000000
0!
0%
#279235000000
1!
1%
#279240000000
0!
0%
#279245000000
1!
1%
#279250000000
0!
0%
#279255000000
1!
1%
#279260000000
0!
0%
#279265000000
1!
1%
#279270000000
0!
0%
#279275000000
1!
1%
#279280000000
0!
0%
#279285000000
1!
1%
#279290000000
0!
0%
#279295000000
1!
1%
#279300000000
0!
0%
#279305000000
1!
1%
#279310000000
0!
0%
#279315000000
1!
1%
#279320000000
0!
0%
#279325000000
1!
1%
#279330000000
0!
0%
#279335000000
1!
1%
#279340000000
0!
0%
#279345000000
1!
1%
#279350000000
0!
0%
#279355000000
1!
1%
#279360000000
0!
0%
#279365000000
1!
1%
#279370000000
0!
0%
#279375000000
1!
1%
#279380000000
0!
0%
#279385000000
1!
1%
#279390000000
0!
0%
#279395000000
1!
1%
#279400000000
0!
0%
#279405000000
1!
1%
#279410000000
0!
0%
#279415000000
1!
1%
#279420000000
0!
0%
#279425000000
1!
1%
#279430000000
0!
0%
#279435000000
1!
1%
#279440000000
0!
0%
#279445000000
1!
1%
#279450000000
0!
0%
#279455000000
1!
1%
#279460000000
0!
0%
#279465000000
1!
1%
#279470000000
0!
0%
#279475000000
1!
1%
#279480000000
0!
0%
#279485000000
1!
1%
#279490000000
0!
0%
#279495000000
1!
1%
#279500000000
0!
0%
#279505000000
1!
1%
#279510000000
0!
0%
#279515000000
1!
1%
#279520000000
0!
0%
#279525000000
1!
1%
#279530000000
0!
0%
#279535000000
1!
1%
#279540000000
0!
0%
#279545000000
1!
1%
#279550000000
0!
0%
#279555000000
1!
1%
#279560000000
0!
0%
#279565000000
1!
1%
#279570000000
0!
0%
#279575000000
1!
1%
#279580000000
0!
0%
#279585000000
1!
1%
#279590000000
0!
0%
#279595000000
1!
1%
#279600000000
0!
0%
#279605000000
1!
1%
#279610000000
0!
0%
#279615000000
1!
1%
#279620000000
0!
0%
#279625000000
1!
1%
#279630000000
0!
0%
#279635000000
1!
1%
#279640000000
0!
0%
#279645000000
1!
1%
#279650000000
0!
0%
#279655000000
1!
1%
#279660000000
0!
0%
#279665000000
1!
1%
#279670000000
0!
0%
#279675000000
1!
1%
#279680000000
0!
0%
#279685000000
1!
1%
#279690000000
0!
0%
#279695000000
1!
1%
#279700000000
0!
0%
#279705000000
1!
1%
#279710000000
0!
0%
#279715000000
1!
1%
#279720000000
0!
0%
#279725000000
1!
1%
#279730000000
0!
0%
#279735000000
1!
1%
#279740000000
0!
0%
#279745000000
1!
1%
#279750000000
0!
0%
#279755000000
1!
1%
#279760000000
0!
0%
#279765000000
1!
1%
#279770000000
0!
0%
#279775000000
1!
1%
#279780000000
0!
0%
#279785000000
1!
1%
#279790000000
0!
0%
#279795000000
1!
1%
#279800000000
0!
0%
#279805000000
1!
1%
#279810000000
0!
0%
#279815000000
1!
1%
#279820000000
0!
0%
#279825000000
1!
1%
#279830000000
0!
0%
#279835000000
1!
1%
#279840000000
0!
0%
#279845000000
1!
1%
#279850000000
0!
0%
#279855000000
1!
1%
#279860000000
0!
0%
#279865000000
1!
1%
#279870000000
0!
0%
#279875000000
1!
1%
#279880000000
0!
0%
#279885000000
1!
1%
#279890000000
0!
0%
#279895000000
1!
1%
#279900000000
0!
0%
#279905000000
1!
1%
#279910000000
0!
0%
#279915000000
1!
1%
#279920000000
0!
0%
#279925000000
1!
1%
#279930000000
0!
0%
#279935000000
1!
1%
#279940000000
0!
0%
#279945000000
1!
1%
#279950000000
0!
0%
#279955000000
1!
1%
#279960000000
0!
0%
#279965000000
1!
1%
#279970000000
0!
0%
#279975000000
1!
1%
#279980000000
0!
0%
#279985000000
1!
1%
#279990000000
0!
0%
#279995000000
1!
1%
#280000000000
0!
0%
#280005000000
1!
1%
#280010000000
0!
0%
#280015000000
1!
1%
#280020000000
0!
0%
#280025000000
1!
1%
#280030000000
0!
0%
#280035000000
1!
1%
#280040000000
0!
0%
#280045000000
1!
1%
#280050000000
0!
0%
#280055000000
1!
1%
#280060000000
0!
0%
#280065000000
1!
1%
#280070000000
0!
0%
#280075000000
1!
1%
#280080000000
0!
0%
#280085000000
1!
1%
#280090000000
0!
0%
#280095000000
1!
1%
#280100000000
0!
0%
#280105000000
1!
1%
#280110000000
0!
0%
#280115000000
1!
1%
#280120000000
0!
0%
#280125000000
1!
1%
#280130000000
0!
0%
#280135000000
1!
1%
#280140000000
0!
0%
#280145000000
1!
1%
#280150000000
0!
0%
#280155000000
1!
1%
#280160000000
0!
0%
#280165000000
1!
1%
#280170000000
0!
0%
#280175000000
1!
1%
#280180000000
0!
0%
#280185000000
1!
1%
#280190000000
0!
0%
#280195000000
1!
1%
#280200000000
0!
0%
#280205000000
1!
1%
#280210000000
0!
0%
#280215000000
1!
1%
#280220000000
0!
0%
#280225000000
1!
1%
#280230000000
0!
0%
#280235000000
1!
1%
#280240000000
0!
0%
#280245000000
1!
1%
#280250000000
0!
0%
#280255000000
1!
1%
#280260000000
0!
0%
#280265000000
1!
1%
#280270000000
0!
0%
#280275000000
1!
1%
#280280000000
0!
0%
#280285000000
1!
1%
#280290000000
0!
0%
#280295000000
1!
1%
#280300000000
0!
0%
#280305000000
1!
1%
#280310000000
0!
0%
#280315000000
1!
1%
#280320000000
0!
0%
#280325000000
1!
1%
#280330000000
0!
0%
#280335000000
1!
1%
#280340000000
0!
0%
#280345000000
1!
1%
#280350000000
0!
0%
#280355000000
1!
1%
#280360000000
0!
0%
#280365000000
1!
1%
#280370000000
0!
0%
#280375000000
1!
1%
#280380000000
0!
0%
#280385000000
1!
1%
#280390000000
0!
0%
#280395000000
1!
1%
#280400000000
0!
0%
#280405000000
1!
1%
#280410000000
0!
0%
#280415000000
1!
1%
#280420000000
0!
0%
#280425000000
1!
1%
#280430000000
0!
0%
#280435000000
1!
1%
#280440000000
0!
0%
#280445000000
1!
1%
#280450000000
0!
0%
#280455000000
1!
1%
#280460000000
0!
0%
#280465000000
1!
1%
#280470000000
0!
0%
#280475000000
1!
1%
#280480000000
0!
0%
#280485000000
1!
1%
#280490000000
0!
0%
#280495000000
1!
1%
#280500000000
0!
0%
#280505000000
1!
1%
#280510000000
0!
0%
#280515000000
1!
1%
#280520000000
0!
0%
#280525000000
1!
1%
#280530000000
0!
0%
#280535000000
1!
1%
#280540000000
0!
0%
#280545000000
1!
1%
#280550000000
0!
0%
#280555000000
1!
1%
#280560000000
0!
0%
#280565000000
1!
1%
#280570000000
0!
0%
#280575000000
1!
1%
#280580000000
0!
0%
#280585000000
1!
1%
#280590000000
0!
0%
#280595000000
1!
1%
#280600000000
0!
0%
#280605000000
1!
1%
#280610000000
0!
0%
#280615000000
1!
1%
#280620000000
0!
0%
#280625000000
1!
1%
#280630000000
0!
0%
#280635000000
1!
1%
#280640000000
0!
0%
#280645000000
1!
1%
#280650000000
0!
0%
#280655000000
1!
1%
#280660000000
0!
0%
#280665000000
1!
1%
#280670000000
0!
0%
#280675000000
1!
1%
#280680000000
0!
0%
#280685000000
1!
1%
#280690000000
0!
0%
#280695000000
1!
1%
#280700000000
0!
0%
#280705000000
1!
1%
#280710000000
0!
0%
#280715000000
1!
1%
#280720000000
0!
0%
#280725000000
1!
1%
#280730000000
0!
0%
#280735000000
1!
1%
#280740000000
0!
0%
#280745000000
1!
1%
#280750000000
0!
0%
#280755000000
1!
1%
#280760000000
0!
0%
#280765000000
1!
1%
#280770000000
0!
0%
#280775000000
1!
1%
#280780000000
0!
0%
#280785000000
1!
1%
#280790000000
0!
0%
#280795000000
1!
1%
#280800000000
0!
0%
#280805000000
1!
1%
#280810000000
0!
0%
#280815000000
1!
1%
#280820000000
0!
0%
#280825000000
1!
1%
#280830000000
0!
0%
#280835000000
1!
1%
#280840000000
0!
0%
#280845000000
1!
1%
#280850000000
0!
0%
#280855000000
1!
1%
#280860000000
0!
0%
#280865000000
1!
1%
#280870000000
0!
0%
#280875000000
1!
1%
#280880000000
0!
0%
#280885000000
1!
1%
#280890000000
0!
0%
#280895000000
1!
1%
#280900000000
0!
0%
#280905000000
1!
1%
#280910000000
0!
0%
#280915000000
1!
1%
#280920000000
0!
0%
#280925000000
1!
1%
#280930000000
0!
0%
#280935000000
1!
1%
#280940000000
0!
0%
#280945000000
1!
1%
#280950000000
0!
0%
#280955000000
1!
1%
#280960000000
0!
0%
#280965000000
1!
1%
#280970000000
0!
0%
#280975000000
1!
1%
#280980000000
0!
0%
#280985000000
1!
1%
#280990000000
0!
0%
#280995000000
1!
1%
#281000000000
0!
0%
#281005000000
1!
1%
#281010000000
0!
0%
#281015000000
1!
1%
#281020000000
0!
0%
#281025000000
1!
1%
#281030000000
0!
0%
#281035000000
1!
1%
#281040000000
0!
0%
#281045000000
1!
1%
#281050000000
0!
0%
#281055000000
1!
1%
#281060000000
0!
0%
#281065000000
1!
1%
#281070000000
0!
0%
#281075000000
1!
1%
#281080000000
0!
0%
#281085000000
1!
1%
#281090000000
0!
0%
#281095000000
1!
1%
#281100000000
0!
0%
#281105000000
1!
1%
#281110000000
0!
0%
#281115000000
1!
1%
#281120000000
0!
0%
#281125000000
1!
1%
#281130000000
0!
0%
#281135000000
1!
1%
#281140000000
0!
0%
#281145000000
1!
1%
#281150000000
0!
0%
#281155000000
1!
1%
#281160000000
0!
0%
#281165000000
1!
1%
#281170000000
0!
0%
#281175000000
1!
1%
#281180000000
0!
0%
#281185000000
1!
1%
#281190000000
0!
0%
#281195000000
1!
1%
#281200000000
0!
0%
#281205000000
1!
1%
#281210000000
0!
0%
#281215000000
1!
1%
#281220000000
0!
0%
#281225000000
1!
1%
#281230000000
0!
0%
#281235000000
1!
1%
#281240000000
0!
0%
#281245000000
1!
1%
#281250000000
0!
0%
#281255000000
1!
1%
#281260000000
0!
0%
#281265000000
1!
1%
#281270000000
0!
0%
#281275000000
1!
1%
#281280000000
0!
0%
#281285000000
1!
1%
#281290000000
0!
0%
#281295000000
1!
1%
#281300000000
0!
0%
#281305000000
1!
1%
#281310000000
0!
0%
#281315000000
1!
1%
#281320000000
0!
0%
#281325000000
1!
1%
#281330000000
0!
0%
#281335000000
1!
1%
#281340000000
0!
0%
#281345000000
1!
1%
#281350000000
0!
0%
#281355000000
1!
1%
#281360000000
0!
0%
#281365000000
1!
1%
#281370000000
0!
0%
#281375000000
1!
1%
#281380000000
0!
0%
#281385000000
1!
1%
#281390000000
0!
0%
#281395000000
1!
1%
#281400000000
0!
0%
#281405000000
1!
1%
#281410000000
0!
0%
#281415000000
1!
1%
#281420000000
0!
0%
#281425000000
1!
1%
#281430000000
0!
0%
#281435000000
1!
1%
#281440000000
0!
0%
#281445000000
1!
1%
#281450000000
0!
0%
#281455000000
1!
1%
#281460000000
0!
0%
#281465000000
1!
1%
#281470000000
0!
0%
#281475000000
1!
1%
#281480000000
0!
0%
#281485000000
1!
1%
#281490000000
0!
0%
#281495000000
1!
1%
#281500000000
0!
0%
#281505000000
1!
1%
#281510000000
0!
0%
#281515000000
1!
1%
#281520000000
0!
0%
#281525000000
1!
1%
#281530000000
0!
0%
#281535000000
1!
1%
#281540000000
0!
0%
#281545000000
1!
1%
#281550000000
0!
0%
#281555000000
1!
1%
#281560000000
0!
0%
#281565000000
1!
1%
#281570000000
0!
0%
#281575000000
1!
1%
#281580000000
0!
0%
#281585000000
1!
1%
#281590000000
0!
0%
#281595000000
1!
1%
#281600000000
0!
0%
#281605000000
1!
1%
#281610000000
0!
0%
#281615000000
1!
1%
#281620000000
0!
0%
#281625000000
1!
1%
#281630000000
0!
0%
#281635000000
1!
1%
#281640000000
0!
0%
#281645000000
1!
1%
#281650000000
0!
0%
#281655000000
1!
1%
#281660000000
0!
0%
#281665000000
1!
1%
#281670000000
0!
0%
#281675000000
1!
1%
#281680000000
0!
0%
#281685000000
1!
1%
#281690000000
0!
0%
#281695000000
1!
1%
#281700000000
0!
0%
#281705000000
1!
1%
#281710000000
0!
0%
#281715000000
1!
1%
#281720000000
0!
0%
#281725000000
1!
1%
#281730000000
0!
0%
#281735000000
1!
1%
#281740000000
0!
0%
#281745000000
1!
1%
#281750000000
0!
0%
#281755000000
1!
1%
#281760000000
0!
0%
#281765000000
1!
1%
#281770000000
0!
0%
#281775000000
1!
1%
#281780000000
0!
0%
#281785000000
1!
1%
#281790000000
0!
0%
#281795000000
1!
1%
#281800000000
0!
0%
#281805000000
1!
1%
#281810000000
0!
0%
#281815000000
1!
1%
#281820000000
0!
0%
#281825000000
1!
1%
#281830000000
0!
0%
#281835000000
1!
1%
#281840000000
0!
0%
#281845000000
1!
1%
#281850000000
0!
0%
#281855000000
1!
1%
#281860000000
0!
0%
#281865000000
1!
1%
#281870000000
0!
0%
#281875000000
1!
1%
#281880000000
0!
0%
#281885000000
1!
1%
#281890000000
0!
0%
#281895000000
1!
1%
#281900000000
0!
0%
#281905000000
1!
1%
#281910000000
0!
0%
#281915000000
1!
1%
#281920000000
0!
0%
#281925000000
1!
1%
#281930000000
0!
0%
#281935000000
1!
1%
#281940000000
0!
0%
#281945000000
1!
1%
#281950000000
0!
0%
#281955000000
1!
1%
#281960000000
0!
0%
#281965000000
1!
1%
#281970000000
0!
0%
#281975000000
1!
1%
#281980000000
0!
0%
#281985000000
1!
1%
#281990000000
0!
0%
#281995000000
1!
1%
#282000000000
0!
0%
#282005000000
1!
1%
#282010000000
0!
0%
#282015000000
1!
1%
#282020000000
0!
0%
#282025000000
1!
1%
#282030000000
0!
0%
#282035000000
1!
1%
#282040000000
0!
0%
#282045000000
1!
1%
#282050000000
0!
0%
#282055000000
1!
1%
#282060000000
0!
0%
#282065000000
1!
1%
#282070000000
0!
0%
#282075000000
1!
1%
#282080000000
0!
0%
#282085000000
1!
1%
#282090000000
0!
0%
#282095000000
1!
1%
#282100000000
0!
0%
#282105000000
1!
1%
#282110000000
0!
0%
#282115000000
1!
1%
#282120000000
0!
0%
#282125000000
1!
1%
#282130000000
0!
0%
#282135000000
1!
1%
#282140000000
0!
0%
#282145000000
1!
1%
#282150000000
0!
0%
#282155000000
1!
1%
#282160000000
0!
0%
#282165000000
1!
1%
#282170000000
0!
0%
#282175000000
1!
1%
#282180000000
0!
0%
#282185000000
1!
1%
#282190000000
0!
0%
#282195000000
1!
1%
#282200000000
0!
0%
#282205000000
1!
1%
#282210000000
0!
0%
#282215000000
1!
1%
#282220000000
0!
0%
#282225000000
1!
1%
#282230000000
0!
0%
#282235000000
1!
1%
#282240000000
0!
0%
#282245000000
1!
1%
#282250000000
0!
0%
#282255000000
1!
1%
#282260000000
0!
0%
#282265000000
1!
1%
#282270000000
0!
0%
#282275000000
1!
1%
#282280000000
0!
0%
#282285000000
1!
1%
#282290000000
0!
0%
#282295000000
1!
1%
#282300000000
0!
0%
#282305000000
1!
1%
#282310000000
0!
0%
#282315000000
1!
1%
#282320000000
0!
0%
#282325000000
1!
1%
#282330000000
0!
0%
#282335000000
1!
1%
#282340000000
0!
0%
#282345000000
1!
1%
#282350000000
0!
0%
#282355000000
1!
1%
#282360000000
0!
0%
#282365000000
1!
1%
#282370000000
0!
0%
#282375000000
1!
1%
#282380000000
0!
0%
#282385000000
1!
1%
#282390000000
0!
0%
#282395000000
1!
1%
#282400000000
0!
0%
#282405000000
1!
1%
#282410000000
0!
0%
#282415000000
1!
1%
#282420000000
0!
0%
#282425000000
1!
1%
#282430000000
0!
0%
#282435000000
1!
1%
#282440000000
0!
0%
#282445000000
1!
1%
#282450000000
0!
0%
#282455000000
1!
1%
#282460000000
0!
0%
#282465000000
1!
1%
#282470000000
0!
0%
#282475000000
1!
1%
#282480000000
0!
0%
#282485000000
1!
1%
#282490000000
0!
0%
#282495000000
1!
1%
#282500000000
0!
0%
#282505000000
1!
1%
#282510000000
0!
0%
#282515000000
1!
1%
#282520000000
0!
0%
#282525000000
1!
1%
#282530000000
0!
0%
#282535000000
1!
1%
#282540000000
0!
0%
#282545000000
1!
1%
#282550000000
0!
0%
#282555000000
1!
1%
#282560000000
0!
0%
#282565000000
1!
1%
#282570000000
0!
0%
#282575000000
1!
1%
#282580000000
0!
0%
#282585000000
1!
1%
#282590000000
0!
0%
#282595000000
1!
1%
#282600000000
0!
0%
#282605000000
1!
1%
#282610000000
0!
0%
#282615000000
1!
1%
#282620000000
0!
0%
#282625000000
1!
1%
#282630000000
0!
0%
#282635000000
1!
1%
#282640000000
0!
0%
#282645000000
1!
1%
#282650000000
0!
0%
#282655000000
1!
1%
#282660000000
0!
0%
#282665000000
1!
1%
#282670000000
0!
0%
#282675000000
1!
1%
#282680000000
0!
0%
#282685000000
1!
1%
#282690000000
0!
0%
#282695000000
1!
1%
#282700000000
0!
0%
#282705000000
1!
1%
#282710000000
0!
0%
#282715000000
1!
1%
#282720000000
0!
0%
#282725000000
1!
1%
#282730000000
0!
0%
#282735000000
1!
1%
#282740000000
0!
0%
#282745000000
1!
1%
#282750000000
0!
0%
#282755000000
1!
1%
#282760000000
0!
0%
#282765000000
1!
1%
#282770000000
0!
0%
#282775000000
1!
1%
#282780000000
0!
0%
#282785000000
1!
1%
#282790000000
0!
0%
#282795000000
1!
1%
#282800000000
0!
0%
#282805000000
1!
1%
#282810000000
0!
0%
#282815000000
1!
1%
#282820000000
0!
0%
#282825000000
1!
1%
#282830000000
0!
0%
#282835000000
1!
1%
#282840000000
0!
0%
#282845000000
1!
1%
#282850000000
0!
0%
#282855000000
1!
1%
#282860000000
0!
0%
#282865000000
1!
1%
#282870000000
0!
0%
#282875000000
1!
1%
#282880000000
0!
0%
#282885000000
1!
1%
#282890000000
0!
0%
#282895000000
1!
1%
#282900000000
0!
0%
#282905000000
1!
1%
#282910000000
0!
0%
#282915000000
1!
1%
#282920000000
0!
0%
#282925000000
1!
1%
#282930000000
0!
0%
#282935000000
1!
1%
#282940000000
0!
0%
#282945000000
1!
1%
#282950000000
0!
0%
#282955000000
1!
1%
#282960000000
0!
0%
#282965000000
1!
1%
#282970000000
0!
0%
#282975000000
1!
1%
#282980000000
0!
0%
#282985000000
1!
1%
#282990000000
0!
0%
#282995000000
1!
1%
#283000000000
0!
0%
#283005000000
1!
1%
#283010000000
0!
0%
#283015000000
1!
1%
#283020000000
0!
0%
#283025000000
1!
1%
#283030000000
0!
0%
#283035000000
1!
1%
#283040000000
0!
0%
#283045000000
1!
1%
#283050000000
0!
0%
#283055000000
1!
1%
#283060000000
0!
0%
#283065000000
1!
1%
#283070000000
0!
0%
#283075000000
1!
1%
#283080000000
0!
0%
#283085000000
1!
1%
#283090000000
0!
0%
#283095000000
1!
1%
#283100000000
0!
0%
#283105000000
1!
1%
#283110000000
0!
0%
#283115000000
1!
1%
#283120000000
0!
0%
#283125000000
1!
1%
#283130000000
0!
0%
#283135000000
1!
1%
#283140000000
0!
0%
#283145000000
1!
1%
#283150000000
0!
0%
#283155000000
1!
1%
#283160000000
0!
0%
#283165000000
1!
1%
#283170000000
0!
0%
#283175000000
1!
1%
#283180000000
0!
0%
#283185000000
1!
1%
#283190000000
0!
0%
#283195000000
1!
1%
#283200000000
0!
0%
#283205000000
1!
1%
#283210000000
0!
0%
#283215000000
1!
1%
#283220000000
0!
0%
#283225000000
1!
1%
#283230000000
0!
0%
#283235000000
1!
1%
#283240000000
0!
0%
#283245000000
1!
1%
#283250000000
0!
0%
#283255000000
1!
1%
#283260000000
0!
0%
#283265000000
1!
1%
#283270000000
0!
0%
#283275000000
1!
1%
#283280000000
0!
0%
#283285000000
1!
1%
#283290000000
0!
0%
#283295000000
1!
1%
#283300000000
0!
0%
#283305000000
1!
1%
#283310000000
0!
0%
#283315000000
1!
1%
#283320000000
0!
0%
#283325000000
1!
1%
#283330000000
0!
0%
#283335000000
1!
1%
#283340000000
0!
0%
#283345000000
1!
1%
#283350000000
0!
0%
#283355000000
1!
1%
#283360000000
0!
0%
#283365000000
1!
1%
#283370000000
0!
0%
#283375000000
1!
1%
#283380000000
0!
0%
#283385000000
1!
1%
#283390000000
0!
0%
#283395000000
1!
1%
#283400000000
0!
0%
#283405000000
1!
1%
#283410000000
0!
0%
#283415000000
1!
1%
#283420000000
0!
0%
#283425000000
1!
1%
#283430000000
0!
0%
#283435000000
1!
1%
#283440000000
0!
0%
#283445000000
1!
1%
#283450000000
0!
0%
#283455000000
1!
1%
#283460000000
0!
0%
#283465000000
1!
1%
#283470000000
0!
0%
#283475000000
1!
1%
#283480000000
0!
0%
#283485000000
1!
1%
#283490000000
0!
0%
#283495000000
1!
1%
#283500000000
0!
0%
#283505000000
1!
1%
#283510000000
0!
0%
#283515000000
1!
1%
#283520000000
0!
0%
#283525000000
1!
1%
#283530000000
0!
0%
#283535000000
1!
1%
#283540000000
0!
0%
#283545000000
1!
1%
#283550000000
0!
0%
#283555000000
1!
1%
#283560000000
0!
0%
#283565000000
1!
1%
#283570000000
0!
0%
#283575000000
1!
1%
#283580000000
0!
0%
#283585000000
1!
1%
#283590000000
0!
0%
#283595000000
1!
1%
#283600000000
0!
0%
#283605000000
1!
1%
#283610000000
0!
0%
#283615000000
1!
1%
#283620000000
0!
0%
#283625000000
1!
1%
#283630000000
0!
0%
#283635000000
1!
1%
#283640000000
0!
0%
#283645000000
1!
1%
#283650000000
0!
0%
#283655000000
1!
1%
#283660000000
0!
0%
#283665000000
1!
1%
#283670000000
0!
0%
#283675000000
1!
1%
#283680000000
0!
0%
#283685000000
1!
1%
#283690000000
0!
0%
#283695000000
1!
1%
#283700000000
0!
0%
#283705000000
1!
1%
#283710000000
0!
0%
#283715000000
1!
1%
#283720000000
0!
0%
#283725000000
1!
1%
#283730000000
0!
0%
#283735000000
1!
1%
#283740000000
0!
0%
#283745000000
1!
1%
#283750000000
0!
0%
#283755000000
1!
1%
#283760000000
0!
0%
#283765000000
1!
1%
#283770000000
0!
0%
#283775000000
1!
1%
#283780000000
0!
0%
#283785000000
1!
1%
#283790000000
0!
0%
#283795000000
1!
1%
#283800000000
0!
0%
#283805000000
1!
1%
#283810000000
0!
0%
#283815000000
1!
1%
#283820000000
0!
0%
#283825000000
1!
1%
#283830000000
0!
0%
#283835000000
1!
1%
#283840000000
0!
0%
#283845000000
1!
1%
#283850000000
0!
0%
#283855000000
1!
1%
#283860000000
0!
0%
#283865000000
1!
1%
#283870000000
0!
0%
#283875000000
1!
1%
#283880000000
0!
0%
#283885000000
1!
1%
#283890000000
0!
0%
#283895000000
1!
1%
#283900000000
0!
0%
#283905000000
1!
1%
#283910000000
0!
0%
#283915000000
1!
1%
#283920000000
0!
0%
#283925000000
1!
1%
#283930000000
0!
0%
#283935000000
1!
1%
#283940000000
0!
0%
#283945000000
1!
1%
#283950000000
0!
0%
#283955000000
1!
1%
#283960000000
0!
0%
#283965000000
1!
1%
#283970000000
0!
0%
#283975000000
1!
1%
#283980000000
0!
0%
#283985000000
1!
1%
#283990000000
0!
0%
#283995000000
1!
1%
#284000000000
0!
0%
#284005000000
1!
1%
#284010000000
0!
0%
#284015000000
1!
1%
#284020000000
0!
0%
#284025000000
1!
1%
#284030000000
0!
0%
#284035000000
1!
1%
#284040000000
0!
0%
#284045000000
1!
1%
#284050000000
0!
0%
#284055000000
1!
1%
#284060000000
0!
0%
#284065000000
1!
1%
#284070000000
0!
0%
#284075000000
1!
1%
#284080000000
0!
0%
#284085000000
1!
1%
#284090000000
0!
0%
#284095000000
1!
1%
#284100000000
0!
0%
#284105000000
1!
1%
#284110000000
0!
0%
#284115000000
1!
1%
#284120000000
0!
0%
#284125000000
1!
1%
#284130000000
0!
0%
#284135000000
1!
1%
#284140000000
0!
0%
#284145000000
1!
1%
#284150000000
0!
0%
#284155000000
1!
1%
#284160000000
0!
0%
#284165000000
1!
1%
#284170000000
0!
0%
#284175000000
1!
1%
#284180000000
0!
0%
#284185000000
1!
1%
#284190000000
0!
0%
#284195000000
1!
1%
#284200000000
0!
0%
#284205000000
1!
1%
#284210000000
0!
0%
#284215000000
1!
1%
#284220000000
0!
0%
#284225000000
1!
1%
#284230000000
0!
0%
#284235000000
1!
1%
#284240000000
0!
0%
#284245000000
1!
1%
#284250000000
0!
0%
#284255000000
1!
1%
#284260000000
0!
0%
#284265000000
1!
1%
#284270000000
0!
0%
#284275000000
1!
1%
#284280000000
0!
0%
#284285000000
1!
1%
#284290000000
0!
0%
#284295000000
1!
1%
#284300000000
0!
0%
#284305000000
1!
1%
#284310000000
0!
0%
#284315000000
1!
1%
#284320000000
0!
0%
#284325000000
1!
1%
#284330000000
0!
0%
#284335000000
1!
1%
#284340000000
0!
0%
#284345000000
1!
1%
#284350000000
0!
0%
#284355000000
1!
1%
#284360000000
0!
0%
#284365000000
1!
1%
#284370000000
0!
0%
#284375000000
1!
1%
#284380000000
0!
0%
#284385000000
1!
1%
#284390000000
0!
0%
#284395000000
1!
1%
#284400000000
0!
0%
#284405000000
1!
1%
#284410000000
0!
0%
#284415000000
1!
1%
#284420000000
0!
0%
#284425000000
1!
1%
#284430000000
0!
0%
#284435000000
1!
1%
#284440000000
0!
0%
#284445000000
1!
1%
#284450000000
0!
0%
#284455000000
1!
1%
#284460000000
0!
0%
#284465000000
1!
1%
#284470000000
0!
0%
#284475000000
1!
1%
#284480000000
0!
0%
#284485000000
1!
1%
#284490000000
0!
0%
#284495000000
1!
1%
#284500000000
0!
0%
#284505000000
1!
1%
#284510000000
0!
0%
#284515000000
1!
1%
#284520000000
0!
0%
#284525000000
1!
1%
#284530000000
0!
0%
#284535000000
1!
1%
#284540000000
0!
0%
#284545000000
1!
1%
#284550000000
0!
0%
#284555000000
1!
1%
#284560000000
0!
0%
#284565000000
1!
1%
#284570000000
0!
0%
#284575000000
1!
1%
#284580000000
0!
0%
#284585000000
1!
1%
#284590000000
0!
0%
#284595000000
1!
1%
#284600000000
0!
0%
#284605000000
1!
1%
#284610000000
0!
0%
#284615000000
1!
1%
#284620000000
0!
0%
#284625000000
1!
1%
#284630000000
0!
0%
#284635000000
1!
1%
#284640000000
0!
0%
#284645000000
1!
1%
#284650000000
0!
0%
#284655000000
1!
1%
#284660000000
0!
0%
#284665000000
1!
1%
#284670000000
0!
0%
#284675000000
1!
1%
#284680000000
0!
0%
#284685000000
1!
1%
#284690000000
0!
0%
#284695000000
1!
1%
#284700000000
0!
0%
#284705000000
1!
1%
#284710000000
0!
0%
#284715000000
1!
1%
#284720000000
0!
0%
#284725000000
1!
1%
#284730000000
0!
0%
#284735000000
1!
1%
#284740000000
0!
0%
#284745000000
1!
1%
#284750000000
0!
0%
#284755000000
1!
1%
#284760000000
0!
0%
#284765000000
1!
1%
#284770000000
0!
0%
#284775000000
1!
1%
#284780000000
0!
0%
#284785000000
1!
1%
#284790000000
0!
0%
#284795000000
1!
1%
#284800000000
0!
0%
#284805000000
1!
1%
#284810000000
0!
0%
#284815000000
1!
1%
#284820000000
0!
0%
#284825000000
1!
1%
#284830000000
0!
0%
#284835000000
1!
1%
#284840000000
0!
0%
#284845000000
1!
1%
#284850000000
0!
0%
#284855000000
1!
1%
#284860000000
0!
0%
#284865000000
1!
1%
#284870000000
0!
0%
#284875000000
1!
1%
#284880000000
0!
0%
#284885000000
1!
1%
#284890000000
0!
0%
#284895000000
1!
1%
#284900000000
0!
0%
#284905000000
1!
1%
#284910000000
0!
0%
#284915000000
1!
1%
#284920000000
0!
0%
#284925000000
1!
1%
#284930000000
0!
0%
#284935000000
1!
1%
#284940000000
0!
0%
#284945000000
1!
1%
#284950000000
0!
0%
#284955000000
1!
1%
#284960000000
0!
0%
#284965000000
1!
1%
#284970000000
0!
0%
#284975000000
1!
1%
#284980000000
0!
0%
#284985000000
1!
1%
#284990000000
0!
0%
#284995000000
1!
1%
#285000000000
0!
0%
#285005000000
1!
1%
#285010000000
0!
0%
#285015000000
1!
1%
#285020000000
0!
0%
#285025000000
1!
1%
#285030000000
0!
0%
#285035000000
1!
1%
#285040000000
0!
0%
#285045000000
1!
1%
#285050000000
0!
0%
#285055000000
1!
1%
#285060000000
0!
0%
#285065000000
1!
1%
#285070000000
0!
0%
#285075000000
1!
1%
#285080000000
0!
0%
#285085000000
1!
1%
#285090000000
0!
0%
#285095000000
1!
1%
#285100000000
0!
0%
#285105000000
1!
1%
#285110000000
0!
0%
#285115000000
1!
1%
#285120000000
0!
0%
#285125000000
1!
1%
#285130000000
0!
0%
#285135000000
1!
1%
#285140000000
0!
0%
#285145000000
1!
1%
#285150000000
0!
0%
#285155000000
1!
1%
#285160000000
0!
0%
#285165000000
1!
1%
#285170000000
0!
0%
#285175000000
1!
1%
#285180000000
0!
0%
#285185000000
1!
1%
#285190000000
0!
0%
#285195000000
1!
1%
#285200000000
0!
0%
#285205000000
1!
1%
#285210000000
0!
0%
#285215000000
1!
1%
#285220000000
0!
0%
#285225000000
1!
1%
#285230000000
0!
0%
#285235000000
1!
1%
#285240000000
0!
0%
#285245000000
1!
1%
#285250000000
0!
0%
#285255000000
1!
1%
#285260000000
0!
0%
#285265000000
1!
1%
#285270000000
0!
0%
#285275000000
1!
1%
#285280000000
0!
0%
#285285000000
1!
1%
#285290000000
0!
0%
#285295000000
1!
1%
#285300000000
0!
0%
#285305000000
1!
1%
#285310000000
0!
0%
#285315000000
1!
1%
#285320000000
0!
0%
#285325000000
1!
1%
#285330000000
0!
0%
#285335000000
1!
1%
#285340000000
0!
0%
#285345000000
1!
1%
#285350000000
0!
0%
#285355000000
1!
1%
#285360000000
0!
0%
#285365000000
1!
1%
#285370000000
0!
0%
#285375000000
1!
1%
#285380000000
0!
0%
#285385000000
1!
1%
#285390000000
0!
0%
#285395000000
1!
1%
#285400000000
0!
0%
#285405000000
1!
1%
#285410000000
0!
0%
#285415000000
1!
1%
#285420000000
0!
0%
#285425000000
1!
1%
#285430000000
0!
0%
#285435000000
1!
1%
#285440000000
0!
0%
#285445000000
1!
1%
#285450000000
0!
0%
#285455000000
1!
1%
#285460000000
0!
0%
#285465000000
1!
1%
#285470000000
0!
0%
#285475000000
1!
1%
#285480000000
0!
0%
#285485000000
1!
1%
#285490000000
0!
0%
#285495000000
1!
1%
#285500000000
0!
0%
#285505000000
1!
1%
#285510000000
0!
0%
#285515000000
1!
1%
#285520000000
0!
0%
#285525000000
1!
1%
#285530000000
0!
0%
#285535000000
1!
1%
#285540000000
0!
0%
#285545000000
1!
1%
#285550000000
0!
0%
#285555000000
1!
1%
#285560000000
0!
0%
#285565000000
1!
1%
#285570000000
0!
0%
#285575000000
1!
1%
#285580000000
0!
0%
#285585000000
1!
1%
#285590000000
0!
0%
#285595000000
1!
1%
#285600000000
0!
0%
#285605000000
1!
1%
#285610000000
0!
0%
#285615000000
1!
1%
#285620000000
0!
0%
#285625000000
1!
1%
#285630000000
0!
0%
#285635000000
1!
1%
#285640000000
0!
0%
#285645000000
1!
1%
#285650000000
0!
0%
#285655000000
1!
1%
#285660000000
0!
0%
#285665000000
1!
1%
#285670000000
0!
0%
#285675000000
1!
1%
#285680000000
0!
0%
#285685000000
1!
1%
#285690000000
0!
0%
#285695000000
1!
1%
#285700000000
0!
0%
#285705000000
1!
1%
#285710000000
0!
0%
#285715000000
1!
1%
#285720000000
0!
0%
#285725000000
1!
1%
#285730000000
0!
0%
#285735000000
1!
1%
#285740000000
0!
0%
#285745000000
1!
1%
#285750000000
0!
0%
#285755000000
1!
1%
#285760000000
0!
0%
#285765000000
1!
1%
#285770000000
0!
0%
#285775000000
1!
1%
#285780000000
0!
0%
#285785000000
1!
1%
#285790000000
0!
0%
#285795000000
1!
1%
#285800000000
0!
0%
#285805000000
1!
1%
#285810000000
0!
0%
#285815000000
1!
1%
#285820000000
0!
0%
#285825000000
1!
1%
#285830000000
0!
0%
#285835000000
1!
1%
#285840000000
0!
0%
#285845000000
1!
1%
#285850000000
0!
0%
#285855000000
1!
1%
#285860000000
0!
0%
#285865000000
1!
1%
#285870000000
0!
0%
#285875000000
1!
1%
#285880000000
0!
0%
#285885000000
1!
1%
#285890000000
0!
0%
#285895000000
1!
1%
#285900000000
0!
0%
#285905000000
1!
1%
#285910000000
0!
0%
#285915000000
1!
1%
#285920000000
0!
0%
#285925000000
1!
1%
#285930000000
0!
0%
#285935000000
1!
1%
#285940000000
0!
0%
#285945000000
1!
1%
#285950000000
0!
0%
#285955000000
1!
1%
#285960000000
0!
0%
#285965000000
1!
1%
#285970000000
0!
0%
#285975000000
1!
1%
#285980000000
0!
0%
#285985000000
1!
1%
#285990000000
0!
0%
#285995000000
1!
1%
#286000000000
0!
0%
#286005000000
1!
1%
#286010000000
0!
0%
#286015000000
1!
1%
#286020000000
0!
0%
#286025000000
1!
1%
#286030000000
0!
0%
#286035000000
1!
1%
#286040000000
0!
0%
#286045000000
1!
1%
#286050000000
0!
0%
#286055000000
1!
1%
#286060000000
0!
0%
#286065000000
1!
1%
#286070000000
0!
0%
#286075000000
1!
1%
#286080000000
0!
0%
#286085000000
1!
1%
#286090000000
0!
0%
#286095000000
1!
1%
#286100000000
0!
0%
#286105000000
1!
1%
#286110000000
0!
0%
#286115000000
1!
1%
#286120000000
0!
0%
#286125000000
1!
1%
#286130000000
0!
0%
#286135000000
1!
1%
#286140000000
0!
0%
#286145000000
1!
1%
#286150000000
0!
0%
#286155000000
1!
1%
#286160000000
0!
0%
#286165000000
1!
1%
#286170000000
0!
0%
#286175000000
1!
1%
#286180000000
0!
0%
#286185000000
1!
1%
#286190000000
0!
0%
#286195000000
1!
1%
#286200000000
0!
0%
#286205000000
1!
1%
#286210000000
0!
0%
#286215000000
1!
1%
#286220000000
0!
0%
#286225000000
1!
1%
#286230000000
0!
0%
#286235000000
1!
1%
#286240000000
0!
0%
#286245000000
1!
1%
#286250000000
0!
0%
#286255000000
1!
1%
#286260000000
0!
0%
#286265000000
1!
1%
#286270000000
0!
0%
#286275000000
1!
1%
#286280000000
0!
0%
#286285000000
1!
1%
#286290000000
0!
0%
#286295000000
1!
1%
#286300000000
0!
0%
#286305000000
1!
1%
#286310000000
0!
0%
#286315000000
1!
1%
#286320000000
0!
0%
#286325000000
1!
1%
#286330000000
0!
0%
#286335000000
1!
1%
#286340000000
0!
0%
#286345000000
1!
1%
#286350000000
0!
0%
#286355000000
1!
1%
#286360000000
0!
0%
#286365000000
1!
1%
#286370000000
0!
0%
#286375000000
1!
1%
#286380000000
0!
0%
#286385000000
1!
1%
#286390000000
0!
0%
#286395000000
1!
1%
#286400000000
0!
0%
#286405000000
1!
1%
#286410000000
0!
0%
#286415000000
1!
1%
#286420000000
0!
0%
#286425000000
1!
1%
#286430000000
0!
0%
#286435000000
1!
1%
#286440000000
0!
0%
#286445000000
1!
1%
#286450000000
0!
0%
#286455000000
1!
1%
#286460000000
0!
0%
#286465000000
1!
1%
#286470000000
0!
0%
#286475000000
1!
1%
#286480000000
0!
0%
#286485000000
1!
1%
#286490000000
0!
0%
#286495000000
1!
1%
#286500000000
0!
0%
#286505000000
1!
1%
#286510000000
0!
0%
#286515000000
1!
1%
#286520000000
0!
0%
#286525000000
1!
1%
#286530000000
0!
0%
#286535000000
1!
1%
#286540000000
0!
0%
#286545000000
1!
1%
#286550000000
0!
0%
#286555000000
1!
1%
#286560000000
0!
0%
#286565000000
1!
1%
#286570000000
0!
0%
#286575000000
1!
1%
#286580000000
0!
0%
#286585000000
1!
1%
#286590000000
0!
0%
#286595000000
1!
1%
#286600000000
0!
0%
#286605000000
1!
1%
#286610000000
0!
0%
#286615000000
1!
1%
#286620000000
0!
0%
#286625000000
1!
1%
#286630000000
0!
0%
#286635000000
1!
1%
#286640000000
0!
0%
#286645000000
1!
1%
#286650000000
0!
0%
#286655000000
1!
1%
#286660000000
0!
0%
#286665000000
1!
1%
#286670000000
0!
0%
#286675000000
1!
1%
#286680000000
0!
0%
#286685000000
1!
1%
#286690000000
0!
0%
#286695000000
1!
1%
#286700000000
0!
0%
#286705000000
1!
1%
#286710000000
0!
0%
#286715000000
1!
1%
#286720000000
0!
0%
#286725000000
1!
1%
#286730000000
0!
0%
#286735000000
1!
1%
#286740000000
0!
0%
#286745000000
1!
1%
#286750000000
0!
0%
#286755000000
1!
1%
#286760000000
0!
0%
#286765000000
1!
1%
#286770000000
0!
0%
#286775000000
1!
1%
#286780000000
0!
0%
#286785000000
1!
1%
#286790000000
0!
0%
#286795000000
1!
1%
#286800000000
0!
0%
#286805000000
1!
1%
#286810000000
0!
0%
#286815000000
1!
1%
#286820000000
0!
0%
#286825000000
1!
1%
#286830000000
0!
0%
#286835000000
1!
1%
#286840000000
0!
0%
#286845000000
1!
1%
#286850000000
0!
0%
#286855000000
1!
1%
#286860000000
0!
0%
#286865000000
1!
1%
#286870000000
0!
0%
#286875000000
1!
1%
#286880000000
0!
0%
#286885000000
1!
1%
#286890000000
0!
0%
#286895000000
1!
1%
#286900000000
0!
0%
#286905000000
1!
1%
#286910000000
0!
0%
#286915000000
1!
1%
#286920000000
0!
0%
#286925000000
1!
1%
#286930000000
0!
0%
#286935000000
1!
1%
#286940000000
0!
0%
#286945000000
1!
1%
#286950000000
0!
0%
#286955000000
1!
1%
#286960000000
0!
0%
#286965000000
1!
1%
#286970000000
0!
0%
#286975000000
1!
1%
#286980000000
0!
0%
#286985000000
1!
1%
#286990000000
0!
0%
#286995000000
1!
1%
#287000000000
0!
0%
#287005000000
1!
1%
#287010000000
0!
0%
#287015000000
1!
1%
#287020000000
0!
0%
#287025000000
1!
1%
#287030000000
0!
0%
#287035000000
1!
1%
#287040000000
0!
0%
#287045000000
1!
1%
#287050000000
0!
0%
#287055000000
1!
1%
#287060000000
0!
0%
#287065000000
1!
1%
#287070000000
0!
0%
#287075000000
1!
1%
#287080000000
0!
0%
#287085000000
1!
1%
#287090000000
0!
0%
#287095000000
1!
1%
#287100000000
0!
0%
#287105000000
1!
1%
#287110000000
0!
0%
#287115000000
1!
1%
#287120000000
0!
0%
#287125000000
1!
1%
#287130000000
0!
0%
#287135000000
1!
1%
#287140000000
0!
0%
#287145000000
1!
1%
#287150000000
0!
0%
#287155000000
1!
1%
#287160000000
0!
0%
#287165000000
1!
1%
#287170000000
0!
0%
#287175000000
1!
1%
#287180000000
0!
0%
#287185000000
1!
1%
#287190000000
0!
0%
#287195000000
1!
1%
#287200000000
0!
0%
#287205000000
1!
1%
#287210000000
0!
0%
#287215000000
1!
1%
#287220000000
0!
0%
#287225000000
1!
1%
#287230000000
0!
0%
#287235000000
1!
1%
#287240000000
0!
0%
#287245000000
1!
1%
#287250000000
0!
0%
#287255000000
1!
1%
#287260000000
0!
0%
#287265000000
1!
1%
#287270000000
0!
0%
#287275000000
1!
1%
#287280000000
0!
0%
#287285000000
1!
1%
#287290000000
0!
0%
#287295000000
1!
1%
#287300000000
0!
0%
#287305000000
1!
1%
#287310000000
0!
0%
#287315000000
1!
1%
#287320000000
0!
0%
#287325000000
1!
1%
#287330000000
0!
0%
#287335000000
1!
1%
#287340000000
0!
0%
#287345000000
1!
1%
#287350000000
0!
0%
#287355000000
1!
1%
#287360000000
0!
0%
#287365000000
1!
1%
#287370000000
0!
0%
#287375000000
1!
1%
#287380000000
0!
0%
#287385000000
1!
1%
#287390000000
0!
0%
#287395000000
1!
1%
#287400000000
0!
0%
#287405000000
1!
1%
#287410000000
0!
0%
#287415000000
1!
1%
#287420000000
0!
0%
#287425000000
1!
1%
#287430000000
0!
0%
#287435000000
1!
1%
#287440000000
0!
0%
#287445000000
1!
1%
#287450000000
0!
0%
#287455000000
1!
1%
#287460000000
0!
0%
#287465000000
1!
1%
#287470000000
0!
0%
#287475000000
1!
1%
#287480000000
0!
0%
#287485000000
1!
1%
#287490000000
0!
0%
#287495000000
1!
1%
#287500000000
0!
0%
#287505000000
1!
1%
#287510000000
0!
0%
#287515000000
1!
1%
#287520000000
0!
0%
#287525000000
1!
1%
#287530000000
0!
0%
#287535000000
1!
1%
#287540000000
0!
0%
#287545000000
1!
1%
#287550000000
0!
0%
#287555000000
1!
1%
#287560000000
0!
0%
#287565000000
1!
1%
#287570000000
0!
0%
#287575000000
1!
1%
#287580000000
0!
0%
#287585000000
1!
1%
#287590000000
0!
0%
#287595000000
1!
1%
#287600000000
0!
0%
#287605000000
1!
1%
#287610000000
0!
0%
#287615000000
1!
1%
#287620000000
0!
0%
#287625000000
1!
1%
#287630000000
0!
0%
#287635000000
1!
1%
#287640000000
0!
0%
#287645000000
1!
1%
#287650000000
0!
0%
#287655000000
1!
1%
#287660000000
0!
0%
#287665000000
1!
1%
#287670000000
0!
0%
#287675000000
1!
1%
#287680000000
0!
0%
#287685000000
1!
1%
#287690000000
0!
0%
#287695000000
1!
1%
#287700000000
0!
0%
#287705000000
1!
1%
#287710000000
0!
0%
#287715000000
1!
1%
#287720000000
0!
0%
#287725000000
1!
1%
#287730000000
0!
0%
#287735000000
1!
1%
#287740000000
0!
0%
#287745000000
1!
1%
#287750000000
0!
0%
#287755000000
1!
1%
#287760000000
0!
0%
#287765000000
1!
1%
#287770000000
0!
0%
#287775000000
1!
1%
#287780000000
0!
0%
#287785000000
1!
1%
#287790000000
0!
0%
#287795000000
1!
1%
#287800000000
0!
0%
#287805000000
1!
1%
#287810000000
0!
0%
#287815000000
1!
1%
#287820000000
0!
0%
#287825000000
1!
1%
#287830000000
0!
0%
#287835000000
1!
1%
#287840000000
0!
0%
#287845000000
1!
1%
#287850000000
0!
0%
#287855000000
1!
1%
#287860000000
0!
0%
#287865000000
1!
1%
#287870000000
0!
0%
#287875000000
1!
1%
#287880000000
0!
0%
#287885000000
1!
1%
#287890000000
0!
0%
#287895000000
1!
1%
#287900000000
0!
0%
#287905000000
1!
1%
#287910000000
0!
0%
#287915000000
1!
1%
#287920000000
0!
0%
#287925000000
1!
1%
#287930000000
0!
0%
#287935000000
1!
1%
#287940000000
0!
0%
#287945000000
1!
1%
#287950000000
0!
0%
#287955000000
1!
1%
#287960000000
0!
0%
#287965000000
1!
1%
#287970000000
0!
0%
#287975000000
1!
1%
#287980000000
0!
0%
#287985000000
1!
1%
#287990000000
0!
0%
#287995000000
1!
1%
#288000000000
0!
0%
#288005000000
1!
1%
#288010000000
0!
0%
#288015000000
1!
1%
#288020000000
0!
0%
#288025000000
1!
1%
#288030000000
0!
0%
#288035000000
1!
1%
#288040000000
0!
0%
#288045000000
1!
1%
#288050000000
0!
0%
#288055000000
1!
1%
#288060000000
0!
0%
#288065000000
1!
1%
#288070000000
0!
0%
#288075000000
1!
1%
#288080000000
0!
0%
#288085000000
1!
1%
#288090000000
0!
0%
#288095000000
1!
1%
#288100000000
0!
0%
#288105000000
1!
1%
#288110000000
0!
0%
#288115000000
1!
1%
#288120000000
0!
0%
#288125000000
1!
1%
#288130000000
0!
0%
#288135000000
1!
1%
#288140000000
0!
0%
#288145000000
1!
1%
#288150000000
0!
0%
#288155000000
1!
1%
#288160000000
0!
0%
#288165000000
1!
1%
#288170000000
0!
0%
#288175000000
1!
1%
#288180000000
0!
0%
#288185000000
1!
1%
#288190000000
0!
0%
#288195000000
1!
1%
#288200000000
0!
0%
#288205000000
1!
1%
#288210000000
0!
0%
#288215000000
1!
1%
#288220000000
0!
0%
#288225000000
1!
1%
#288230000000
0!
0%
#288235000000
1!
1%
#288240000000
0!
0%
#288245000000
1!
1%
#288250000000
0!
0%
#288255000000
1!
1%
#288260000000
0!
0%
#288265000000
1!
1%
#288270000000
0!
0%
#288275000000
1!
1%
#288280000000
0!
0%
#288285000000
1!
1%
#288290000000
0!
0%
#288295000000
1!
1%
#288300000000
0!
0%
#288305000000
1!
1%
#288310000000
0!
0%
#288315000000
1!
1%
#288320000000
0!
0%
#288325000000
1!
1%
#288330000000
0!
0%
#288335000000
1!
1%
#288340000000
0!
0%
#288345000000
1!
1%
#288350000000
0!
0%
#288355000000
1!
1%
#288360000000
0!
0%
#288365000000
1!
1%
#288370000000
0!
0%
#288375000000
1!
1%
#288380000000
0!
0%
#288385000000
1!
1%
#288390000000
0!
0%
#288395000000
1!
1%
#288400000000
0!
0%
#288405000000
1!
1%
#288410000000
0!
0%
#288415000000
1!
1%
#288420000000
0!
0%
#288425000000
1!
1%
#288430000000
0!
0%
#288435000000
1!
1%
#288440000000
0!
0%
#288445000000
1!
1%
#288450000000
0!
0%
#288455000000
1!
1%
#288460000000
0!
0%
#288465000000
1!
1%
#288470000000
0!
0%
#288475000000
1!
1%
#288480000000
0!
0%
#288485000000
1!
1%
#288490000000
0!
0%
#288495000000
1!
1%
#288500000000
0!
0%
#288505000000
1!
1%
#288510000000
0!
0%
#288515000000
1!
1%
#288520000000
0!
0%
#288525000000
1!
1%
#288530000000
0!
0%
#288535000000
1!
1%
#288540000000
0!
0%
#288545000000
1!
1%
#288550000000
0!
0%
#288555000000
1!
1%
#288560000000
0!
0%
#288565000000
1!
1%
#288570000000
0!
0%
#288575000000
1!
1%
#288580000000
0!
0%
#288585000000
1!
1%
#288590000000
0!
0%
#288595000000
1!
1%
#288600000000
0!
0%
#288605000000
1!
1%
#288610000000
0!
0%
#288615000000
1!
1%
#288620000000
0!
0%
#288625000000
1!
1%
#288630000000
0!
0%
#288635000000
1!
1%
#288640000000
0!
0%
#288645000000
1!
1%
#288650000000
0!
0%
#288655000000
1!
1%
#288660000000
0!
0%
#288665000000
1!
1%
#288670000000
0!
0%
#288675000000
1!
1%
#288680000000
0!
0%
#288685000000
1!
1%
#288690000000
0!
0%
#288695000000
1!
1%
#288700000000
0!
0%
#288705000000
1!
1%
#288710000000
0!
0%
#288715000000
1!
1%
#288720000000
0!
0%
#288725000000
1!
1%
#288730000000
0!
0%
#288735000000
1!
1%
#288740000000
0!
0%
#288745000000
1!
1%
#288750000000
0!
0%
#288755000000
1!
1%
#288760000000
0!
0%
#288765000000
1!
1%
#288770000000
0!
0%
#288775000000
1!
1%
#288780000000
0!
0%
#288785000000
1!
1%
#288790000000
0!
0%
#288795000000
1!
1%
#288800000000
0!
0%
#288805000000
1!
1%
#288810000000
0!
0%
#288815000000
1!
1%
#288820000000
0!
0%
#288825000000
1!
1%
#288830000000
0!
0%
#288835000000
1!
1%
#288840000000
0!
0%
#288845000000
1!
1%
#288850000000
0!
0%
#288855000000
1!
1%
#288860000000
0!
0%
#288865000000
1!
1%
#288870000000
0!
0%
#288875000000
1!
1%
#288880000000
0!
0%
#288885000000
1!
1%
#288890000000
0!
0%
#288895000000
1!
1%
#288900000000
0!
0%
#288905000000
1!
1%
#288910000000
0!
0%
#288915000000
1!
1%
#288920000000
0!
0%
#288925000000
1!
1%
#288930000000
0!
0%
#288935000000
1!
1%
#288940000000
0!
0%
#288945000000
1!
1%
#288950000000
0!
0%
#288955000000
1!
1%
#288960000000
0!
0%
#288965000000
1!
1%
#288970000000
0!
0%
#288975000000
1!
1%
#288980000000
0!
0%
#288985000000
1!
1%
#288990000000
0!
0%
#288995000000
1!
1%
#289000000000
0!
0%
#289005000000
1!
1%
#289010000000
0!
0%
#289015000000
1!
1%
#289020000000
0!
0%
#289025000000
1!
1%
#289030000000
0!
0%
#289035000000
1!
1%
#289040000000
0!
0%
#289045000000
1!
1%
#289050000000
0!
0%
#289055000000
1!
1%
#289060000000
0!
0%
#289065000000
1!
1%
#289070000000
0!
0%
#289075000000
1!
1%
#289080000000
0!
0%
#289085000000
1!
1%
#289090000000
0!
0%
#289095000000
1!
1%
#289100000000
0!
0%
#289105000000
1!
1%
#289110000000
0!
0%
#289115000000
1!
1%
#289120000000
0!
0%
#289125000000
1!
1%
#289130000000
0!
0%
#289135000000
1!
1%
#289140000000
0!
0%
#289145000000
1!
1%
#289150000000
0!
0%
#289155000000
1!
1%
#289160000000
0!
0%
#289165000000
1!
1%
#289170000000
0!
0%
#289175000000
1!
1%
#289180000000
0!
0%
#289185000000
1!
1%
#289190000000
0!
0%
#289195000000
1!
1%
#289200000000
0!
0%
#289205000000
1!
1%
#289210000000
0!
0%
#289215000000
1!
1%
#289220000000
0!
0%
#289225000000
1!
1%
#289230000000
0!
0%
#289235000000
1!
1%
#289240000000
0!
0%
#289245000000
1!
1%
#289250000000
0!
0%
#289255000000
1!
1%
#289260000000
0!
0%
#289265000000
1!
1%
#289270000000
0!
0%
#289275000000
1!
1%
#289280000000
0!
0%
#289285000000
1!
1%
#289290000000
0!
0%
#289295000000
1!
1%
#289300000000
0!
0%
#289305000000
1!
1%
#289310000000
0!
0%
#289315000000
1!
1%
#289320000000
0!
0%
#289325000000
1!
1%
#289330000000
0!
0%
#289335000000
1!
1%
#289340000000
0!
0%
#289345000000
1!
1%
#289350000000
0!
0%
#289355000000
1!
1%
#289360000000
0!
0%
#289365000000
1!
1%
#289370000000
0!
0%
#289375000000
1!
1%
#289380000000
0!
0%
#289385000000
1!
1%
#289390000000
0!
0%
#289395000000
1!
1%
#289400000000
0!
0%
#289405000000
1!
1%
#289410000000
0!
0%
#289415000000
1!
1%
#289420000000
0!
0%
#289425000000
1!
1%
#289430000000
0!
0%
#289435000000
1!
1%
#289440000000
0!
0%
#289445000000
1!
1%
#289450000000
0!
0%
#289455000000
1!
1%
#289460000000
0!
0%
#289465000000
1!
1%
#289470000000
0!
0%
#289475000000
1!
1%
#289480000000
0!
0%
#289485000000
1!
1%
#289490000000
0!
0%
#289495000000
1!
1%
#289500000000
0!
0%
#289505000000
1!
1%
#289510000000
0!
0%
#289515000000
1!
1%
#289520000000
0!
0%
#289525000000
1!
1%
#289530000000
0!
0%
#289535000000
1!
1%
#289540000000
0!
0%
#289545000000
1!
1%
#289550000000
0!
0%
#289555000000
1!
1%
#289560000000
0!
0%
#289565000000
1!
1%
#289570000000
0!
0%
#289575000000
1!
1%
#289580000000
0!
0%
#289585000000
1!
1%
#289590000000
0!
0%
#289595000000
1!
1%
#289600000000
0!
0%
#289605000000
1!
1%
#289610000000
0!
0%
#289615000000
1!
1%
#289620000000
0!
0%
#289625000000
1!
1%
#289630000000
0!
0%
#289635000000
1!
1%
#289640000000
0!
0%
#289645000000
1!
1%
#289650000000
0!
0%
#289655000000
1!
1%
#289660000000
0!
0%
#289665000000
1!
1%
#289670000000
0!
0%
#289675000000
1!
1%
#289680000000
0!
0%
#289685000000
1!
1%
#289690000000
0!
0%
#289695000000
1!
1%
#289700000000
0!
0%
#289705000000
1!
1%
#289710000000
0!
0%
#289715000000
1!
1%
#289720000000
0!
0%
#289725000000
1!
1%
#289730000000
0!
0%
#289735000000
1!
1%
#289740000000
0!
0%
#289745000000
1!
1%
#289750000000
0!
0%
#289755000000
1!
1%
#289760000000
0!
0%
#289765000000
1!
1%
#289770000000
0!
0%
#289775000000
1!
1%
#289780000000
0!
0%
#289785000000
1!
1%
#289790000000
0!
0%
#289795000000
1!
1%
#289800000000
0!
0%
#289805000000
1!
1%
#289810000000
0!
0%
#289815000000
1!
1%
#289820000000
0!
0%
#289825000000
1!
1%
#289830000000
0!
0%
#289835000000
1!
1%
#289840000000
0!
0%
#289845000000
1!
1%
#289850000000
0!
0%
#289855000000
1!
1%
#289860000000
0!
0%
#289865000000
1!
1%
#289870000000
0!
0%
#289875000000
1!
1%
#289880000000
0!
0%
#289885000000
1!
1%
#289890000000
0!
0%
#289895000000
1!
1%
#289900000000
0!
0%
#289905000000
1!
1%
#289910000000
0!
0%
#289915000000
1!
1%
#289920000000
0!
0%
#289925000000
1!
1%
#289930000000
0!
0%
#289935000000
1!
1%
#289940000000
0!
0%
#289945000000
1!
1%
#289950000000
0!
0%
#289955000000
1!
1%
#289960000000
0!
0%
#289965000000
1!
1%
#289970000000
0!
0%
#289975000000
1!
1%
#289980000000
0!
0%
#289985000000
1!
1%
#289990000000
0!
0%
#289995000000
1!
1%
#290000000000
0!
0%
#290005000000
1!
1%
#290010000000
0!
0%
#290015000000
1!
1%
#290020000000
0!
0%
#290025000000
1!
1%
#290030000000
0!
0%
#290035000000
1!
1%
#290040000000
0!
0%
#290045000000
1!
1%
#290050000000
0!
0%
#290055000000
1!
1%
#290060000000
0!
0%
#290065000000
1!
1%
#290070000000
0!
0%
#290075000000
1!
1%
#290080000000
0!
0%
#290085000000
1!
1%
#290090000000
0!
0%
#290095000000
1!
1%
#290100000000
0!
0%
#290105000000
1!
1%
#290110000000
0!
0%
#290115000000
1!
1%
#290120000000
0!
0%
#290125000000
1!
1%
#290130000000
0!
0%
#290135000000
1!
1%
#290140000000
0!
0%
#290145000000
1!
1%
#290150000000
0!
0%
#290155000000
1!
1%
#290160000000
0!
0%
#290165000000
1!
1%
#290170000000
0!
0%
#290175000000
1!
1%
#290180000000
0!
0%
#290185000000
1!
1%
#290190000000
0!
0%
#290195000000
1!
1%
#290200000000
0!
0%
#290205000000
1!
1%
#290210000000
0!
0%
#290215000000
1!
1%
#290220000000
0!
0%
#290225000000
1!
1%
#290230000000
0!
0%
#290235000000
1!
1%
#290240000000
0!
0%
#290245000000
1!
1%
#290250000000
0!
0%
#290255000000
1!
1%
#290260000000
0!
0%
#290265000000
1!
1%
#290270000000
0!
0%
#290275000000
1!
1%
#290280000000
0!
0%
#290285000000
1!
1%
#290290000000
0!
0%
#290295000000
1!
1%
#290300000000
0!
0%
#290305000000
1!
1%
#290310000000
0!
0%
#290315000000
1!
1%
#290320000000
0!
0%
#290325000000
1!
1%
#290330000000
0!
0%
#290335000000
1!
1%
#290340000000
0!
0%
#290345000000
1!
1%
#290350000000
0!
0%
#290355000000
1!
1%
#290360000000
0!
0%
#290365000000
1!
1%
#290370000000
0!
0%
#290375000000
1!
1%
#290380000000
0!
0%
#290385000000
1!
1%
#290390000000
0!
0%
#290395000000
1!
1%
#290400000000
0!
0%
#290405000000
1!
1%
#290410000000
0!
0%
#290415000000
1!
1%
#290420000000
0!
0%
#290425000000
1!
1%
#290430000000
0!
0%
#290435000000
1!
1%
#290440000000
0!
0%
#290445000000
1!
1%
#290450000000
0!
0%
#290455000000
1!
1%
#290460000000
0!
0%
#290465000000
1!
1%
#290470000000
0!
0%
#290475000000
1!
1%
#290480000000
0!
0%
#290485000000
1!
1%
#290490000000
0!
0%
#290495000000
1!
1%
#290500000000
0!
0%
#290505000000
1!
1%
#290510000000
0!
0%
#290515000000
1!
1%
#290520000000
0!
0%
#290525000000
1!
1%
#290530000000
0!
0%
#290535000000
1!
1%
#290540000000
0!
0%
#290545000000
1!
1%
#290550000000
0!
0%
#290555000000
1!
1%
#290560000000
0!
0%
#290565000000
1!
1%
#290570000000
0!
0%
#290575000000
1!
1%
#290580000000
0!
0%
#290585000000
1!
1%
#290590000000
0!
0%
#290595000000
1!
1%
#290600000000
0!
0%
#290605000000
1!
1%
#290610000000
0!
0%
#290615000000
1!
1%
#290620000000
0!
0%
#290625000000
1!
1%
#290630000000
0!
0%
#290635000000
1!
1%
#290640000000
0!
0%
#290645000000
1!
1%
#290650000000
0!
0%
#290655000000
1!
1%
#290660000000
0!
0%
#290665000000
1!
1%
#290670000000
0!
0%
#290675000000
1!
1%
#290680000000
0!
0%
#290685000000
1!
1%
#290690000000
0!
0%
#290695000000
1!
1%
#290700000000
0!
0%
#290705000000
1!
1%
#290710000000
0!
0%
#290715000000
1!
1%
#290720000000
0!
0%
#290725000000
1!
1%
#290730000000
0!
0%
#290735000000
1!
1%
#290740000000
0!
0%
#290745000000
1!
1%
#290750000000
0!
0%
#290755000000
1!
1%
#290760000000
0!
0%
#290765000000
1!
1%
#290770000000
0!
0%
#290775000000
1!
1%
#290780000000
0!
0%
#290785000000
1!
1%
#290790000000
0!
0%
#290795000000
1!
1%
#290800000000
0!
0%
#290805000000
1!
1%
#290810000000
0!
0%
#290815000000
1!
1%
#290820000000
0!
0%
#290825000000
1!
1%
#290830000000
0!
0%
#290835000000
1!
1%
#290840000000
0!
0%
#290845000000
1!
1%
#290850000000
0!
0%
#290855000000
1!
1%
#290860000000
0!
0%
#290865000000
1!
1%
#290870000000
0!
0%
#290875000000
1!
1%
#290880000000
0!
0%
#290885000000
1!
1%
#290890000000
0!
0%
#290895000000
1!
1%
#290900000000
0!
0%
#290905000000
1!
1%
#290910000000
0!
0%
#290915000000
1!
1%
#290920000000
0!
0%
#290925000000
1!
1%
#290930000000
0!
0%
#290935000000
1!
1%
#290940000000
0!
0%
#290945000000
1!
1%
#290950000000
0!
0%
#290955000000
1!
1%
#290960000000
0!
0%
#290965000000
1!
1%
#290970000000
0!
0%
#290975000000
1!
1%
#290980000000
0!
0%
#290985000000
1!
1%
#290990000000
0!
0%
#290995000000
1!
1%
#291000000000
0!
0%
#291005000000
1!
1%
#291010000000
0!
0%
#291015000000
1!
1%
#291020000000
0!
0%
#291025000000
1!
1%
#291030000000
0!
0%
#291035000000
1!
1%
#291040000000
0!
0%
#291045000000
1!
1%
#291050000000
0!
0%
#291055000000
1!
1%
#291060000000
0!
0%
#291065000000
1!
1%
#291070000000
0!
0%
#291075000000
1!
1%
#291080000000
0!
0%
#291085000000
1!
1%
#291090000000
0!
0%
#291095000000
1!
1%
#291100000000
0!
0%
#291105000000
1!
1%
#291110000000
0!
0%
#291115000000
1!
1%
#291120000000
0!
0%
#291125000000
1!
1%
#291130000000
0!
0%
#291135000000
1!
1%
#291140000000
0!
0%
#291145000000
1!
1%
#291150000000
0!
0%
#291155000000
1!
1%
#291160000000
0!
0%
#291165000000
1!
1%
#291170000000
0!
0%
#291175000000
1!
1%
#291180000000
0!
0%
#291185000000
1!
1%
#291190000000
0!
0%
#291195000000
1!
1%
#291200000000
0!
0%
#291205000000
1!
1%
#291210000000
0!
0%
#291215000000
1!
1%
#291220000000
0!
0%
#291225000000
1!
1%
#291230000000
0!
0%
#291235000000
1!
1%
#291240000000
0!
0%
#291245000000
1!
1%
#291250000000
0!
0%
#291255000000
1!
1%
#291260000000
0!
0%
#291265000000
1!
1%
#291270000000
0!
0%
#291275000000
1!
1%
#291280000000
0!
0%
#291285000000
1!
1%
#291290000000
0!
0%
#291295000000
1!
1%
#291300000000
0!
0%
#291305000000
1!
1%
#291310000000
0!
0%
#291315000000
1!
1%
#291320000000
0!
0%
#291325000000
1!
1%
#291330000000
0!
0%
#291335000000
1!
1%
#291340000000
0!
0%
#291345000000
1!
1%
#291350000000
0!
0%
#291355000000
1!
1%
#291360000000
0!
0%
#291365000000
1!
1%
#291370000000
0!
0%
#291375000000
1!
1%
#291380000000
0!
0%
#291385000000
1!
1%
#291390000000
0!
0%
#291395000000
1!
1%
#291400000000
0!
0%
#291405000000
1!
1%
#291410000000
0!
0%
#291415000000
1!
1%
#291420000000
0!
0%
#291425000000
1!
1%
#291430000000
0!
0%
#291435000000
1!
1%
#291440000000
0!
0%
#291445000000
1!
1%
#291450000000
0!
0%
#291455000000
1!
1%
#291460000000
0!
0%
#291465000000
1!
1%
#291470000000
0!
0%
#291475000000
1!
1%
#291480000000
0!
0%
#291485000000
1!
1%
#291490000000
0!
0%
#291495000000
1!
1%
#291500000000
0!
0%
#291505000000
1!
1%
#291510000000
0!
0%
#291515000000
1!
1%
#291520000000
0!
0%
#291525000000
1!
1%
#291530000000
0!
0%
#291535000000
1!
1%
#291540000000
0!
0%
#291545000000
1!
1%
#291550000000
0!
0%
#291555000000
1!
1%
#291560000000
0!
0%
#291565000000
1!
1%
#291570000000
0!
0%
#291575000000
1!
1%
#291580000000
0!
0%
#291585000000
1!
1%
#291590000000
0!
0%
#291595000000
1!
1%
#291600000000
0!
0%
#291605000000
1!
1%
#291610000000
0!
0%
#291615000000
1!
1%
#291620000000
0!
0%
#291625000000
1!
1%
#291630000000
0!
0%
#291635000000
1!
1%
#291640000000
0!
0%
#291645000000
1!
1%
#291650000000
0!
0%
#291655000000
1!
1%
#291660000000
0!
0%
#291665000000
1!
1%
#291670000000
0!
0%
#291675000000
1!
1%
#291680000000
0!
0%
#291685000000
1!
1%
#291690000000
0!
0%
#291695000000
1!
1%
#291700000000
0!
0%
#291705000000
1!
1%
#291710000000
0!
0%
#291715000000
1!
1%
#291720000000
0!
0%
#291725000000
1!
1%
#291730000000
0!
0%
#291735000000
1!
1%
#291740000000
0!
0%
#291745000000
1!
1%
#291750000000
0!
0%
#291755000000
1!
1%
#291760000000
0!
0%
#291765000000
1!
1%
#291770000000
0!
0%
#291775000000
1!
1%
#291780000000
0!
0%
#291785000000
1!
1%
#291790000000
0!
0%
#291795000000
1!
1%
#291800000000
0!
0%
#291805000000
1!
1%
#291810000000
0!
0%
#291815000000
1!
1%
#291820000000
0!
0%
#291825000000
1!
1%
#291830000000
0!
0%
#291835000000
1!
1%
#291840000000
0!
0%
#291845000000
1!
1%
#291850000000
0!
0%
#291855000000
1!
1%
#291860000000
0!
0%
#291865000000
1!
1%
#291870000000
0!
0%
#291875000000
1!
1%
#291880000000
0!
0%
#291885000000
1!
1%
#291890000000
0!
0%
#291895000000
1!
1%
#291900000000
0!
0%
#291905000000
1!
1%
#291910000000
0!
0%
#291915000000
1!
1%
#291920000000
0!
0%
#291925000000
1!
1%
#291930000000
0!
0%
#291935000000
1!
1%
#291940000000
0!
0%
#291945000000
1!
1%
#291950000000
0!
0%
#291955000000
1!
1%
#291960000000
0!
0%
#291965000000
1!
1%
#291970000000
0!
0%
#291975000000
1!
1%
#291980000000
0!
0%
#291985000000
1!
1%
#291990000000
0!
0%
#291995000000
1!
1%
#292000000000
0!
0%
#292005000000
1!
1%
#292010000000
0!
0%
#292015000000
1!
1%
#292020000000
0!
0%
#292025000000
1!
1%
#292030000000
0!
0%
#292035000000
1!
1%
#292040000000
0!
0%
#292045000000
1!
1%
#292050000000
0!
0%
#292055000000
1!
1%
#292060000000
0!
0%
#292065000000
1!
1%
#292070000000
0!
0%
#292075000000
1!
1%
#292080000000
0!
0%
#292085000000
1!
1%
#292090000000
0!
0%
#292095000000
1!
1%
#292100000000
0!
0%
#292105000000
1!
1%
#292110000000
0!
0%
#292115000000
1!
1%
#292120000000
0!
0%
#292125000000
1!
1%
#292130000000
0!
0%
#292135000000
1!
1%
#292140000000
0!
0%
#292145000000
1!
1%
#292150000000
0!
0%
#292155000000
1!
1%
#292160000000
0!
0%
#292165000000
1!
1%
#292170000000
0!
0%
#292175000000
1!
1%
#292180000000
0!
0%
#292185000000
1!
1%
#292190000000
0!
0%
#292195000000
1!
1%
#292200000000
0!
0%
#292205000000
1!
1%
#292210000000
0!
0%
#292215000000
1!
1%
#292220000000
0!
0%
#292225000000
1!
1%
#292230000000
0!
0%
#292235000000
1!
1%
#292240000000
0!
0%
#292245000000
1!
1%
#292250000000
0!
0%
#292255000000
1!
1%
#292260000000
0!
0%
#292265000000
1!
1%
#292270000000
0!
0%
#292275000000
1!
1%
#292280000000
0!
0%
#292285000000
1!
1%
#292290000000
0!
0%
#292295000000
1!
1%
#292300000000
0!
0%
#292305000000
1!
1%
#292310000000
0!
0%
#292315000000
1!
1%
#292320000000
0!
0%
#292325000000
1!
1%
#292330000000
0!
0%
#292335000000
1!
1%
#292340000000
0!
0%
#292345000000
1!
1%
#292350000000
0!
0%
#292355000000
1!
1%
#292360000000
0!
0%
#292365000000
1!
1%
#292370000000
0!
0%
#292375000000
1!
1%
#292380000000
0!
0%
#292385000000
1!
1%
#292390000000
0!
0%
#292395000000
1!
1%
#292400000000
0!
0%
#292405000000
1!
1%
#292410000000
0!
0%
#292415000000
1!
1%
#292420000000
0!
0%
#292425000000
1!
1%
#292430000000
0!
0%
#292435000000
1!
1%
#292440000000
0!
0%
#292445000000
1!
1%
#292450000000
0!
0%
#292455000000
1!
1%
#292460000000
0!
0%
#292465000000
1!
1%
#292470000000
0!
0%
#292475000000
1!
1%
#292480000000
0!
0%
#292485000000
1!
1%
#292490000000
0!
0%
#292495000000
1!
1%
#292500000000
0!
0%
#292505000000
1!
1%
#292510000000
0!
0%
#292515000000
1!
1%
#292520000000
0!
0%
#292525000000
1!
1%
#292530000000
0!
0%
#292535000000
1!
1%
#292540000000
0!
0%
#292545000000
1!
1%
#292550000000
0!
0%
#292555000000
1!
1%
#292560000000
0!
0%
#292565000000
1!
1%
#292570000000
0!
0%
#292575000000
1!
1%
#292580000000
0!
0%
#292585000000
1!
1%
#292590000000
0!
0%
#292595000000
1!
1%
#292600000000
0!
0%
#292605000000
1!
1%
#292610000000
0!
0%
#292615000000
1!
1%
#292620000000
0!
0%
#292625000000
1!
1%
#292630000000
0!
0%
#292635000000
1!
1%
#292640000000
0!
0%
#292645000000
1!
1%
#292650000000
0!
0%
#292655000000
1!
1%
#292660000000
0!
0%
#292665000000
1!
1%
#292670000000
0!
0%
#292675000000
1!
1%
#292680000000
0!
0%
#292685000000
1!
1%
#292690000000
0!
0%
#292695000000
1!
1%
#292700000000
0!
0%
#292705000000
1!
1%
#292710000000
0!
0%
#292715000000
1!
1%
#292720000000
0!
0%
#292725000000
1!
1%
#292730000000
0!
0%
#292735000000
1!
1%
#292740000000
0!
0%
#292745000000
1!
1%
#292750000000
0!
0%
#292755000000
1!
1%
#292760000000
0!
0%
#292765000000
1!
1%
#292770000000
0!
0%
#292775000000
1!
1%
#292780000000
0!
0%
#292785000000
1!
1%
#292790000000
0!
0%
#292795000000
1!
1%
#292800000000
0!
0%
#292805000000
1!
1%
#292810000000
0!
0%
#292815000000
1!
1%
#292820000000
0!
0%
#292825000000
1!
1%
#292830000000
0!
0%
#292835000000
1!
1%
#292840000000
0!
0%
#292845000000
1!
1%
#292850000000
0!
0%
#292855000000
1!
1%
#292860000000
0!
0%
#292865000000
1!
1%
#292870000000
0!
0%
#292875000000
1!
1%
#292880000000
0!
0%
#292885000000
1!
1%
#292890000000
0!
0%
#292895000000
1!
1%
#292900000000
0!
0%
#292905000000
1!
1%
#292910000000
0!
0%
#292915000000
1!
1%
#292920000000
0!
0%
#292925000000
1!
1%
#292930000000
0!
0%
#292935000000
1!
1%
#292940000000
0!
0%
#292945000000
1!
1%
#292950000000
0!
0%
#292955000000
1!
1%
#292960000000
0!
0%
#292965000000
1!
1%
#292970000000
0!
0%
#292975000000
1!
1%
#292980000000
0!
0%
#292985000000
1!
1%
#292990000000
0!
0%
#292995000000
1!
1%
#293000000000
0!
0%
#293005000000
1!
1%
#293010000000
0!
0%
#293015000000
1!
1%
#293020000000
0!
0%
#293025000000
1!
1%
#293030000000
0!
0%
#293035000000
1!
1%
#293040000000
0!
0%
#293045000000
1!
1%
#293050000000
0!
0%
#293055000000
1!
1%
#293060000000
0!
0%
#293065000000
1!
1%
#293070000000
0!
0%
#293075000000
1!
1%
#293080000000
0!
0%
#293085000000
1!
1%
#293090000000
0!
0%
#293095000000
1!
1%
#293100000000
0!
0%
#293105000000
1!
1%
#293110000000
0!
0%
#293115000000
1!
1%
#293120000000
0!
0%
#293125000000
1!
1%
#293130000000
0!
0%
#293135000000
1!
1%
#293140000000
0!
0%
#293145000000
1!
1%
#293150000000
0!
0%
#293155000000
1!
1%
#293160000000
0!
0%
#293165000000
1!
1%
#293170000000
0!
0%
#293175000000
1!
1%
#293180000000
0!
0%
#293185000000
1!
1%
#293190000000
0!
0%
#293195000000
1!
1%
#293200000000
0!
0%
#293205000000
1!
1%
#293210000000
0!
0%
#293215000000
1!
1%
#293220000000
0!
0%
#293225000000
1!
1%
#293230000000
0!
0%
#293235000000
1!
1%
#293240000000
0!
0%
#293245000000
1!
1%
#293250000000
0!
0%
#293255000000
1!
1%
#293260000000
0!
0%
#293265000000
1!
1%
#293270000000
0!
0%
#293275000000
1!
1%
#293280000000
0!
0%
#293285000000
1!
1%
#293290000000
0!
0%
#293295000000
1!
1%
#293300000000
0!
0%
#293305000000
1!
1%
#293310000000
0!
0%
#293315000000
1!
1%
#293320000000
0!
0%
#293325000000
1!
1%
#293330000000
0!
0%
#293335000000
1!
1%
#293340000000
0!
0%
#293345000000
1!
1%
#293350000000
0!
0%
#293355000000
1!
1%
#293360000000
0!
0%
#293365000000
1!
1%
#293370000000
0!
0%
#293375000000
1!
1%
#293380000000
0!
0%
#293385000000
1!
1%
#293390000000
0!
0%
#293395000000
1!
1%
#293400000000
0!
0%
#293405000000
1!
1%
#293410000000
0!
0%
#293415000000
1!
1%
#293420000000
0!
0%
#293425000000
1!
1%
#293430000000
0!
0%
#293435000000
1!
1%
#293440000000
0!
0%
#293445000000
1!
1%
#293450000000
0!
0%
#293455000000
1!
1%
#293460000000
0!
0%
#293465000000
1!
1%
#293470000000
0!
0%
#293475000000
1!
1%
#293480000000
0!
0%
#293485000000
1!
1%
#293490000000
0!
0%
#293495000000
1!
1%
#293500000000
0!
0%
#293505000000
1!
1%
#293510000000
0!
0%
#293515000000
1!
1%
#293520000000
0!
0%
#293525000000
1!
1%
#293530000000
0!
0%
#293535000000
1!
1%
#293540000000
0!
0%
#293545000000
1!
1%
#293550000000
0!
0%
#293555000000
1!
1%
#293560000000
0!
0%
#293565000000
1!
1%
#293570000000
0!
0%
#293575000000
1!
1%
#293580000000
0!
0%
#293585000000
1!
1%
#293590000000
0!
0%
#293595000000
1!
1%
#293600000000
0!
0%
#293605000000
1!
1%
#293610000000
0!
0%
#293615000000
1!
1%
#293620000000
0!
0%
#293625000000
1!
1%
#293630000000
0!
0%
#293635000000
1!
1%
#293640000000
0!
0%
#293645000000
1!
1%
#293650000000
0!
0%
#293655000000
1!
1%
#293660000000
0!
0%
#293665000000
1!
1%
#293670000000
0!
0%
#293675000000
1!
1%
#293680000000
0!
0%
#293685000000
1!
1%
#293690000000
0!
0%
#293695000000
1!
1%
#293700000000
0!
0%
#293705000000
1!
1%
#293710000000
0!
0%
#293715000000
1!
1%
#293720000000
0!
0%
#293725000000
1!
1%
#293730000000
0!
0%
#293735000000
1!
1%
#293740000000
0!
0%
#293745000000
1!
1%
#293750000000
0!
0%
#293755000000
1!
1%
#293760000000
0!
0%
#293765000000
1!
1%
#293770000000
0!
0%
#293775000000
1!
1%
#293780000000
0!
0%
#293785000000
1!
1%
#293790000000
0!
0%
#293795000000
1!
1%
#293800000000
0!
0%
#293805000000
1!
1%
#293810000000
0!
0%
#293815000000
1!
1%
#293820000000
0!
0%
#293825000000
1!
1%
#293830000000
0!
0%
#293835000000
1!
1%
#293840000000
0!
0%
#293845000000
1!
1%
#293850000000
0!
0%
#293855000000
1!
1%
#293860000000
0!
0%
#293865000000
1!
1%
#293870000000
0!
0%
#293875000000
1!
1%
#293880000000
0!
0%
#293885000000
1!
1%
#293890000000
0!
0%
#293895000000
1!
1%
#293900000000
0!
0%
#293905000000
1!
1%
#293910000000
0!
0%
#293915000000
1!
1%
#293920000000
0!
0%
#293925000000
1!
1%
#293930000000
0!
0%
#293935000000
1!
1%
#293940000000
0!
0%
#293945000000
1!
1%
#293950000000
0!
0%
#293955000000
1!
1%
#293960000000
0!
0%
#293965000000
1!
1%
#293970000000
0!
0%
#293975000000
1!
1%
#293980000000
0!
0%
#293985000000
1!
1%
#293990000000
0!
0%
#293995000000
1!
1%
#294000000000
0!
0%
#294005000000
1!
1%
#294010000000
0!
0%
#294015000000
1!
1%
#294020000000
0!
0%
#294025000000
1!
1%
#294030000000
0!
0%
#294035000000
1!
1%
#294040000000
0!
0%
#294045000000
1!
1%
#294050000000
0!
0%
#294055000000
1!
1%
#294060000000
0!
0%
#294065000000
1!
1%
#294070000000
0!
0%
#294075000000
1!
1%
#294080000000
0!
0%
#294085000000
1!
1%
#294090000000
0!
0%
#294095000000
1!
1%
#294100000000
0!
0%
#294105000000
1!
1%
#294110000000
0!
0%
#294115000000
1!
1%
#294120000000
0!
0%
#294125000000
1!
1%
#294130000000
0!
0%
#294135000000
1!
1%
#294140000000
0!
0%
#294145000000
1!
1%
#294150000000
0!
0%
#294155000000
1!
1%
#294160000000
0!
0%
#294165000000
1!
1%
#294170000000
0!
0%
#294175000000
1!
1%
#294180000000
0!
0%
#294185000000
1!
1%
#294190000000
0!
0%
#294195000000
1!
1%
#294200000000
0!
0%
#294205000000
1!
1%
#294210000000
0!
0%
#294215000000
1!
1%
#294220000000
0!
0%
#294225000000
1!
1%
#294230000000
0!
0%
#294235000000
1!
1%
#294240000000
0!
0%
#294245000000
1!
1%
#294250000000
0!
0%
#294255000000
1!
1%
#294260000000
0!
0%
#294265000000
1!
1%
#294270000000
0!
0%
#294275000000
1!
1%
#294280000000
0!
0%
#294285000000
1!
1%
#294290000000
0!
0%
#294295000000
1!
1%
#294300000000
0!
0%
#294305000000
1!
1%
#294310000000
0!
0%
#294315000000
1!
1%
#294320000000
0!
0%
#294325000000
1!
1%
#294330000000
0!
0%
#294335000000
1!
1%
#294340000000
0!
0%
#294345000000
1!
1%
#294350000000
0!
0%
#294355000000
1!
1%
#294360000000
0!
0%
#294365000000
1!
1%
#294370000000
0!
0%
#294375000000
1!
1%
#294380000000
0!
0%
#294385000000
1!
1%
#294390000000
0!
0%
#294395000000
1!
1%
#294400000000
0!
0%
#294405000000
1!
1%
#294410000000
0!
0%
#294415000000
1!
1%
#294420000000
0!
0%
#294425000000
1!
1%
#294430000000
0!
0%
#294435000000
1!
1%
#294440000000
0!
0%
#294445000000
1!
1%
#294450000000
0!
0%
#294455000000
1!
1%
#294460000000
0!
0%
#294465000000
1!
1%
#294470000000
0!
0%
#294475000000
1!
1%
#294480000000
0!
0%
#294485000000
1!
1%
#294490000000
0!
0%
#294495000000
1!
1%
#294500000000
0!
0%
#294505000000
1!
1%
#294510000000
0!
0%
#294515000000
1!
1%
#294520000000
0!
0%
#294525000000
1!
1%
#294530000000
0!
0%
#294535000000
1!
1%
#294540000000
0!
0%
#294545000000
1!
1%
#294550000000
0!
0%
#294555000000
1!
1%
#294560000000
0!
0%
#294565000000
1!
1%
#294570000000
0!
0%
#294575000000
1!
1%
#294580000000
0!
0%
#294585000000
1!
1%
#294590000000
0!
0%
#294595000000
1!
1%
#294600000000
0!
0%
#294605000000
1!
1%
#294610000000
0!
0%
#294615000000
1!
1%
#294620000000
0!
0%
#294625000000
1!
1%
#294630000000
0!
0%
#294635000000
1!
1%
#294640000000
0!
0%
#294645000000
1!
1%
#294650000000
0!
0%
#294655000000
1!
1%
#294660000000
0!
0%
#294665000000
1!
1%
#294670000000
0!
0%
#294675000000
1!
1%
#294680000000
0!
0%
#294685000000
1!
1%
#294690000000
0!
0%
#294695000000
1!
1%
#294700000000
0!
0%
#294705000000
1!
1%
#294710000000
0!
0%
#294715000000
1!
1%
#294720000000
0!
0%
#294725000000
1!
1%
#294730000000
0!
0%
#294735000000
1!
1%
#294740000000
0!
0%
#294745000000
1!
1%
#294750000000
0!
0%
#294755000000
1!
1%
#294760000000
0!
0%
#294765000000
1!
1%
#294770000000
0!
0%
#294775000000
1!
1%
#294780000000
0!
0%
#294785000000
1!
1%
#294790000000
0!
0%
#294795000000
1!
1%
#294800000000
0!
0%
#294805000000
1!
1%
#294810000000
0!
0%
#294815000000
1!
1%
#294820000000
0!
0%
#294825000000
1!
1%
#294830000000
0!
0%
#294835000000
1!
1%
#294840000000
0!
0%
#294845000000
1!
1%
#294850000000
0!
0%
#294855000000
1!
1%
#294860000000
0!
0%
#294865000000
1!
1%
#294870000000
0!
0%
#294875000000
1!
1%
#294880000000
0!
0%
#294885000000
1!
1%
#294890000000
0!
0%
#294895000000
1!
1%
#294900000000
0!
0%
#294905000000
1!
1%
#294910000000
0!
0%
#294915000000
1!
1%
#294920000000
0!
0%
#294925000000
1!
1%
#294930000000
0!
0%
#294935000000
1!
1%
#294940000000
0!
0%
#294945000000
1!
1%
#294950000000
0!
0%
#294955000000
1!
1%
#294960000000
0!
0%
#294965000000
1!
1%
#294970000000
0!
0%
#294975000000
1!
1%
#294980000000
0!
0%
#294985000000
1!
1%
#294990000000
0!
0%
#294995000000
1!
1%
#295000000000
0!
0%
#295005000000
1!
1%
#295010000000
0!
0%
#295015000000
1!
1%
#295020000000
0!
0%
#295025000000
1!
1%
#295030000000
0!
0%
#295035000000
1!
1%
#295040000000
0!
0%
#295045000000
1!
1%
#295050000000
0!
0%
#295055000000
1!
1%
#295060000000
0!
0%
#295065000000
1!
1%
#295070000000
0!
0%
#295075000000
1!
1%
#295080000000
0!
0%
#295085000000
1!
1%
#295090000000
0!
0%
#295095000000
1!
1%
#295100000000
0!
0%
#295105000000
1!
1%
#295110000000
0!
0%
#295115000000
1!
1%
#295120000000
0!
0%
#295125000000
1!
1%
#295130000000
0!
0%
#295135000000
1!
1%
#295140000000
0!
0%
#295145000000
1!
1%
#295150000000
0!
0%
#295155000000
1!
1%
#295160000000
0!
0%
#295165000000
1!
1%
#295170000000
0!
0%
#295175000000
1!
1%
#295180000000
0!
0%
#295185000000
1!
1%
#295190000000
0!
0%
#295195000000
1!
1%
#295200000000
0!
0%
#295205000000
1!
1%
#295210000000
0!
0%
#295215000000
1!
1%
#295220000000
0!
0%
#295225000000
1!
1%
#295230000000
0!
0%
#295235000000
1!
1%
#295240000000
0!
0%
#295245000000
1!
1%
#295250000000
0!
0%
#295255000000
1!
1%
#295260000000
0!
0%
#295265000000
1!
1%
#295270000000
0!
0%
#295275000000
1!
1%
#295280000000
0!
0%
#295285000000
1!
1%
#295290000000
0!
0%
#295295000000
1!
1%
#295300000000
0!
0%
#295305000000
1!
1%
#295310000000
0!
0%
#295315000000
1!
1%
#295320000000
0!
0%
#295325000000
1!
1%
#295330000000
0!
0%
#295335000000
1!
1%
#295340000000
0!
0%
#295345000000
1!
1%
#295350000000
0!
0%
#295355000000
1!
1%
#295360000000
0!
0%
#295365000000
1!
1%
#295370000000
0!
0%
#295375000000
1!
1%
#295380000000
0!
0%
#295385000000
1!
1%
#295390000000
0!
0%
#295395000000
1!
1%
#295400000000
0!
0%
#295405000000
1!
1%
#295410000000
0!
0%
#295415000000
1!
1%
#295420000000
0!
0%
#295425000000
1!
1%
#295430000000
0!
0%
#295435000000
1!
1%
#295440000000
0!
0%
#295445000000
1!
1%
#295450000000
0!
0%
#295455000000
1!
1%
#295460000000
0!
0%
#295465000000
1!
1%
#295470000000
0!
0%
#295475000000
1!
1%
#295480000000
0!
0%
#295485000000
1!
1%
#295490000000
0!
0%
#295495000000
1!
1%
#295500000000
0!
0%
#295505000000
1!
1%
#295510000000
0!
0%
#295515000000
1!
1%
#295520000000
0!
0%
#295525000000
1!
1%
#295530000000
0!
0%
#295535000000
1!
1%
#295540000000
0!
0%
#295545000000
1!
1%
#295550000000
0!
0%
#295555000000
1!
1%
#295560000000
0!
0%
#295565000000
1!
1%
#295570000000
0!
0%
#295575000000
1!
1%
#295580000000
0!
0%
#295585000000
1!
1%
#295590000000
0!
0%
#295595000000
1!
1%
#295600000000
0!
0%
#295605000000
1!
1%
#295610000000
0!
0%
#295615000000
1!
1%
#295620000000
0!
0%
#295625000000
1!
1%
#295630000000
0!
0%
#295635000000
1!
1%
#295640000000
0!
0%
#295645000000
1!
1%
#295650000000
0!
0%
#295655000000
1!
1%
#295660000000
0!
0%
#295665000000
1!
1%
#295670000000
0!
0%
#295675000000
1!
1%
#295680000000
0!
0%
#295685000000
1!
1%
#295690000000
0!
0%
#295695000000
1!
1%
#295700000000
0!
0%
#295705000000
1!
1%
#295710000000
0!
0%
#295715000000
1!
1%
#295720000000
0!
0%
#295725000000
1!
1%
#295730000000
0!
0%
#295735000000
1!
1%
#295740000000
0!
0%
#295745000000
1!
1%
#295750000000
0!
0%
#295755000000
1!
1%
#295760000000
0!
0%
#295765000000
1!
1%
#295770000000
0!
0%
#295775000000
1!
1%
#295780000000
0!
0%
#295785000000
1!
1%
#295790000000
0!
0%
#295795000000
1!
1%
#295800000000
0!
0%
#295805000000
1!
1%
#295810000000
0!
0%
#295815000000
1!
1%
#295820000000
0!
0%
#295825000000
1!
1%
#295830000000
0!
0%
#295835000000
1!
1%
#295840000000
0!
0%
#295845000000
1!
1%
#295850000000
0!
0%
#295855000000
1!
1%
#295860000000
0!
0%
#295865000000
1!
1%
#295870000000
0!
0%
#295875000000
1!
1%
#295880000000
0!
0%
#295885000000
1!
1%
#295890000000
0!
0%
#295895000000
1!
1%
#295900000000
0!
0%
#295905000000
1!
1%
#295910000000
0!
0%
#295915000000
1!
1%
#295920000000
0!
0%
#295925000000
1!
1%
#295930000000
0!
0%
#295935000000
1!
1%
#295940000000
0!
0%
#295945000000
1!
1%
#295950000000
0!
0%
#295955000000
1!
1%
#295960000000
0!
0%
#295965000000
1!
1%
#295970000000
0!
0%
#295975000000
1!
1%
#295980000000
0!
0%
#295985000000
1!
1%
#295990000000
0!
0%
#295995000000
1!
1%
#296000000000
0!
0%
#296005000000
1!
1%
#296010000000
0!
0%
#296015000000
1!
1%
#296020000000
0!
0%
#296025000000
1!
1%
#296030000000
0!
0%
#296035000000
1!
1%
#296040000000
0!
0%
#296045000000
1!
1%
#296050000000
0!
0%
#296055000000
1!
1%
#296060000000
0!
0%
#296065000000
1!
1%
#296070000000
0!
0%
#296075000000
1!
1%
#296080000000
0!
0%
#296085000000
1!
1%
#296090000000
0!
0%
#296095000000
1!
1%
#296100000000
0!
0%
#296105000000
1!
1%
#296110000000
0!
0%
#296115000000
1!
1%
#296120000000
0!
0%
#296125000000
1!
1%
#296130000000
0!
0%
#296135000000
1!
1%
#296140000000
0!
0%
#296145000000
1!
1%
#296150000000
0!
0%
#296155000000
1!
1%
#296160000000
0!
0%
#296165000000
1!
1%
#296170000000
0!
0%
#296175000000
1!
1%
#296180000000
0!
0%
#296185000000
1!
1%
#296190000000
0!
0%
#296195000000
1!
1%
#296200000000
0!
0%
#296205000000
1!
1%
#296210000000
0!
0%
#296215000000
1!
1%
#296220000000
0!
0%
#296225000000
1!
1%
#296230000000
0!
0%
#296235000000
1!
1%
#296240000000
0!
0%
#296245000000
1!
1%
#296250000000
0!
0%
#296255000000
1!
1%
#296260000000
0!
0%
#296265000000
1!
1%
#296270000000
0!
0%
#296275000000
1!
1%
#296280000000
0!
0%
#296285000000
1!
1%
#296290000000
0!
0%
#296295000000
1!
1%
#296300000000
0!
0%
#296305000000
1!
1%
#296310000000
0!
0%
#296315000000
1!
1%
#296320000000
0!
0%
#296325000000
1!
1%
#296330000000
0!
0%
#296335000000
1!
1%
#296340000000
0!
0%
#296345000000
1!
1%
#296350000000
0!
0%
#296355000000
1!
1%
#296360000000
0!
0%
#296365000000
1!
1%
#296370000000
0!
0%
#296375000000
1!
1%
#296380000000
0!
0%
#296385000000
1!
1%
#296390000000
0!
0%
#296395000000
1!
1%
#296400000000
0!
0%
#296405000000
1!
1%
#296410000000
0!
0%
#296415000000
1!
1%
#296420000000
0!
0%
#296425000000
1!
1%
#296430000000
0!
0%
#296435000000
1!
1%
#296440000000
0!
0%
#296445000000
1!
1%
#296450000000
0!
0%
#296455000000
1!
1%
#296460000000
0!
0%
#296465000000
1!
1%
#296470000000
0!
0%
#296475000000
1!
1%
#296480000000
0!
0%
#296485000000
1!
1%
#296490000000
0!
0%
#296495000000
1!
1%
#296500000000
0!
0%
#296505000000
1!
1%
#296510000000
0!
0%
#296515000000
1!
1%
#296520000000
0!
0%
#296525000000
1!
1%
#296530000000
0!
0%
#296535000000
1!
1%
#296540000000
0!
0%
#296545000000
1!
1%
#296550000000
0!
0%
#296555000000
1!
1%
#296560000000
0!
0%
#296565000000
1!
1%
#296570000000
0!
0%
#296575000000
1!
1%
#296580000000
0!
0%
#296585000000
1!
1%
#296590000000
0!
0%
#296595000000
1!
1%
#296600000000
0!
0%
#296605000000
1!
1%
#296610000000
0!
0%
#296615000000
1!
1%
#296620000000
0!
0%
#296625000000
1!
1%
#296630000000
0!
0%
#296635000000
1!
1%
#296640000000
0!
0%
#296645000000
1!
1%
#296650000000
0!
0%
#296655000000
1!
1%
#296660000000
0!
0%
#296665000000
1!
1%
#296670000000
0!
0%
#296675000000
1!
1%
#296680000000
0!
0%
#296685000000
1!
1%
#296690000000
0!
0%
#296695000000
1!
1%
#296700000000
0!
0%
#296705000000
1!
1%
#296710000000
0!
0%
#296715000000
1!
1%
#296720000000
0!
0%
#296725000000
1!
1%
#296730000000
0!
0%
#296735000000
1!
1%
#296740000000
0!
0%
#296745000000
1!
1%
#296750000000
0!
0%
#296755000000
1!
1%
#296760000000
0!
0%
#296765000000
1!
1%
#296770000000
0!
0%
#296775000000
1!
1%
#296780000000
0!
0%
#296785000000
1!
1%
#296790000000
0!
0%
#296795000000
1!
1%
#296800000000
0!
0%
#296805000000
1!
1%
#296810000000
0!
0%
#296815000000
1!
1%
#296820000000
0!
0%
#296825000000
1!
1%
#296830000000
0!
0%
#296835000000
1!
1%
#296840000000
0!
0%
#296845000000
1!
1%
#296850000000
0!
0%
#296855000000
1!
1%
#296860000000
0!
0%
#296865000000
1!
1%
#296870000000
0!
0%
#296875000000
1!
1%
#296880000000
0!
0%
#296885000000
1!
1%
#296890000000
0!
0%
#296895000000
1!
1%
#296900000000
0!
0%
#296905000000
1!
1%
#296910000000
0!
0%
#296915000000
1!
1%
#296920000000
0!
0%
#296925000000
1!
1%
#296930000000
0!
0%
#296935000000
1!
1%
#296940000000
0!
0%
#296945000000
1!
1%
#296950000000
0!
0%
#296955000000
1!
1%
#296960000000
0!
0%
#296965000000
1!
1%
#296970000000
0!
0%
#296975000000
1!
1%
#296980000000
0!
0%
#296985000000
1!
1%
#296990000000
0!
0%
#296995000000
1!
1%
#297000000000
0!
0%
#297005000000
1!
1%
#297010000000
0!
0%
#297015000000
1!
1%
#297020000000
0!
0%
#297025000000
1!
1%
#297030000000
0!
0%
#297035000000
1!
1%
#297040000000
0!
0%
#297045000000
1!
1%
#297050000000
0!
0%
#297055000000
1!
1%
#297060000000
0!
0%
#297065000000
1!
1%
#297070000000
0!
0%
#297075000000
1!
1%
#297080000000
0!
0%
#297085000000
1!
1%
#297090000000
0!
0%
#297095000000
1!
1%
#297100000000
0!
0%
#297105000000
1!
1%
#297110000000
0!
0%
#297115000000
1!
1%
#297120000000
0!
0%
#297125000000
1!
1%
#297130000000
0!
0%
#297135000000
1!
1%
#297140000000
0!
0%
#297145000000
1!
1%
#297150000000
0!
0%
#297155000000
1!
1%
#297160000000
0!
0%
#297165000000
1!
1%
#297170000000
0!
0%
#297175000000
1!
1%
#297180000000
0!
0%
#297185000000
1!
1%
#297190000000
0!
0%
#297195000000
1!
1%
#297200000000
0!
0%
#297205000000
1!
1%
#297210000000
0!
0%
#297215000000
1!
1%
#297220000000
0!
0%
#297225000000
1!
1%
#297230000000
0!
0%
#297235000000
1!
1%
#297240000000
0!
0%
#297245000000
1!
1%
#297250000000
0!
0%
#297255000000
1!
1%
#297260000000
0!
0%
#297265000000
1!
1%
#297270000000
0!
0%
#297275000000
1!
1%
#297280000000
0!
0%
#297285000000
1!
1%
#297290000000
0!
0%
#297295000000
1!
1%
#297300000000
0!
0%
#297305000000
1!
1%
#297310000000
0!
0%
#297315000000
1!
1%
#297320000000
0!
0%
#297325000000
1!
1%
#297330000000
0!
0%
#297335000000
1!
1%
#297340000000
0!
0%
#297345000000
1!
1%
#297350000000
0!
0%
#297355000000
1!
1%
#297360000000
0!
0%
#297365000000
1!
1%
#297370000000
0!
0%
#297375000000
1!
1%
#297380000000
0!
0%
#297385000000
1!
1%
#297390000000
0!
0%
#297395000000
1!
1%
#297400000000
0!
0%
#297405000000
1!
1%
#297410000000
0!
0%
#297415000000
1!
1%
#297420000000
0!
0%
#297425000000
1!
1%
#297430000000
0!
0%
#297435000000
1!
1%
#297440000000
0!
0%
#297445000000
1!
1%
#297450000000
0!
0%
#297455000000
1!
1%
#297460000000
0!
0%
#297465000000
1!
1%
#297470000000
0!
0%
#297475000000
1!
1%
#297480000000
0!
0%
#297485000000
1!
1%
#297490000000
0!
0%
#297495000000
1!
1%
#297500000000
0!
0%
#297505000000
1!
1%
#297510000000
0!
0%
#297515000000
1!
1%
#297520000000
0!
0%
#297525000000
1!
1%
#297530000000
0!
0%
#297535000000
1!
1%
#297540000000
0!
0%
#297545000000
1!
1%
#297550000000
0!
0%
#297555000000
1!
1%
#297560000000
0!
0%
#297565000000
1!
1%
#297570000000
0!
0%
#297575000000
1!
1%
#297580000000
0!
0%
#297585000000
1!
1%
#297590000000
0!
0%
#297595000000
1!
1%
#297600000000
0!
0%
#297605000000
1!
1%
#297610000000
0!
0%
#297615000000
1!
1%
#297620000000
0!
0%
#297625000000
1!
1%
#297630000000
0!
0%
#297635000000
1!
1%
#297640000000
0!
0%
#297645000000
1!
1%
#297650000000
0!
0%
#297655000000
1!
1%
#297660000000
0!
0%
#297665000000
1!
1%
#297670000000
0!
0%
#297675000000
1!
1%
#297680000000
0!
0%
#297685000000
1!
1%
#297690000000
0!
0%
#297695000000
1!
1%
#297700000000
0!
0%
#297705000000
1!
1%
#297710000000
0!
0%
#297715000000
1!
1%
#297720000000
0!
0%
#297725000000
1!
1%
#297730000000
0!
0%
#297735000000
1!
1%
#297740000000
0!
0%
#297745000000
1!
1%
#297750000000
0!
0%
#297755000000
1!
1%
#297760000000
0!
0%
#297765000000
1!
1%
#297770000000
0!
0%
#297775000000
1!
1%
#297780000000
0!
0%
#297785000000
1!
1%
#297790000000
0!
0%
#297795000000
1!
1%
#297800000000
0!
0%
#297805000000
1!
1%
#297810000000
0!
0%
#297815000000
1!
1%
#297820000000
0!
0%
#297825000000
1!
1%
#297830000000
0!
0%
#297835000000
1!
1%
#297840000000
0!
0%
#297845000000
1!
1%
#297850000000
0!
0%
#297855000000
1!
1%
#297860000000
0!
0%
#297865000000
1!
1%
#297870000000
0!
0%
#297875000000
1!
1%
#297880000000
0!
0%
#297885000000
1!
1%
#297890000000
0!
0%
#297895000000
1!
1%
#297900000000
0!
0%
#297905000000
1!
1%
#297910000000
0!
0%
#297915000000
1!
1%
#297920000000
0!
0%
#297925000000
1!
1%
#297930000000
0!
0%
#297935000000
1!
1%
#297940000000
0!
0%
#297945000000
1!
1%
#297950000000
0!
0%
#297955000000
1!
1%
#297960000000
0!
0%
#297965000000
1!
1%
#297970000000
0!
0%
#297975000000
1!
1%
#297980000000
0!
0%
#297985000000
1!
1%
#297990000000
0!
0%
#297995000000
1!
1%
#298000000000
0!
0%
#298005000000
1!
1%
#298010000000
0!
0%
#298015000000
1!
1%
#298020000000
0!
0%
#298025000000
1!
1%
#298030000000
0!
0%
#298035000000
1!
1%
#298040000000
0!
0%
#298045000000
1!
1%
#298050000000
0!
0%
#298055000000
1!
1%
#298060000000
0!
0%
#298065000000
1!
1%
#298070000000
0!
0%
#298075000000
1!
1%
#298080000000
0!
0%
#298085000000
1!
1%
#298090000000
0!
0%
#298095000000
1!
1%
#298100000000
0!
0%
#298105000000
1!
1%
#298110000000
0!
0%
#298115000000
1!
1%
#298120000000
0!
0%
#298125000000
1!
1%
#298130000000
0!
0%
#298135000000
1!
1%
#298140000000
0!
0%
#298145000000
1!
1%
#298150000000
0!
0%
#298155000000
1!
1%
#298160000000
0!
0%
#298165000000
1!
1%
#298170000000
0!
0%
#298175000000
1!
1%
#298180000000
0!
0%
#298185000000
1!
1%
#298190000000
0!
0%
#298195000000
1!
1%
#298200000000
0!
0%
#298205000000
1!
1%
#298210000000
0!
0%
#298215000000
1!
1%
#298220000000
0!
0%
#298225000000
1!
1%
#298230000000
0!
0%
#298235000000
1!
1%
#298240000000
0!
0%
#298245000000
1!
1%
#298250000000
0!
0%
#298255000000
1!
1%
#298260000000
0!
0%
#298265000000
1!
1%
#298270000000
0!
0%
#298275000000
1!
1%
#298280000000
0!
0%
#298285000000
1!
1%
#298290000000
0!
0%
#298295000000
1!
1%
#298300000000
0!
0%
#298305000000
1!
1%
#298310000000
0!
0%
#298315000000
1!
1%
#298320000000
0!
0%
#298325000000
1!
1%
#298330000000
0!
0%
#298335000000
1!
1%
#298340000000
0!
0%
#298345000000
1!
1%
#298350000000
0!
0%
#298355000000
1!
1%
#298360000000
0!
0%
#298365000000
1!
1%
#298370000000
0!
0%
#298375000000
1!
1%
#298380000000
0!
0%
#298385000000
1!
1%
#298390000000
0!
0%
#298395000000
1!
1%
#298400000000
0!
0%
#298405000000
1!
1%
#298410000000
0!
0%
#298415000000
1!
1%
#298420000000
0!
0%
#298425000000
1!
1%
#298430000000
0!
0%
#298435000000
1!
1%
#298440000000
0!
0%
#298445000000
1!
1%
#298450000000
0!
0%
#298455000000
1!
1%
#298460000000
0!
0%
#298465000000
1!
1%
#298470000000
0!
0%
#298475000000
1!
1%
#298480000000
0!
0%
#298485000000
1!
1%
#298490000000
0!
0%
#298495000000
1!
1%
#298500000000
0!
0%
#298505000000
1!
1%
#298510000000
0!
0%
#298515000000
1!
1%
#298520000000
0!
0%
#298525000000
1!
1%
#298530000000
0!
0%
#298535000000
1!
1%
#298540000000
0!
0%
#298545000000
1!
1%
#298550000000
0!
0%
#298555000000
1!
1%
#298560000000
0!
0%
#298565000000
1!
1%
#298570000000
0!
0%
#298575000000
1!
1%
#298580000000
0!
0%
#298585000000
1!
1%
#298590000000
0!
0%
#298595000000
1!
1%
#298600000000
0!
0%
#298605000000
1!
1%
#298610000000
0!
0%
#298615000000
1!
1%
#298620000000
0!
0%
#298625000000
1!
1%
#298630000000
0!
0%
#298635000000
1!
1%
#298640000000
0!
0%
#298645000000
1!
1%
#298650000000
0!
0%
#298655000000
1!
1%
#298660000000
0!
0%
#298665000000
1!
1%
#298670000000
0!
0%
#298675000000
1!
1%
#298680000000
0!
0%
#298685000000
1!
1%
#298690000000
0!
0%
#298695000000
1!
1%
#298700000000
0!
0%
#298705000000
1!
1%
#298710000000
0!
0%
#298715000000
1!
1%
#298720000000
0!
0%
#298725000000
1!
1%
#298730000000
0!
0%
#298735000000
1!
1%
#298740000000
0!
0%
#298745000000
1!
1%
#298750000000
0!
0%
#298755000000
1!
1%
#298760000000
0!
0%
#298765000000
1!
1%
#298770000000
0!
0%
#298775000000
1!
1%
#298780000000
0!
0%
#298785000000
1!
1%
#298790000000
0!
0%
#298795000000
1!
1%
#298800000000
0!
0%
#298805000000
1!
1%
#298810000000
0!
0%
#298815000000
1!
1%
#298820000000
0!
0%
#298825000000
1!
1%
#298830000000
0!
0%
#298835000000
1!
1%
#298840000000
0!
0%
#298845000000
1!
1%
#298850000000
0!
0%
#298855000000
1!
1%
#298860000000
0!
0%
#298865000000
1!
1%
#298870000000
0!
0%
#298875000000
1!
1%
#298880000000
0!
0%
#298885000000
1!
1%
#298890000000
0!
0%
#298895000000
1!
1%
#298900000000
0!
0%
#298905000000
1!
1%
#298910000000
0!
0%
#298915000000
1!
1%
#298920000000
0!
0%
#298925000000
1!
1%
#298930000000
0!
0%
#298935000000
1!
1%
#298940000000
0!
0%
#298945000000
1!
1%
#298950000000
0!
0%
#298955000000
1!
1%
#298960000000
0!
0%
#298965000000
1!
1%
#298970000000
0!
0%
#298975000000
1!
1%
#298980000000
0!
0%
#298985000000
1!
1%
#298990000000
0!
0%
#298995000000
1!
1%
#299000000000
0!
0%
#299005000000
1!
1%
#299010000000
0!
0%
#299015000000
1!
1%
#299020000000
0!
0%
#299025000000
1!
1%
#299030000000
0!
0%
#299035000000
1!
1%
#299040000000
0!
0%
#299045000000
1!
1%
#299050000000
0!
0%
#299055000000
1!
1%
#299060000000
0!
0%
#299065000000
1!
1%
#299070000000
0!
0%
#299075000000
1!
1%
#299080000000
0!
0%
#299085000000
1!
1%
#299090000000
0!
0%
#299095000000
1!
1%
#299100000000
0!
0%
#299105000000
1!
1%
#299110000000
0!
0%
#299115000000
1!
1%
#299120000000
0!
0%
#299125000000
1!
1%
#299130000000
0!
0%
#299135000000
1!
1%
#299140000000
0!
0%
#299145000000
1!
1%
#299150000000
0!
0%
#299155000000
1!
1%
#299160000000
0!
0%
#299165000000
1!
1%
#299170000000
0!
0%
#299175000000
1!
1%
#299180000000
0!
0%
#299185000000
1!
1%
#299190000000
0!
0%
#299195000000
1!
1%
#299200000000
0!
0%
#299205000000
1!
1%
#299210000000
0!
0%
#299215000000
1!
1%
#299220000000
0!
0%
#299225000000
1!
1%
#299230000000
0!
0%
#299235000000
1!
1%
#299240000000
0!
0%
#299245000000
1!
1%
#299250000000
0!
0%
#299255000000
1!
1%
#299260000000
0!
0%
#299265000000
1!
1%
#299270000000
0!
0%
#299275000000
1!
1%
#299280000000
0!
0%
#299285000000
1!
1%
#299290000000
0!
0%
#299295000000
1!
1%
#299300000000
0!
0%
#299305000000
1!
1%
#299310000000
0!
0%
#299315000000
1!
1%
#299320000000
0!
0%
#299325000000
1!
1%
#299330000000
0!
0%
#299335000000
1!
1%
#299340000000
0!
0%
#299345000000
1!
1%
#299350000000
0!
0%
#299355000000
1!
1%
#299360000000
0!
0%
#299365000000
1!
1%
#299370000000
0!
0%
#299375000000
1!
1%
#299380000000
0!
0%
#299385000000
1!
1%
#299390000000
0!
0%
#299395000000
1!
1%
#299400000000
0!
0%
#299405000000
1!
1%
#299410000000
0!
0%
#299415000000
1!
1%
#299420000000
0!
0%
#299425000000
1!
1%
#299430000000
0!
0%
#299435000000
1!
1%
#299440000000
0!
0%
#299445000000
1!
1%
#299450000000
0!
0%
#299455000000
1!
1%
#299460000000
0!
0%
#299465000000
1!
1%
#299470000000
0!
0%
#299475000000
1!
1%
#299480000000
0!
0%
#299485000000
1!
1%
#299490000000
0!
0%
#299495000000
1!
1%
#299500000000
0!
0%
#299505000000
1!
1%
#299510000000
0!
0%
#299515000000
1!
1%
#299520000000
0!
0%
#299525000000
1!
1%
#299530000000
0!
0%
#299535000000
1!
1%
#299540000000
0!
0%
#299545000000
1!
1%
#299550000000
0!
0%
#299555000000
1!
1%
#299560000000
0!
0%
#299565000000
1!
1%
#299570000000
0!
0%
#299575000000
1!
1%
#299580000000
0!
0%
#299585000000
1!
1%
#299590000000
0!
0%
#299595000000
1!
1%
#299600000000
0!
0%
#299605000000
1!
1%
#299610000000
0!
0%
#299615000000
1!
1%
#299620000000
0!
0%
#299625000000
1!
1%
#299630000000
0!
0%
#299635000000
1!
1%
#299640000000
0!
0%
#299645000000
1!
1%
#299650000000
0!
0%
#299655000000
1!
1%
#299660000000
0!
0%
#299665000000
1!
1%
#299670000000
0!
0%
#299675000000
1!
1%
#299680000000
0!
0%
#299685000000
1!
1%
#299690000000
0!
0%
#299695000000
1!
1%
#299700000000
0!
0%
#299705000000
1!
1%
#299710000000
0!
0%
#299715000000
1!
1%
#299720000000
0!
0%
#299725000000
1!
1%
#299730000000
0!
0%
#299735000000
1!
1%
#299740000000
0!
0%
#299745000000
1!
1%
#299750000000
0!
0%
#299755000000
1!
1%
#299760000000
0!
0%
#299765000000
1!
1%
#299770000000
0!
0%
#299775000000
1!
1%
#299780000000
0!
0%
#299785000000
1!
1%
#299790000000
0!
0%
#299795000000
1!
1%
#299800000000
0!
0%
#299805000000
1!
1%
#299810000000
0!
0%
#299815000000
1!
1%
#299820000000
0!
0%
#299825000000
1!
1%
#299830000000
0!
0%
#299835000000
1!
1%
#299840000000
0!
0%
#299845000000
1!
1%
#299850000000
0!
0%
#299855000000
1!
1%
#299860000000
0!
0%
#299865000000
1!
1%
#299870000000
0!
0%
#299875000000
1!
1%
#299880000000
0!
0%
#299885000000
1!
1%
#299890000000
0!
0%
#299895000000
1!
1%
#299900000000
0!
0%
#299905000000
1!
1%
#299910000000
0!
0%
#299915000000
1!
1%
#299920000000
0!
0%
#299925000000
1!
1%
#299930000000
0!
0%
#299935000000
1!
1%
#299940000000
0!
0%
#299945000000
1!
1%
#299950000000
0!
0%
#299955000000
1!
1%
#299960000000
0!
0%
#299965000000
1!
1%
#299970000000
0!
0%
#299975000000
1!
1%
#299980000000
0!
0%
#299985000000
1!
1%
#299990000000
0!
0%
#299995000000
1!
1%
#300000000000
0!
0%
#300005000000
1!
1%
#300010000000
0!
0%
#300015000000
1!
1%
#300020000000
0!
0%
#300025000000
1!
1%
#300030000000
0!
0%
#300035000000
1!
1%
#300040000000
0!
0%
#300045000000
1!
1%
#300050000000
0!
0%
#300055000000
1!
1%
#300060000000
0!
0%
#300065000000
1!
1%
#300070000000
0!
0%
#300075000000
1!
1%
#300080000000
0!
0%
#300085000000
1!
1%
#300090000000
0!
0%
#300095000000
1!
1%
#300100000000
0!
0%
#300105000000
1!
1%
#300110000000
0!
0%
#300115000000
1!
1%
#300120000000
0!
0%
#300125000000
1!
1%
#300130000000
0!
0%
#300135000000
1!
1%
#300140000000
0!
0%
#300145000000
1!
1%
#300150000000
0!
0%
#300155000000
1!
1%
#300160000000
0!
0%
#300165000000
1!
1%
#300170000000
0!
0%
#300175000000
1!
1%
#300180000000
0!
0%
#300185000000
1!
1%
#300190000000
0!
0%
#300195000000
1!
1%
#300200000000
0!
0%
#300205000000
1!
1%
#300210000000
0!
0%
#300215000000
1!
1%
#300220000000
0!
0%
#300225000000
1!
1%
#300230000000
0!
0%
#300235000000
1!
1%
#300240000000
0!
0%
#300245000000
1!
1%
#300250000000
0!
0%
#300255000000
1!
1%
#300260000000
0!
0%
#300265000000
1!
1%
#300270000000
0!
0%
#300275000000
1!
1%
#300280000000
0!
0%
#300285000000
1!
1%
#300290000000
0!
0%
#300295000000
1!
1%
#300300000000
0!
0%
#300305000000
1!
1%
#300310000000
0!
0%
#300315000000
1!
1%
#300320000000
0!
0%
#300325000000
1!
1%
#300330000000
0!
0%
#300335000000
1!
1%
#300340000000
0!
0%
#300345000000
1!
1%
#300350000000
0!
0%
#300355000000
1!
1%
#300360000000
0!
0%
#300365000000
1!
1%
#300370000000
0!
0%
#300375000000
1!
1%
#300380000000
0!
0%
#300385000000
1!
1%
#300390000000
0!
0%
#300395000000
1!
1%
#300400000000
0!
0%
#300405000000
1!
1%
#300410000000
0!
0%
#300415000000
1!
1%
#300420000000
0!
0%
#300425000000
1!
1%
#300430000000
0!
0%
#300435000000
1!
1%
#300440000000
0!
0%
#300445000000
1!
1%
#300450000000
0!
0%
#300455000000
1!
1%
#300460000000
0!
0%
#300465000000
1!
1%
#300470000000
0!
0%
#300475000000
1!
1%
#300480000000
0!
0%
#300485000000
1!
1%
#300490000000
0!
0%
#300495000000
1!
1%
#300500000000
0!
0%
#300505000000
1!
1%
#300510000000
0!
0%
#300515000000
1!
1%
#300520000000
0!
0%
#300525000000
1!
1%
#300530000000
0!
0%
#300535000000
1!
1%
#300540000000
0!
0%
#300545000000
1!
1%
#300550000000
0!
0%
#300555000000
1!
1%
#300560000000
0!
0%
#300565000000
1!
1%
#300570000000
0!
0%
#300575000000
1!
1%
#300580000000
0!
0%
#300585000000
1!
1%
#300590000000
0!
0%
#300595000000
1!
1%
#300600000000
0!
0%
#300605000000
1!
1%
#300610000000
0!
0%
#300615000000
1!
1%
#300620000000
0!
0%
#300625000000
1!
1%
#300630000000
0!
0%
#300635000000
1!
1%
#300640000000
0!
0%
#300645000000
1!
1%
#300650000000
0!
0%
#300655000000
1!
1%
#300660000000
0!
0%
#300665000000
1!
1%
#300670000000
0!
0%
#300675000000
1!
1%
#300680000000
0!
0%
#300685000000
1!
1%
#300690000000
0!
0%
#300695000000
1!
1%
#300700000000
0!
0%
#300705000000
1!
1%
#300710000000
0!
0%
#300715000000
1!
1%
#300720000000
0!
0%
#300725000000
1!
1%
#300730000000
0!
0%
#300735000000
1!
1%
#300740000000
0!
0%
#300745000000
1!
1%
#300750000000
0!
0%
#300755000000
1!
1%
#300760000000
0!
0%
#300765000000
1!
1%
#300770000000
0!
0%
#300775000000
1!
1%
#300780000000
0!
0%
#300785000000
1!
1%
#300790000000
0!
0%
#300795000000
1!
1%
#300800000000
0!
0%
#300805000000
1!
1%
#300810000000
0!
0%
#300815000000
1!
1%
#300820000000
0!
0%
#300825000000
1!
1%
#300830000000
0!
0%
#300835000000
1!
1%
#300840000000
0!
0%
#300845000000
1!
1%
#300850000000
0!
0%
#300855000000
1!
1%
#300860000000
0!
0%
#300865000000
1!
1%
#300870000000
0!
0%
#300875000000
1!
1%
#300880000000
0!
0%
#300885000000
1!
1%
#300890000000
0!
0%
#300895000000
1!
1%
#300900000000
0!
0%
#300905000000
1!
1%
#300910000000
0!
0%
#300915000000
1!
1%
#300920000000
0!
0%
#300925000000
1!
1%
#300930000000
0!
0%
#300935000000
1!
1%
#300940000000
0!
0%
#300945000000
1!
1%
#300950000000
0!
0%
#300955000000
1!
1%
#300960000000
0!
0%
#300965000000
1!
1%
#300970000000
0!
0%
#300975000000
1!
1%
#300980000000
0!
0%
#300985000000
1!
1%
#300990000000
0!
0%
#300995000000
1!
1%
#301000000000
0!
0%
#301005000000
1!
1%
#301010000000
0!
0%
#301015000000
1!
1%
#301020000000
0!
0%
#301025000000
1!
1%
#301030000000
0!
0%
#301035000000
1!
1%
#301040000000
0!
0%
#301045000000
1!
1%
#301050000000
0!
0%
#301055000000
1!
1%
#301060000000
0!
0%
#301065000000
1!
1%
#301070000000
0!
0%
#301075000000
1!
1%
#301080000000
0!
0%
#301085000000
1!
1%
#301090000000
0!
0%
#301095000000
1!
1%
#301100000000
0!
0%
#301105000000
1!
1%
#301110000000
0!
0%
#301115000000
1!
1%
#301120000000
0!
0%
#301125000000
1!
1%
#301130000000
0!
0%
#301135000000
1!
1%
#301140000000
0!
0%
#301145000000
1!
1%
#301150000000
0!
0%
#301155000000
1!
1%
#301160000000
0!
0%
#301165000000
1!
1%
#301170000000
0!
0%
#301175000000
1!
1%
#301180000000
0!
0%
#301185000000
1!
1%
#301190000000
0!
0%
#301195000000
1!
1%
#301200000000
0!
0%
#301205000000
1!
1%
#301210000000
0!
0%
#301215000000
1!
1%
#301220000000
0!
0%
#301225000000
1!
1%
#301230000000
0!
0%
#301235000000
1!
1%
#301240000000
0!
0%
#301245000000
1!
1%
#301250000000
0!
0%
#301255000000
1!
1%
#301260000000
0!
0%
#301265000000
1!
1%
#301270000000
0!
0%
#301275000000
1!
1%
#301280000000
0!
0%
#301285000000
1!
1%
#301290000000
0!
0%
#301295000000
1!
1%
#301300000000
0!
0%
#301305000000
1!
1%
#301310000000
0!
0%
#301315000000
1!
1%
#301320000000
0!
0%
#301325000000
1!
1%
#301330000000
0!
0%
#301335000000
1!
1%
#301340000000
0!
0%
#301345000000
1!
1%
#301350000000
0!
0%
#301355000000
1!
1%
#301360000000
0!
0%
#301365000000
1!
1%
#301370000000
0!
0%
#301375000000
1!
1%
#301380000000
0!
0%
#301385000000
1!
1%
#301390000000
0!
0%
#301395000000
1!
1%
#301400000000
0!
0%
#301405000000
1!
1%
#301410000000
0!
0%
#301415000000
1!
1%
#301420000000
0!
0%
#301425000000
1!
1%
#301430000000
0!
0%
#301435000000
1!
1%
#301440000000
0!
0%
#301445000000
1!
1%
#301450000000
0!
0%
#301455000000
1!
1%
#301460000000
0!
0%
#301465000000
1!
1%
#301470000000
0!
0%
#301475000000
1!
1%
#301480000000
0!
0%
#301485000000
1!
1%
#301490000000
0!
0%
#301495000000
1!
1%
#301500000000
0!
0%
#301505000000
1!
1%
#301510000000
0!
0%
#301515000000
1!
1%
#301520000000
0!
0%
#301525000000
1!
1%
#301530000000
0!
0%
#301535000000
1!
1%
#301540000000
0!
0%
#301545000000
1!
1%
#301550000000
0!
0%
#301555000000
1!
1%
#301560000000
0!
0%
#301565000000
1!
1%
#301570000000
0!
0%
#301575000000
1!
1%
#301580000000
0!
0%
#301585000000
1!
1%
#301590000000
0!
0%
#301595000000
1!
1%
#301600000000
0!
0%
#301605000000
1!
1%
#301610000000
0!
0%
#301615000000
1!
1%
#301620000000
0!
0%
#301625000000
1!
1%
#301630000000
0!
0%
#301635000000
1!
1%
#301640000000
0!
0%
#301645000000
1!
1%
#301650000000
0!
0%
#301655000000
1!
1%
#301660000000
0!
0%
#301665000000
1!
1%
#301670000000
0!
0%
#301675000000
1!
1%
#301680000000
0!
0%
#301685000000
1!
1%
#301690000000
0!
0%
#301695000000
1!
1%
#301700000000
0!
0%
#301705000000
1!
1%
#301710000000
0!
0%
#301715000000
1!
1%
#301720000000
0!
0%
#301725000000
1!
1%
#301730000000
0!
0%
#301735000000
1!
1%
#301740000000
0!
0%
#301745000000
1!
1%
#301750000000
0!
0%
#301755000000
1!
1%
#301760000000
0!
0%
#301765000000
1!
1%
#301770000000
0!
0%
#301775000000
1!
1%
#301780000000
0!
0%
#301785000000
1!
1%
#301790000000
0!
0%
#301795000000
1!
1%
#301800000000
0!
0%
#301805000000
1!
1%
#301810000000
0!
0%
#301815000000
1!
1%
#301820000000
0!
0%
#301825000000
1!
1%
#301830000000
0!
0%
#301835000000
1!
1%
#301840000000
0!
0%
#301845000000
1!
1%
#301850000000
0!
0%
#301855000000
1!
1%
#301860000000
0!
0%
#301865000000
1!
1%
#301870000000
0!
0%
#301875000000
1!
1%
#301880000000
0!
0%
#301885000000
1!
1%
#301890000000
0!
0%
#301895000000
1!
1%
#301900000000
0!
0%
#301905000000
1!
1%
#301910000000
0!
0%
#301915000000
1!
1%
#301920000000
0!
0%
#301925000000
1!
1%
#301930000000
0!
0%
#301935000000
1!
1%
#301940000000
0!
0%
#301945000000
1!
1%
#301950000000
0!
0%
#301955000000
1!
1%
#301960000000
0!
0%
#301965000000
1!
1%
#301970000000
0!
0%
#301975000000
1!
1%
#301980000000
0!
0%
#301985000000
1!
1%
#301990000000
0!
0%
#301995000000
1!
1%
#302000000000
0!
0%
#302005000000
1!
1%
#302010000000
0!
0%
#302015000000
1!
1%
#302020000000
0!
0%
#302025000000
1!
1%
#302030000000
0!
0%
#302035000000
1!
1%
#302040000000
0!
0%
#302045000000
1!
1%
#302050000000
0!
0%
#302055000000
1!
1%
#302060000000
0!
0%
#302065000000
1!
1%
#302070000000
0!
0%
#302075000000
1!
1%
#302080000000
0!
0%
#302085000000
1!
1%
#302090000000
0!
0%
#302095000000
1!
1%
#302100000000
0!
0%
#302105000000
1!
1%
#302110000000
0!
0%
#302115000000
1!
1%
#302120000000
0!
0%
#302125000000
1!
1%
#302130000000
0!
0%
#302135000000
1!
1%
#302140000000
0!
0%
#302145000000
1!
1%
#302150000000
0!
0%
#302155000000
1!
1%
#302160000000
0!
0%
#302165000000
1!
1%
#302170000000
0!
0%
#302175000000
1!
1%
#302180000000
0!
0%
#302185000000
1!
1%
#302190000000
0!
0%
#302195000000
1!
1%
#302200000000
0!
0%
#302205000000
1!
1%
#302210000000
0!
0%
#302215000000
1!
1%
#302220000000
0!
0%
#302225000000
1!
1%
#302230000000
0!
0%
#302235000000
1!
1%
#302240000000
0!
0%
#302245000000
1!
1%
#302250000000
0!
0%
#302255000000
1!
1%
#302260000000
0!
0%
#302265000000
1!
1%
#302270000000
0!
0%
#302275000000
1!
1%
#302280000000
0!
0%
#302285000000
1!
1%
#302290000000
0!
0%
#302295000000
1!
1%
#302300000000
0!
0%
#302305000000
1!
1%
#302310000000
0!
0%
#302315000000
1!
1%
#302320000000
0!
0%
#302325000000
1!
1%
#302330000000
0!
0%
#302335000000
1!
1%
#302340000000
0!
0%
#302345000000
1!
1%
#302350000000
0!
0%
#302355000000
1!
1%
#302360000000
0!
0%
#302365000000
1!
1%
#302370000000
0!
0%
#302375000000
1!
1%
#302380000000
0!
0%
#302385000000
1!
1%
#302390000000
0!
0%
#302395000000
1!
1%
#302400000000
0!
0%
#302405000000
1!
1%
#302410000000
0!
0%
#302415000000
1!
1%
#302420000000
0!
0%
#302425000000
1!
1%
#302430000000
0!
0%
#302435000000
1!
1%
#302440000000
0!
0%
#302445000000
1!
1%
#302450000000
0!
0%
#302455000000
1!
1%
#302460000000
0!
0%
#302465000000
1!
1%
#302470000000
0!
0%
#302475000000
1!
1%
#302480000000
0!
0%
#302485000000
1!
1%
#302490000000
0!
0%
#302495000000
1!
1%
#302500000000
0!
0%
#302505000000
1!
1%
#302510000000
0!
0%
#302515000000
1!
1%
#302520000000
0!
0%
#302525000000
1!
1%
#302530000000
0!
0%
#302535000000
1!
1%
#302540000000
0!
0%
#302545000000
1!
1%
#302550000000
0!
0%
#302555000000
1!
1%
#302560000000
0!
0%
#302565000000
1!
1%
#302570000000
0!
0%
#302575000000
1!
1%
#302580000000
0!
0%
#302585000000
1!
1%
#302590000000
0!
0%
#302595000000
1!
1%
#302600000000
0!
0%
#302605000000
1!
1%
#302610000000
0!
0%
#302615000000
1!
1%
#302620000000
0!
0%
#302625000000
1!
1%
#302630000000
0!
0%
#302635000000
1!
1%
#302640000000
0!
0%
#302645000000
1!
1%
#302650000000
0!
0%
#302655000000
1!
1%
#302660000000
0!
0%
#302665000000
1!
1%
#302670000000
0!
0%
#302675000000
1!
1%
#302680000000
0!
0%
#302685000000
1!
1%
#302690000000
0!
0%
#302695000000
1!
1%
#302700000000
0!
0%
#302705000000
1!
1%
#302710000000
0!
0%
#302715000000
1!
1%
#302720000000
0!
0%
#302725000000
1!
1%
#302730000000
0!
0%
#302735000000
1!
1%
#302740000000
0!
0%
#302745000000
1!
1%
#302750000000
0!
0%
#302755000000
1!
1%
#302760000000
0!
0%
#302765000000
1!
1%
#302770000000
0!
0%
#302775000000
1!
1%
#302780000000
0!
0%
#302785000000
1!
1%
#302790000000
0!
0%
#302795000000
1!
1%
#302800000000
0!
0%
#302805000000
1!
1%
#302810000000
0!
0%
#302815000000
1!
1%
#302820000000
0!
0%
#302825000000
1!
1%
#302830000000
0!
0%
#302835000000
1!
1%
#302840000000
0!
0%
#302845000000
1!
1%
#302850000000
0!
0%
#302855000000
1!
1%
#302860000000
0!
0%
#302865000000
1!
1%
#302870000000
0!
0%
#302875000000
1!
1%
#302880000000
0!
0%
#302885000000
1!
1%
#302890000000
0!
0%
#302895000000
1!
1%
#302900000000
0!
0%
#302905000000
1!
1%
#302910000000
0!
0%
#302915000000
1!
1%
#302920000000
0!
0%
#302925000000
1!
1%
#302930000000
0!
0%
#302935000000
1!
1%
#302940000000
0!
0%
#302945000000
1!
1%
#302950000000
0!
0%
#302955000000
1!
1%
#302960000000
0!
0%
#302965000000
1!
1%
#302970000000
0!
0%
#302975000000
1!
1%
#302980000000
0!
0%
#302985000000
1!
1%
#302990000000
0!
0%
#302995000000
1!
1%
#303000000000
0!
0%
#303005000000
1!
1%
#303010000000
0!
0%
#303015000000
1!
1%
#303020000000
0!
0%
#303025000000
1!
1%
#303030000000
0!
0%
#303035000000
1!
1%
#303040000000
0!
0%
#303045000000
1!
1%
#303050000000
0!
0%
#303055000000
1!
1%
#303060000000
0!
0%
#303065000000
1!
1%
#303070000000
0!
0%
#303075000000
1!
1%
#303080000000
0!
0%
#303085000000
1!
1%
#303090000000
0!
0%
#303095000000
1!
1%
#303100000000
0!
0%
#303105000000
1!
1%
#303110000000
0!
0%
#303115000000
1!
1%
#303120000000
0!
0%
#303125000000
1!
1%
#303130000000
0!
0%
#303135000000
1!
1%
#303140000000
0!
0%
#303145000000
1!
1%
#303150000000
0!
0%
#303155000000
1!
1%
#303160000000
0!
0%
#303165000000
1!
1%
#303170000000
0!
0%
#303175000000
1!
1%
#303180000000
0!
0%
#303185000000
1!
1%
#303190000000
0!
0%
#303195000000
1!
1%
#303200000000
0!
0%
#303205000000
1!
1%
#303210000000
0!
0%
#303215000000
1!
1%
#303220000000
0!
0%
#303225000000
1!
1%
#303230000000
0!
0%
#303235000000
1!
1%
#303240000000
0!
0%
#303245000000
1!
1%
#303250000000
0!
0%
#303255000000
1!
1%
#303260000000
0!
0%
#303265000000
1!
1%
#303270000000
0!
0%
#303275000000
1!
1%
#303280000000
0!
0%
#303285000000
1!
1%
#303290000000
0!
0%
#303295000000
1!
1%
#303300000000
0!
0%
#303305000000
1!
1%
#303310000000
0!
0%
#303315000000
1!
1%
#303320000000
0!
0%
#303325000000
1!
1%
#303330000000
0!
0%
#303335000000
1!
1%
#303340000000
0!
0%
#303345000000
1!
1%
#303350000000
0!
0%
#303355000000
1!
1%
#303360000000
0!
0%
#303365000000
1!
1%
#303370000000
0!
0%
#303375000000
1!
1%
#303380000000
0!
0%
#303385000000
1!
1%
#303390000000
0!
0%
#303395000000
1!
1%
#303400000000
0!
0%
#303405000000
1!
1%
#303410000000
0!
0%
#303415000000
1!
1%
#303420000000
0!
0%
#303425000000
1!
1%
#303430000000
0!
0%
#303435000000
1!
1%
#303440000000
0!
0%
#303445000000
1!
1%
#303450000000
0!
0%
#303455000000
1!
1%
#303460000000
0!
0%
#303465000000
1!
1%
#303470000000
0!
0%
#303475000000
1!
1%
#303480000000
0!
0%
#303485000000
1!
1%
#303490000000
0!
0%
#303495000000
1!
1%
#303500000000
0!
0%
#303505000000
1!
1%
#303510000000
0!
0%
#303515000000
1!
1%
#303520000000
0!
0%
#303525000000
1!
1%
#303530000000
0!
0%
#303535000000
1!
1%
#303540000000
0!
0%
#303545000000
1!
1%
#303550000000
0!
0%
#303555000000
1!
1%
#303560000000
0!
0%
#303565000000
1!
1%
#303570000000
0!
0%
#303575000000
1!
1%
#303580000000
0!
0%
#303585000000
1!
1%
#303590000000
0!
0%
#303595000000
1!
1%
#303600000000
0!
0%
#303605000000
1!
1%
#303610000000
0!
0%
#303615000000
1!
1%
#303620000000
0!
0%
#303625000000
1!
1%
#303630000000
0!
0%
#303635000000
1!
1%
#303640000000
0!
0%
#303645000000
1!
1%
#303650000000
0!
0%
#303655000000
1!
1%
#303660000000
0!
0%
#303665000000
1!
1%
#303670000000
0!
0%
#303675000000
1!
1%
#303680000000
0!
0%
#303685000000
1!
1%
#303690000000
0!
0%
#303695000000
1!
1%
#303700000000
0!
0%
#303705000000
1!
1%
#303710000000
0!
0%
#303715000000
1!
1%
#303720000000
0!
0%
#303725000000
1!
1%
#303730000000
0!
0%
#303735000000
1!
1%
#303740000000
0!
0%
#303745000000
1!
1%
#303750000000
0!
0%
#303755000000
1!
1%
#303760000000
0!
0%
#303765000000
1!
1%
#303770000000
0!
0%
#303775000000
1!
1%
#303780000000
0!
0%
#303785000000
1!
1%
#303790000000
0!
0%
#303795000000
1!
1%
#303800000000
0!
0%
#303805000000
1!
1%
#303810000000
0!
0%
#303815000000
1!
1%
#303820000000
0!
0%
#303825000000
1!
1%
#303830000000
0!
0%
#303835000000
1!
1%
#303840000000
0!
0%
#303845000000
1!
1%
#303850000000
0!
0%
#303855000000
1!
1%
#303860000000
0!
0%
#303865000000
1!
1%
#303870000000
0!
0%
#303875000000
1!
1%
#303880000000
0!
0%
#303885000000
1!
1%
#303890000000
0!
0%
#303895000000
1!
1%
#303900000000
0!
0%
#303905000000
1!
1%
#303910000000
0!
0%
#303915000000
1!
1%
#303920000000
0!
0%
#303925000000
1!
1%
#303930000000
0!
0%
#303935000000
1!
1%
#303940000000
0!
0%
#303945000000
1!
1%
#303950000000
0!
0%
#303955000000
1!
1%
#303960000000
0!
0%
#303965000000
1!
1%
#303970000000
0!
0%
#303975000000
1!
1%
#303980000000
0!
0%
#303985000000
1!
1%
#303990000000
0!
0%
#303995000000
1!
1%
#304000000000
0!
0%
#304005000000
1!
1%
#304010000000
0!
0%
#304015000000
1!
1%
#304020000000
0!
0%
#304025000000
1!
1%
#304030000000
0!
0%
#304035000000
1!
1%
#304040000000
0!
0%
#304045000000
1!
1%
#304050000000
0!
0%
#304055000000
1!
1%
#304060000000
0!
0%
#304065000000
1!
1%
#304070000000
0!
0%
#304075000000
1!
1%
#304080000000
0!
0%
#304085000000
1!
1%
#304090000000
0!
0%
#304095000000
1!
1%
#304100000000
0!
0%
#304105000000
1!
1%
#304110000000
0!
0%
#304115000000
1!
1%
#304120000000
0!
0%
#304125000000
1!
1%
#304130000000
0!
0%
#304135000000
1!
1%
#304140000000
0!
0%
#304145000000
1!
1%
#304150000000
0!
0%
#304155000000
1!
1%
#304160000000
0!
0%
#304165000000
1!
1%
#304170000000
0!
0%
#304175000000
1!
1%
#304180000000
0!
0%
#304185000000
1!
1%
#304190000000
0!
0%
#304195000000
1!
1%
#304200000000
0!
0%
#304205000000
1!
1%
#304210000000
0!
0%
#304215000000
1!
1%
#304220000000
0!
0%
#304225000000
1!
1%
#304230000000
0!
0%
#304235000000
1!
1%
#304240000000
0!
0%
#304245000000
1!
1%
#304250000000
0!
0%
#304255000000
1!
1%
#304260000000
0!
0%
#304265000000
1!
1%
#304270000000
0!
0%
#304275000000
1!
1%
#304280000000
0!
0%
#304285000000
1!
1%
#304290000000
0!
0%
#304295000000
1!
1%
#304300000000
0!
0%
#304305000000
1!
1%
#304310000000
0!
0%
#304315000000
1!
1%
#304320000000
0!
0%
#304325000000
1!
1%
#304330000000
0!
0%
#304335000000
1!
1%
#304340000000
0!
0%
#304345000000
1!
1%
#304350000000
0!
0%
#304355000000
1!
1%
#304360000000
0!
0%
#304365000000
1!
1%
#304370000000
0!
0%
#304375000000
1!
1%
#304380000000
0!
0%
#304385000000
1!
1%
#304390000000
0!
0%
#304395000000
1!
1%
#304400000000
0!
0%
#304405000000
1!
1%
#304410000000
0!
0%
#304415000000
1!
1%
#304420000000
0!
0%
#304425000000
1!
1%
#304430000000
0!
0%
#304435000000
1!
1%
#304440000000
0!
0%
#304445000000
1!
1%
#304450000000
0!
0%
#304455000000
1!
1%
#304460000000
0!
0%
#304465000000
1!
1%
#304470000000
0!
0%
#304475000000
1!
1%
#304480000000
0!
0%
#304485000000
1!
1%
#304490000000
0!
0%
#304495000000
1!
1%
#304500000000
0!
0%
#304505000000
1!
1%
#304510000000
0!
0%
#304515000000
1!
1%
#304520000000
0!
0%
#304525000000
1!
1%
#304530000000
0!
0%
#304535000000
1!
1%
#304540000000
0!
0%
#304545000000
1!
1%
#304550000000
0!
0%
#304555000000
1!
1%
#304560000000
0!
0%
#304565000000
1!
1%
#304570000000
0!
0%
#304575000000
1!
1%
#304580000000
0!
0%
#304585000000
1!
1%
#304590000000
0!
0%
#304595000000
1!
1%
#304600000000
0!
0%
#304605000000
1!
1%
#304610000000
0!
0%
#304615000000
1!
1%
#304620000000
0!
0%
#304625000000
1!
1%
#304630000000
0!
0%
#304635000000
1!
1%
#304640000000
0!
0%
#304645000000
1!
1%
#304650000000
0!
0%
#304655000000
1!
1%
#304660000000
0!
0%
#304665000000
1!
1%
#304670000000
0!
0%
#304675000000
1!
1%
#304680000000
0!
0%
#304685000000
1!
1%
#304690000000
0!
0%
#304695000000
1!
1%
#304700000000
0!
0%
#304705000000
1!
1%
#304710000000
0!
0%
#304715000000
1!
1%
#304720000000
0!
0%
#304725000000
1!
1%
#304730000000
0!
0%
#304735000000
1!
1%
#304740000000
0!
0%
#304745000000
1!
1%
#304750000000
0!
0%
#304755000000
1!
1%
#304760000000
0!
0%
#304765000000
1!
1%
#304770000000
0!
0%
#304775000000
1!
1%
#304780000000
0!
0%
#304785000000
1!
1%
#304790000000
0!
0%
#304795000000
1!
1%
#304800000000
0!
0%
#304805000000
1!
1%
#304810000000
0!
0%
#304815000000
1!
1%
#304820000000
0!
0%
#304825000000
1!
1%
#304830000000
0!
0%
#304835000000
1!
1%
#304840000000
0!
0%
#304845000000
1!
1%
#304850000000
0!
0%
#304855000000
1!
1%
#304860000000
0!
0%
#304865000000
1!
1%
#304870000000
0!
0%
#304875000000
1!
1%
#304880000000
0!
0%
#304885000000
1!
1%
#304890000000
0!
0%
#304895000000
1!
1%
#304900000000
0!
0%
#304905000000
1!
1%
#304910000000
0!
0%
#304915000000
1!
1%
#304920000000
0!
0%
#304925000000
1!
1%
#304930000000
0!
0%
#304935000000
1!
1%
#304940000000
0!
0%
#304945000000
1!
1%
#304950000000
0!
0%
#304955000000
1!
1%
#304960000000
0!
0%
#304965000000
1!
1%
#304970000000
0!
0%
#304975000000
1!
1%
#304980000000
0!
0%
#304985000000
1!
1%
#304990000000
0!
0%
#304995000000
1!
1%
#305000000000
0!
0%
#305005000000
1!
1%
#305010000000
0!
0%
#305015000000
1!
1%
#305020000000
0!
0%
#305025000000
1!
1%
#305030000000
0!
0%
#305035000000
1!
1%
#305040000000
0!
0%
#305045000000
1!
1%
#305050000000
0!
0%
#305055000000
1!
1%
#305060000000
0!
0%
#305065000000
1!
1%
#305070000000
0!
0%
#305075000000
1!
1%
#305080000000
0!
0%
#305085000000
1!
1%
#305090000000
0!
0%
#305095000000
1!
1%
#305100000000
0!
0%
#305105000000
1!
1%
#305110000000
0!
0%
#305115000000
1!
1%
#305120000000
0!
0%
#305125000000
1!
1%
#305130000000
0!
0%
#305135000000
1!
1%
#305140000000
0!
0%
#305145000000
1!
1%
#305150000000
0!
0%
#305155000000
1!
1%
#305160000000
0!
0%
#305165000000
1!
1%
#305170000000
0!
0%
#305175000000
1!
1%
#305180000000
0!
0%
#305185000000
1!
1%
#305190000000
0!
0%
#305195000000
1!
1%
#305200000000
0!
0%
#305205000000
1!
1%
#305210000000
0!
0%
#305215000000
1!
1%
#305220000000
0!
0%
#305225000000
1!
1%
#305230000000
0!
0%
#305235000000
1!
1%
#305240000000
0!
0%
#305245000000
1!
1%
#305250000000
0!
0%
#305255000000
1!
1%
#305260000000
0!
0%
#305265000000
1!
1%
#305270000000
0!
0%
#305275000000
1!
1%
#305280000000
0!
0%
#305285000000
1!
1%
#305290000000
0!
0%
#305295000000
1!
1%
#305300000000
0!
0%
#305305000000
1!
1%
#305310000000
0!
0%
#305315000000
1!
1%
#305320000000
0!
0%
#305325000000
1!
1%
#305330000000
0!
0%
#305335000000
1!
1%
#305340000000
0!
0%
#305345000000
1!
1%
#305350000000
0!
0%
#305355000000
1!
1%
#305360000000
0!
0%
#305365000000
1!
1%
#305370000000
0!
0%
#305375000000
1!
1%
#305380000000
0!
0%
#305385000000
1!
1%
#305390000000
0!
0%
#305395000000
1!
1%
#305400000000
0!
0%
#305405000000
1!
1%
#305410000000
0!
0%
#305415000000
1!
1%
#305420000000
0!
0%
#305425000000
1!
1%
#305430000000
0!
0%
#305435000000
1!
1%
#305440000000
0!
0%
#305445000000
1!
1%
#305450000000
0!
0%
#305455000000
1!
1%
#305460000000
0!
0%
#305465000000
1!
1%
#305470000000
0!
0%
#305475000000
1!
1%
#305480000000
0!
0%
#305485000000
1!
1%
#305490000000
0!
0%
#305495000000
1!
1%
#305500000000
0!
0%
#305505000000
1!
1%
#305510000000
0!
0%
#305515000000
1!
1%
#305520000000
0!
0%
#305525000000
1!
1%
#305530000000
0!
0%
#305535000000
1!
1%
#305540000000
0!
0%
#305545000000
1!
1%
#305550000000
0!
0%
#305555000000
1!
1%
#305560000000
0!
0%
#305565000000
1!
1%
#305570000000
0!
0%
#305575000000
1!
1%
#305580000000
0!
0%
#305585000000
1!
1%
#305590000000
0!
0%
#305595000000
1!
1%
#305600000000
0!
0%
#305605000000
1!
1%
#305610000000
0!
0%
#305615000000
1!
1%
#305620000000
0!
0%
#305625000000
1!
1%
#305630000000
0!
0%
#305635000000
1!
1%
#305640000000
0!
0%
#305645000000
1!
1%
#305650000000
0!
0%
#305655000000
1!
1%
#305660000000
0!
0%
#305665000000
1!
1%
#305670000000
0!
0%
#305675000000
1!
1%
#305680000000
0!
0%
#305685000000
1!
1%
#305690000000
0!
0%
#305695000000
1!
1%
#305700000000
0!
0%
#305705000000
1!
1%
#305710000000
0!
0%
#305715000000
1!
1%
#305720000000
0!
0%
#305725000000
1!
1%
#305730000000
0!
0%
#305735000000
1!
1%
#305740000000
0!
0%
#305745000000
1!
1%
#305750000000
0!
0%
#305755000000
1!
1%
#305760000000
0!
0%
#305765000000
1!
1%
#305770000000
0!
0%
#305775000000
1!
1%
#305780000000
0!
0%
#305785000000
1!
1%
#305790000000
0!
0%
#305795000000
1!
1%
#305800000000
0!
0%
#305805000000
1!
1%
#305810000000
0!
0%
#305815000000
1!
1%
#305820000000
0!
0%
#305825000000
1!
1%
#305830000000
0!
0%
#305835000000
1!
1%
#305840000000
0!
0%
#305845000000
1!
1%
#305850000000
0!
0%
#305855000000
1!
1%
#305860000000
0!
0%
#305865000000
1!
1%
#305870000000
0!
0%
#305875000000
1!
1%
#305880000000
0!
0%
#305885000000
1!
1%
#305890000000
0!
0%
#305895000000
1!
1%
#305900000000
0!
0%
#305905000000
1!
1%
#305910000000
0!
0%
#305915000000
1!
1%
#305920000000
0!
0%
#305925000000
1!
1%
#305930000000
0!
0%
#305935000000
1!
1%
#305940000000
0!
0%
#305945000000
1!
1%
#305950000000
0!
0%
#305955000000
1!
1%
#305960000000
0!
0%
#305965000000
1!
1%
#305970000000
0!
0%
#305975000000
1!
1%
#305980000000
0!
0%
#305985000000
1!
1%
#305990000000
0!
0%
#305995000000
1!
1%
#306000000000
0!
0%
#306005000000
1!
1%
#306010000000
0!
0%
#306015000000
1!
1%
#306020000000
0!
0%
#306025000000
1!
1%
#306030000000
0!
0%
#306035000000
1!
1%
#306040000000
0!
0%
#306045000000
1!
1%
#306050000000
0!
0%
#306055000000
1!
1%
#306060000000
0!
0%
#306065000000
1!
1%
#306070000000
0!
0%
#306075000000
1!
1%
#306080000000
0!
0%
#306085000000
1!
1%
#306090000000
0!
0%
#306095000000
1!
1%
#306100000000
0!
0%
#306105000000
1!
1%
#306110000000
0!
0%
#306115000000
1!
1%
#306120000000
0!
0%
#306125000000
1!
1%
#306130000000
0!
0%
#306135000000
1!
1%
#306140000000
0!
0%
#306145000000
1!
1%
#306150000000
0!
0%
#306155000000
1!
1%
#306160000000
0!
0%
#306165000000
1!
1%
#306170000000
0!
0%
#306175000000
1!
1%
#306180000000
0!
0%
#306185000000
1!
1%
#306190000000
0!
0%
#306195000000
1!
1%
#306200000000
0!
0%
#306205000000
1!
1%
#306210000000
0!
0%
#306215000000
1!
1%
#306220000000
0!
0%
#306225000000
1!
1%
#306230000000
0!
0%
#306235000000
1!
1%
#306240000000
0!
0%
#306245000000
1!
1%
#306250000000
0!
0%
#306255000000
1!
1%
#306260000000
0!
0%
#306265000000
1!
1%
#306270000000
0!
0%
#306275000000
1!
1%
#306280000000
0!
0%
#306285000000
1!
1%
#306290000000
0!
0%
#306295000000
1!
1%
#306300000000
0!
0%
#306305000000
1!
1%
#306310000000
0!
0%
#306315000000
1!
1%
#306320000000
0!
0%
#306325000000
1!
1%
#306330000000
0!
0%
#306335000000
1!
1%
#306340000000
0!
0%
#306345000000
1!
1%
#306350000000
0!
0%
#306355000000
1!
1%
#306360000000
0!
0%
#306365000000
1!
1%
#306370000000
0!
0%
#306375000000
1!
1%
#306380000000
0!
0%
#306385000000
1!
1%
#306390000000
0!
0%
#306395000000
1!
1%
#306400000000
0!
0%
#306405000000
1!
1%
#306410000000
0!
0%
#306415000000
1!
1%
#306420000000
0!
0%
#306425000000
1!
1%
#306430000000
0!
0%
#306435000000
1!
1%
#306440000000
0!
0%
#306445000000
1!
1%
#306450000000
0!
0%
#306455000000
1!
1%
#306460000000
0!
0%
#306465000000
1!
1%
#306470000000
0!
0%
#306475000000
1!
1%
#306480000000
0!
0%
#306485000000
1!
1%
#306490000000
0!
0%
#306495000000
1!
1%
#306500000000
0!
0%
#306505000000
1!
1%
#306510000000
0!
0%
#306515000000
1!
1%
#306520000000
0!
0%
#306525000000
1!
1%
#306530000000
0!
0%
#306535000000
1!
1%
#306540000000
0!
0%
#306545000000
1!
1%
#306550000000
0!
0%
#306555000000
1!
1%
#306560000000
0!
0%
#306565000000
1!
1%
#306570000000
0!
0%
#306575000000
1!
1%
#306580000000
0!
0%
#306585000000
1!
1%
#306590000000
0!
0%
#306595000000
1!
1%
#306600000000
0!
0%
#306605000000
1!
1%
#306610000000
0!
0%
#306615000000
1!
1%
#306620000000
0!
0%
#306625000000
1!
1%
#306630000000
0!
0%
#306635000000
1!
1%
#306640000000
0!
0%
#306645000000
1!
1%
#306650000000
0!
0%
#306655000000
1!
1%
#306660000000
0!
0%
#306665000000
1!
1%
#306670000000
0!
0%
#306675000000
1!
1%
#306680000000
0!
0%
#306685000000
1!
1%
#306690000000
0!
0%
#306695000000
1!
1%
#306700000000
0!
0%
#306705000000
1!
1%
#306710000000
0!
0%
#306715000000
1!
1%
#306720000000
0!
0%
#306725000000
1!
1%
#306730000000
0!
0%
#306735000000
1!
1%
#306740000000
0!
0%
#306745000000
1!
1%
#306750000000
0!
0%
#306755000000
1!
1%
#306760000000
0!
0%
#306765000000
1!
1%
#306770000000
0!
0%
#306775000000
1!
1%
#306780000000
0!
0%
#306785000000
1!
1%
#306790000000
0!
0%
#306795000000
1!
1%
#306800000000
0!
0%
#306805000000
1!
1%
#306810000000
0!
0%
#306815000000
1!
1%
#306820000000
0!
0%
#306825000000
1!
1%
#306830000000
0!
0%
#306835000000
1!
1%
#306840000000
0!
0%
#306845000000
1!
1%
#306850000000
0!
0%
#306855000000
1!
1%
#306860000000
0!
0%
#306865000000
1!
1%
#306870000000
0!
0%
#306875000000
1!
1%
#306880000000
0!
0%
#306885000000
1!
1%
#306890000000
0!
0%
#306895000000
1!
1%
#306900000000
0!
0%
#306905000000
1!
1%
#306910000000
0!
0%
#306915000000
1!
1%
#306920000000
0!
0%
#306925000000
1!
1%
#306930000000
0!
0%
#306935000000
1!
1%
#306940000000
0!
0%
#306945000000
1!
1%
#306950000000
0!
0%
#306955000000
1!
1%
#306960000000
0!
0%
#306965000000
1!
1%
#306970000000
0!
0%
#306975000000
1!
1%
#306980000000
0!
0%
#306985000000
1!
1%
#306990000000
0!
0%
#306995000000
1!
1%
#307000000000
0!
0%
#307005000000
1!
1%
#307010000000
0!
0%
#307015000000
1!
1%
#307020000000
0!
0%
#307025000000
1!
1%
#307030000000
0!
0%
#307035000000
1!
1%
#307040000000
0!
0%
#307045000000
1!
1%
#307050000000
0!
0%
#307055000000
1!
1%
#307060000000
0!
0%
#307065000000
1!
1%
#307070000000
0!
0%
#307075000000
1!
1%
#307080000000
0!
0%
#307085000000
1!
1%
#307090000000
0!
0%
#307095000000
1!
1%
#307100000000
0!
0%
#307105000000
1!
1%
#307110000000
0!
0%
#307115000000
1!
1%
#307120000000
0!
0%
#307125000000
1!
1%
#307130000000
0!
0%
#307135000000
1!
1%
#307140000000
0!
0%
#307145000000
1!
1%
#307150000000
0!
0%
#307155000000
1!
1%
#307160000000
0!
0%
#307165000000
1!
1%
#307170000000
0!
0%
#307175000000
1!
1%
#307180000000
0!
0%
#307185000000
1!
1%
#307190000000
0!
0%
#307195000000
1!
1%
#307200000000
0!
0%
#307205000000
1!
1%
#307210000000
0!
0%
#307215000000
1!
1%
#307220000000
0!
0%
#307225000000
1!
1%
#307230000000
0!
0%
#307235000000
1!
1%
#307240000000
0!
0%
#307245000000
1!
1%
#307250000000
0!
0%
#307255000000
1!
1%
#307260000000
0!
0%
#307265000000
1!
1%
#307270000000
0!
0%
#307275000000
1!
1%
#307280000000
0!
0%
#307285000000
1!
1%
#307290000000
0!
0%
#307295000000
1!
1%
#307300000000
0!
0%
#307305000000
1!
1%
#307310000000
0!
0%
#307315000000
1!
1%
#307320000000
0!
0%
#307325000000
1!
1%
#307330000000
0!
0%
#307335000000
1!
1%
#307340000000
0!
0%
#307345000000
1!
1%
#307350000000
0!
0%
#307355000000
1!
1%
#307360000000
0!
0%
#307365000000
1!
1%
#307370000000
0!
0%
#307375000000
1!
1%
#307380000000
0!
0%
#307385000000
1!
1%
#307390000000
0!
0%
#307395000000
1!
1%
#307400000000
0!
0%
#307405000000
1!
1%
#307410000000
0!
0%
#307415000000
1!
1%
#307420000000
0!
0%
#307425000000
1!
1%
#307430000000
0!
0%
#307435000000
1!
1%
#307440000000
0!
0%
#307445000000
1!
1%
#307450000000
0!
0%
#307455000000
1!
1%
#307460000000
0!
0%
#307465000000
1!
1%
#307470000000
0!
0%
#307475000000
1!
1%
#307480000000
0!
0%
#307485000000
1!
1%
#307490000000
0!
0%
#307495000000
1!
1%
#307500000000
0!
0%
#307505000000
1!
1%
#307510000000
0!
0%
#307515000000
1!
1%
#307520000000
0!
0%
#307525000000
1!
1%
#307530000000
0!
0%
#307535000000
1!
1%
#307540000000
0!
0%
#307545000000
1!
1%
#307550000000
0!
0%
#307555000000
1!
1%
#307560000000
0!
0%
#307565000000
1!
1%
#307570000000
0!
0%
#307575000000
1!
1%
#307580000000
0!
0%
#307585000000
1!
1%
#307590000000
0!
0%
#307595000000
1!
1%
#307600000000
0!
0%
#307605000000
1!
1%
#307610000000
0!
0%
#307615000000
1!
1%
#307620000000
0!
0%
#307625000000
1!
1%
#307630000000
0!
0%
#307635000000
1!
1%
#307640000000
0!
0%
#307645000000
1!
1%
#307650000000
0!
0%
#307655000000
1!
1%
#307660000000
0!
0%
#307665000000
1!
1%
#307670000000
0!
0%
#307675000000
1!
1%
#307680000000
0!
0%
#307685000000
1!
1%
#307690000000
0!
0%
#307695000000
1!
1%
#307700000000
0!
0%
#307705000000
1!
1%
#307710000000
0!
0%
#307715000000
1!
1%
#307720000000
0!
0%
#307725000000
1!
1%
#307730000000
0!
0%
#307735000000
1!
1%
#307740000000
0!
0%
#307745000000
1!
1%
#307750000000
0!
0%
#307755000000
1!
1%
#307760000000
0!
0%
#307765000000
1!
1%
#307770000000
0!
0%
#307775000000
1!
1%
#307780000000
0!
0%
#307785000000
1!
1%
#307790000000
0!
0%
#307795000000
1!
1%
#307800000000
0!
0%
#307805000000
1!
1%
#307810000000
0!
0%
#307815000000
1!
1%
#307820000000
0!
0%
#307825000000
1!
1%
#307830000000
0!
0%
#307835000000
1!
1%
#307840000000
0!
0%
#307845000000
1!
1%
#307850000000
0!
0%
#307855000000
1!
1%
#307860000000
0!
0%
#307865000000
1!
1%
#307870000000
0!
0%
#307875000000
1!
1%
#307880000000
0!
0%
#307885000000
1!
1%
#307890000000
0!
0%
#307895000000
1!
1%
#307900000000
0!
0%
#307905000000
1!
1%
#307910000000
0!
0%
#307915000000
1!
1%
#307920000000
0!
0%
#307925000000
1!
1%
#307930000000
0!
0%
#307935000000
1!
1%
#307940000000
0!
0%
#307945000000
1!
1%
#307950000000
0!
0%
#307955000000
1!
1%
#307960000000
0!
0%
#307965000000
1!
1%
#307970000000
0!
0%
#307975000000
1!
1%
#307980000000
0!
0%
#307985000000
1!
1%
#307990000000
0!
0%
#307995000000
1!
1%
#308000000000
0!
0%
#308005000000
1!
1%
#308010000000
0!
0%
#308015000000
1!
1%
#308020000000
0!
0%
#308025000000
1!
1%
#308030000000
0!
0%
#308035000000
1!
1%
#308040000000
0!
0%
#308045000000
1!
1%
#308050000000
0!
0%
#308055000000
1!
1%
#308060000000
0!
0%
#308065000000
1!
1%
#308070000000
0!
0%
#308075000000
1!
1%
#308080000000
0!
0%
#308085000000
1!
1%
#308090000000
0!
0%
#308095000000
1!
1%
#308100000000
0!
0%
#308105000000
1!
1%
#308110000000
0!
0%
#308115000000
1!
1%
#308120000000
0!
0%
#308125000000
1!
1%
#308130000000
0!
0%
#308135000000
1!
1%
#308140000000
0!
0%
#308145000000
1!
1%
#308150000000
0!
0%
#308155000000
1!
1%
#308160000000
0!
0%
#308165000000
1!
1%
#308170000000
0!
0%
#308175000000
1!
1%
#308180000000
0!
0%
#308185000000
1!
1%
#308190000000
0!
0%
#308195000000
1!
1%
#308200000000
0!
0%
#308205000000
1!
1%
#308210000000
0!
0%
#308215000000
1!
1%
#308220000000
0!
0%
#308225000000
1!
1%
#308230000000
0!
0%
#308235000000
1!
1%
#308240000000
0!
0%
#308245000000
1!
1%
#308250000000
0!
0%
#308255000000
1!
1%
#308260000000
0!
0%
#308265000000
1!
1%
#308270000000
0!
0%
#308275000000
1!
1%
#308280000000
0!
0%
#308285000000
1!
1%
#308290000000
0!
0%
#308295000000
1!
1%
#308300000000
0!
0%
#308305000000
1!
1%
#308310000000
0!
0%
#308315000000
1!
1%
#308320000000
0!
0%
#308325000000
1!
1%
#308330000000
0!
0%
#308335000000
1!
1%
#308340000000
0!
0%
#308345000000
1!
1%
#308350000000
0!
0%
#308355000000
1!
1%
#308360000000
0!
0%
#308365000000
1!
1%
#308370000000
0!
0%
#308375000000
1!
1%
#308380000000
0!
0%
#308385000000
1!
1%
#308390000000
0!
0%
#308395000000
1!
1%
#308400000000
0!
0%
#308405000000
1!
1%
#308410000000
0!
0%
#308415000000
1!
1%
#308420000000
0!
0%
#308425000000
1!
1%
#308430000000
0!
0%
#308435000000
1!
1%
#308440000000
0!
0%
#308445000000
1!
1%
#308450000000
0!
0%
#308455000000
1!
1%
#308460000000
0!
0%
#308465000000
1!
1%
#308470000000
0!
0%
#308475000000
1!
1%
#308480000000
0!
0%
#308485000000
1!
1%
#308490000000
0!
0%
#308495000000
1!
1%
#308500000000
0!
0%
#308505000000
1!
1%
#308510000000
0!
0%
#308515000000
1!
1%
#308520000000
0!
0%
#308525000000
1!
1%
#308530000000
0!
0%
#308535000000
1!
1%
#308540000000
0!
0%
#308545000000
1!
1%
#308550000000
0!
0%
#308555000000
1!
1%
#308560000000
0!
0%
#308565000000
1!
1%
#308570000000
0!
0%
#308575000000
1!
1%
#308580000000
0!
0%
#308585000000
1!
1%
#308590000000
0!
0%
#308595000000
1!
1%
#308600000000
0!
0%
#308605000000
1!
1%
#308610000000
0!
0%
#308615000000
1!
1%
#308620000000
0!
0%
#308625000000
1!
1%
#308630000000
0!
0%
#308635000000
1!
1%
#308640000000
0!
0%
#308645000000
1!
1%
#308650000000
0!
0%
#308655000000
1!
1%
#308660000000
0!
0%
#308665000000
1!
1%
#308670000000
0!
0%
#308675000000
1!
1%
#308680000000
0!
0%
#308685000000
1!
1%
#308690000000
0!
0%
#308695000000
1!
1%
#308700000000
0!
0%
#308705000000
1!
1%
#308710000000
0!
0%
#308715000000
1!
1%
#308720000000
0!
0%
#308725000000
1!
1%
#308730000000
0!
0%
#308735000000
1!
1%
#308740000000
0!
0%
#308745000000
1!
1%
#308750000000
0!
0%
#308755000000
1!
1%
#308760000000
0!
0%
#308765000000
1!
1%
#308770000000
0!
0%
#308775000000
1!
1%
#308780000000
0!
0%
#308785000000
1!
1%
#308790000000
0!
0%
#308795000000
1!
1%
#308800000000
0!
0%
#308805000000
1!
1%
#308810000000
0!
0%
#308815000000
1!
1%
#308820000000
0!
0%
#308825000000
1!
1%
#308830000000
0!
0%
#308835000000
1!
1%
#308840000000
0!
0%
#308845000000
1!
1%
#308850000000
0!
0%
#308855000000
1!
1%
#308860000000
0!
0%
#308865000000
1!
1%
#308870000000
0!
0%
#308875000000
1!
1%
#308880000000
0!
0%
#308885000000
1!
1%
#308890000000
0!
0%
#308895000000
1!
1%
#308900000000
0!
0%
#308905000000
1!
1%
#308910000000
0!
0%
#308915000000
1!
1%
#308920000000
0!
0%
#308925000000
1!
1%
#308930000000
0!
0%
#308935000000
1!
1%
#308940000000
0!
0%
#308945000000
1!
1%
#308950000000
0!
0%
#308955000000
1!
1%
#308960000000
0!
0%
#308965000000
1!
1%
#308970000000
0!
0%
#308975000000
1!
1%
#308980000000
0!
0%
#308985000000
1!
1%
#308990000000
0!
0%
#308995000000
1!
1%
#309000000000
0!
0%
#309005000000
1!
1%
#309010000000
0!
0%
#309015000000
1!
1%
#309020000000
0!
0%
#309025000000
1!
1%
#309030000000
0!
0%
#309035000000
1!
1%
#309040000000
0!
0%
#309045000000
1!
1%
#309050000000
0!
0%
#309055000000
1!
1%
#309060000000
0!
0%
#309065000000
1!
1%
#309070000000
0!
0%
#309075000000
1!
1%
#309080000000
0!
0%
#309085000000
1!
1%
#309090000000
0!
0%
#309095000000
1!
1%
#309100000000
0!
0%
#309105000000
1!
1%
#309110000000
0!
0%
#309115000000
1!
1%
#309120000000
0!
0%
#309125000000
1!
1%
#309130000000
0!
0%
#309135000000
1!
1%
#309140000000
0!
0%
#309145000000
1!
1%
#309150000000
0!
0%
#309155000000
1!
1%
#309160000000
0!
0%
#309165000000
1!
1%
#309170000000
0!
0%
#309175000000
1!
1%
#309180000000
0!
0%
#309185000000
1!
1%
#309190000000
0!
0%
#309195000000
1!
1%
#309200000000
0!
0%
#309205000000
1!
1%
#309210000000
0!
0%
#309215000000
1!
1%
#309220000000
0!
0%
#309225000000
1!
1%
#309230000000
0!
0%
#309235000000
1!
1%
#309240000000
0!
0%
#309245000000
1!
1%
#309250000000
0!
0%
#309255000000
1!
1%
#309260000000
0!
0%
#309265000000
1!
1%
#309270000000
0!
0%
#309275000000
1!
1%
#309280000000
0!
0%
#309285000000
1!
1%
#309290000000
0!
0%
#309295000000
1!
1%
#309300000000
0!
0%
#309305000000
1!
1%
#309310000000
0!
0%
#309315000000
1!
1%
#309320000000
0!
0%
#309325000000
1!
1%
#309330000000
0!
0%
#309335000000
1!
1%
#309340000000
0!
0%
#309345000000
1!
1%
#309350000000
0!
0%
#309355000000
1!
1%
#309360000000
0!
0%
#309365000000
1!
1%
#309370000000
0!
0%
#309375000000
1!
1%
#309380000000
0!
0%
#309385000000
1!
1%
#309390000000
0!
0%
#309395000000
1!
1%
#309400000000
0!
0%
#309405000000
1!
1%
#309410000000
0!
0%
#309415000000
1!
1%
#309420000000
0!
0%
#309425000000
1!
1%
#309430000000
0!
0%
#309435000000
1!
1%
#309440000000
0!
0%
#309445000000
1!
1%
#309450000000
0!
0%
#309455000000
1!
1%
#309460000000
0!
0%
#309465000000
1!
1%
#309470000000
0!
0%
#309475000000
1!
1%
#309480000000
0!
0%
#309485000000
1!
1%
#309490000000
0!
0%
#309495000000
1!
1%
#309500000000
0!
0%
#309505000000
1!
1%
#309510000000
0!
0%
#309515000000
1!
1%
#309520000000
0!
0%
#309525000000
1!
1%
#309530000000
0!
0%
#309535000000
1!
1%
#309540000000
0!
0%
#309545000000
1!
1%
#309550000000
0!
0%
#309555000000
1!
1%
#309560000000
0!
0%
#309565000000
1!
1%
#309570000000
0!
0%
#309575000000
1!
1%
#309580000000
0!
0%
#309585000000
1!
1%
#309590000000
0!
0%
#309595000000
1!
1%
#309600000000
0!
0%
#309605000000
1!
1%
#309610000000
0!
0%
#309615000000
1!
1%
#309620000000
0!
0%
#309625000000
1!
1%
#309630000000
0!
0%
#309635000000
1!
1%
#309640000000
0!
0%
#309645000000
1!
1%
#309650000000
0!
0%
#309655000000
1!
1%
#309660000000
0!
0%
#309665000000
1!
1%
#309670000000
0!
0%
#309675000000
1!
1%
#309680000000
0!
0%
#309685000000
1!
1%
#309690000000
0!
0%
#309695000000
1!
1%
#309700000000
0!
0%
#309705000000
1!
1%
#309710000000
0!
0%
#309715000000
1!
1%
#309720000000
0!
0%
#309725000000
1!
1%
#309730000000
0!
0%
#309735000000
1!
1%
#309740000000
0!
0%
#309745000000
1!
1%
#309750000000
0!
0%
#309755000000
1!
1%
#309760000000
0!
0%
#309765000000
1!
1%
#309770000000
0!
0%
#309775000000
1!
1%
#309780000000
0!
0%
#309785000000
1!
1%
#309790000000
0!
0%
#309795000000
1!
1%
#309800000000
0!
0%
#309805000000
1!
1%
#309810000000
0!
0%
#309815000000
1!
1%
#309820000000
0!
0%
#309825000000
1!
1%
#309830000000
0!
0%
#309835000000
1!
1%
#309840000000
0!
0%
#309845000000
1!
1%
#309850000000
0!
0%
#309855000000
1!
1%
#309860000000
0!
0%
#309865000000
1!
1%
#309870000000
0!
0%
#309875000000
1!
1%
#309880000000
0!
0%
#309885000000
1!
1%
#309890000000
0!
0%
#309895000000
1!
1%
#309900000000
0!
0%
#309905000000
1!
1%
#309910000000
0!
0%
#309915000000
1!
1%
#309920000000
0!
0%
#309925000000
1!
1%
#309930000000
0!
0%
#309935000000
1!
1%
#309940000000
0!
0%
#309945000000
1!
1%
#309950000000
0!
0%
#309955000000
1!
1%
#309960000000
0!
0%
#309965000000
1!
1%
#309970000000
0!
0%
#309975000000
1!
1%
#309980000000
0!
0%
#309985000000
1!
1%
#309990000000
0!
0%
#309995000000
1!
1%
#310000000000
0!
0%
#310005000000
1!
1%
#310010000000
0!
0%
#310015000000
1!
1%
#310020000000
0!
0%
#310025000000
1!
1%
#310030000000
0!
0%
#310035000000
1!
1%
#310040000000
0!
0%
#310045000000
1!
1%
#310050000000
0!
0%
#310055000000
1!
1%
#310060000000
0!
0%
#310065000000
1!
1%
#310070000000
0!
0%
#310075000000
1!
1%
#310080000000
0!
0%
#310085000000
1!
1%
#310090000000
0!
0%
#310095000000
1!
1%
#310100000000
0!
0%
#310105000000
1!
1%
#310110000000
0!
0%
#310115000000
1!
1%
#310120000000
0!
0%
#310125000000
1!
1%
#310130000000
0!
0%
#310135000000
1!
1%
#310140000000
0!
0%
#310145000000
1!
1%
#310150000000
0!
0%
#310155000000
1!
1%
#310160000000
0!
0%
#310165000000
1!
1%
#310170000000
0!
0%
#310175000000
1!
1%
#310180000000
0!
0%
#310185000000
1!
1%
#310190000000
0!
0%
#310195000000
1!
1%
#310200000000
0!
0%
#310205000000
1!
1%
#310210000000
0!
0%
#310215000000
1!
1%
#310220000000
0!
0%
#310225000000
1!
1%
#310230000000
0!
0%
#310235000000
1!
1%
#310240000000
0!
0%
#310245000000
1!
1%
#310250000000
0!
0%
#310255000000
1!
1%
#310260000000
0!
0%
#310265000000
1!
1%
#310270000000
0!
0%
#310275000000
1!
1%
#310280000000
0!
0%
#310285000000
1!
1%
#310290000000
0!
0%
#310295000000
1!
1%
#310300000000
0!
0%
#310305000000
1!
1%
#310310000000
0!
0%
#310315000000
1!
1%
#310320000000
0!
0%
#310325000000
1!
1%
#310330000000
0!
0%
#310335000000
1!
1%
#310340000000
0!
0%
#310345000000
1!
1%
#310350000000
0!
0%
#310355000000
1!
1%
#310360000000
0!
0%
#310365000000
1!
1%
#310370000000
0!
0%
#310375000000
1!
1%
#310380000000
0!
0%
#310385000000
1!
1%
#310390000000
0!
0%
#310395000000
1!
1%
#310400000000
0!
0%
#310405000000
1!
1%
#310410000000
0!
0%
#310415000000
1!
1%
#310420000000
0!
0%
#310425000000
1!
1%
#310430000000
0!
0%
#310435000000
1!
1%
#310440000000
0!
0%
#310445000000
1!
1%
#310450000000
0!
0%
#310455000000
1!
1%
#310460000000
0!
0%
#310465000000
1!
1%
#310470000000
0!
0%
#310475000000
1!
1%
#310480000000
0!
0%
#310485000000
1!
1%
#310490000000
0!
0%
#310495000000
1!
1%
#310500000000
0!
0%
#310505000000
1!
1%
#310510000000
0!
0%
#310515000000
1!
1%
#310520000000
0!
0%
#310525000000
1!
1%
#310530000000
0!
0%
#310535000000
1!
1%
#310540000000
0!
0%
#310545000000
1!
1%
#310550000000
0!
0%
#310555000000
1!
1%
#310560000000
0!
0%
#310565000000
1!
1%
#310570000000
0!
0%
#310575000000
1!
1%
#310580000000
0!
0%
#310585000000
1!
1%
#310590000000
0!
0%
#310595000000
1!
1%
#310600000000
0!
0%
#310605000000
1!
1%
#310610000000
0!
0%
#310615000000
1!
1%
#310620000000
0!
0%
#310625000000
1!
1%
#310630000000
0!
0%
#310635000000
1!
1%
#310640000000
0!
0%
#310645000000
1!
1%
#310650000000
0!
0%
#310655000000
1!
1%
#310660000000
0!
0%
#310665000000
1!
1%
#310670000000
0!
0%
#310675000000
1!
1%
#310680000000
0!
0%
#310685000000
1!
1%
#310690000000
0!
0%
#310695000000
1!
1%
#310700000000
0!
0%
#310705000000
1!
1%
#310710000000
0!
0%
#310715000000
1!
1%
#310720000000
0!
0%
#310725000000
1!
1%
#310730000000
0!
0%
#310735000000
1!
1%
#310740000000
0!
0%
#310745000000
1!
1%
#310750000000
0!
0%
#310755000000
1!
1%
#310760000000
0!
0%
#310765000000
1!
1%
#310770000000
0!
0%
#310775000000
1!
1%
#310780000000
0!
0%
#310785000000
1!
1%
#310790000000
0!
0%
#310795000000
1!
1%
#310800000000
0!
0%
#310805000000
1!
1%
#310810000000
0!
0%
#310815000000
1!
1%
#310820000000
0!
0%
#310825000000
1!
1%
#310830000000
0!
0%
#310835000000
1!
1%
#310840000000
0!
0%
#310845000000
1!
1%
#310850000000
0!
0%
#310855000000
1!
1%
#310860000000
0!
0%
#310865000000
1!
1%
#310870000000
0!
0%
#310875000000
1!
1%
#310880000000
0!
0%
#310885000000
1!
1%
#310890000000
0!
0%
#310895000000
1!
1%
#310900000000
0!
0%
#310905000000
1!
1%
#310910000000
0!
0%
#310915000000
1!
1%
#310920000000
0!
0%
#310925000000
1!
1%
#310930000000
0!
0%
#310935000000
1!
1%
#310940000000
0!
0%
#310945000000
1!
1%
#310950000000
0!
0%
#310955000000
1!
1%
#310960000000
0!
0%
#310965000000
1!
1%
#310970000000
0!
0%
#310975000000
1!
1%
#310980000000
0!
0%
#310985000000
1!
1%
#310990000000
0!
0%
#310995000000
1!
1%
#311000000000
0!
0%
#311005000000
1!
1%
#311010000000
0!
0%
#311015000000
1!
1%
#311020000000
0!
0%
#311025000000
1!
1%
#311030000000
0!
0%
#311035000000
1!
1%
#311040000000
0!
0%
#311045000000
1!
1%
#311050000000
0!
0%
#311055000000
1!
1%
#311060000000
0!
0%
#311065000000
1!
1%
#311070000000
0!
0%
#311075000000
1!
1%
#311080000000
0!
0%
#311085000000
1!
1%
#311090000000
0!
0%
#311095000000
1!
1%
#311100000000
0!
0%
#311105000000
1!
1%
#311110000000
0!
0%
#311115000000
1!
1%
#311120000000
0!
0%
#311125000000
1!
1%
#311130000000
0!
0%
#311135000000
1!
1%
#311140000000
0!
0%
#311145000000
1!
1%
#311150000000
0!
0%
#311155000000
1!
1%
#311160000000
0!
0%
#311165000000
1!
1%
#311170000000
0!
0%
#311175000000
1!
1%
#311180000000
0!
0%
#311185000000
1!
1%
#311190000000
0!
0%
#311195000000
1!
1%
#311200000000
0!
0%
#311205000000
1!
1%
#311210000000
0!
0%
#311215000000
1!
1%
#311220000000
0!
0%
#311225000000
1!
1%
#311230000000
0!
0%
#311235000000
1!
1%
#311240000000
0!
0%
#311245000000
1!
1%
#311250000000
0!
0%
#311255000000
1!
1%
#311260000000
0!
0%
#311265000000
1!
1%
#311270000000
0!
0%
#311275000000
1!
1%
#311280000000
0!
0%
#311285000000
1!
1%
#311290000000
0!
0%
#311295000000
1!
1%
#311300000000
0!
0%
#311305000000
1!
1%
#311310000000
0!
0%
#311315000000
1!
1%
#311320000000
0!
0%
#311325000000
1!
1%
#311330000000
0!
0%
#311335000000
1!
1%
#311340000000
0!
0%
#311345000000
1!
1%
#311350000000
0!
0%
#311355000000
1!
1%
#311360000000
0!
0%
#311365000000
1!
1%
#311370000000
0!
0%
#311375000000
1!
1%
#311380000000
0!
0%
#311385000000
1!
1%
#311390000000
0!
0%
#311395000000
1!
1%
#311400000000
0!
0%
#311405000000
1!
1%
#311410000000
0!
0%
#311415000000
1!
1%
#311420000000
0!
0%
#311425000000
1!
1%
#311430000000
0!
0%
#311435000000
1!
1%
#311440000000
0!
0%
#311445000000
1!
1%
#311450000000
0!
0%
#311455000000
1!
1%
#311460000000
0!
0%
#311465000000
1!
1%
#311470000000
0!
0%
#311475000000
1!
1%
#311480000000
0!
0%
#311485000000
1!
1%
#311490000000
0!
0%
#311495000000
1!
1%
#311500000000
0!
0%
#311505000000
1!
1%
#311510000000
0!
0%
#311515000000
1!
1%
#311520000000
0!
0%
#311525000000
1!
1%
#311530000000
0!
0%
#311535000000
1!
1%
#311540000000
0!
0%
#311545000000
1!
1%
#311550000000
0!
0%
#311555000000
1!
1%
#311560000000
0!
0%
#311565000000
1!
1%
#311570000000
0!
0%
#311575000000
1!
1%
#311580000000
0!
0%
#311585000000
1!
1%
#311590000000
0!
0%
#311595000000
1!
1%
#311600000000
0!
0%
#311605000000
1!
1%
#311610000000
0!
0%
#311615000000
1!
1%
#311620000000
0!
0%
#311625000000
1!
1%
#311630000000
0!
0%
#311635000000
1!
1%
#311640000000
0!
0%
#311645000000
1!
1%
#311650000000
0!
0%
#311655000000
1!
1%
#311660000000
0!
0%
#311665000000
1!
1%
#311670000000
0!
0%
#311675000000
1!
1%
#311680000000
0!
0%
#311685000000
1!
1%
#311690000000
0!
0%
#311695000000
1!
1%
#311700000000
0!
0%
#311705000000
1!
1%
#311710000000
0!
0%
#311715000000
1!
1%
#311720000000
0!
0%
#311725000000
1!
1%
#311730000000
0!
0%
#311735000000
1!
1%
#311740000000
0!
0%
#311745000000
1!
1%
#311750000000
0!
0%
#311755000000
1!
1%
#311760000000
0!
0%
#311765000000
1!
1%
#311770000000
0!
0%
#311775000000
1!
1%
#311780000000
0!
0%
#311785000000
1!
1%
#311790000000
0!
0%
#311795000000
1!
1%
#311800000000
0!
0%
#311805000000
1!
1%
#311810000000
0!
0%
#311815000000
1!
1%
#311820000000
0!
0%
#311825000000
1!
1%
#311830000000
0!
0%
#311835000000
1!
1%
#311840000000
0!
0%
#311845000000
1!
1%
#311850000000
0!
0%
#311855000000
1!
1%
#311860000000
0!
0%
#311865000000
1!
1%
#311870000000
0!
0%
#311875000000
1!
1%
#311880000000
0!
0%
#311885000000
1!
1%
#311890000000
0!
0%
#311895000000
1!
1%
#311900000000
0!
0%
#311905000000
1!
1%
#311910000000
0!
0%
#311915000000
1!
1%
#311920000000
0!
0%
#311925000000
1!
1%
#311930000000
0!
0%
#311935000000
1!
1%
#311940000000
0!
0%
#311945000000
1!
1%
#311950000000
0!
0%
#311955000000
1!
1%
#311960000000
0!
0%
#311965000000
1!
1%
#311970000000
0!
0%
#311975000000
1!
1%
#311980000000
0!
0%
#311985000000
1!
1%
#311990000000
0!
0%
#311995000000
1!
1%
#312000000000
0!
0%
#312005000000
1!
1%
#312010000000
0!
0%
#312015000000
1!
1%
#312020000000
0!
0%
#312025000000
1!
1%
#312030000000
0!
0%
#312035000000
1!
1%
#312040000000
0!
0%
#312045000000
1!
1%
#312050000000
0!
0%
#312055000000
1!
1%
#312060000000
0!
0%
#312065000000
1!
1%
#312070000000
0!
0%
#312075000000
1!
1%
#312080000000
0!
0%
#312085000000
1!
1%
#312090000000
0!
0%
#312095000000
1!
1%
#312100000000
0!
0%
#312105000000
1!
1%
#312110000000
0!
0%
#312115000000
1!
1%
#312120000000
0!
0%
#312125000000
1!
1%
#312130000000
0!
0%
#312135000000
1!
1%
#312140000000
0!
0%
#312145000000
1!
1%
#312150000000
0!
0%
#312155000000
1!
1%
#312160000000
0!
0%
#312165000000
1!
1%
#312170000000
0!
0%
#312175000000
1!
1%
#312180000000
0!
0%
#312185000000
1!
1%
#312190000000
0!
0%
#312195000000
1!
1%
#312200000000
0!
0%
#312205000000
1!
1%
#312210000000
0!
0%
#312215000000
1!
1%
#312220000000
0!
0%
#312225000000
1!
1%
#312230000000
0!
0%
#312235000000
1!
1%
#312240000000
0!
0%
#312245000000
1!
1%
#312250000000
0!
0%
#312255000000
1!
1%
#312260000000
0!
0%
#312265000000
1!
1%
#312270000000
0!
0%
#312275000000
1!
1%
#312280000000
0!
0%
#312285000000
1!
1%
#312290000000
0!
0%
#312295000000
1!
1%
#312300000000
0!
0%
#312305000000
1!
1%
#312310000000
0!
0%
#312315000000
1!
1%
#312320000000
0!
0%
#312325000000
1!
1%
#312330000000
0!
0%
#312335000000
1!
1%
#312340000000
0!
0%
#312345000000
1!
1%
#312350000000
0!
0%
#312355000000
1!
1%
#312360000000
0!
0%
#312365000000
1!
1%
#312370000000
0!
0%
#312375000000
1!
1%
#312380000000
0!
0%
#312385000000
1!
1%
#312390000000
0!
0%
#312395000000
1!
1%
#312400000000
0!
0%
#312405000000
1!
1%
#312410000000
0!
0%
#312415000000
1!
1%
#312420000000
0!
0%
#312425000000
1!
1%
#312430000000
0!
0%
#312435000000
1!
1%
#312440000000
0!
0%
#312445000000
1!
1%
#312450000000
0!
0%
#312455000000
1!
1%
#312460000000
0!
0%
#312465000000
1!
1%
#312470000000
0!
0%
#312475000000
1!
1%
#312480000000
0!
0%
#312485000000
1!
1%
#312490000000
0!
0%
#312495000000
1!
1%
#312500000000
0!
0%
#312505000000
1!
1%
#312510000000
0!
0%
#312515000000
1!
1%
#312520000000
0!
0%
#312525000000
1!
1%
#312530000000
0!
0%
#312535000000
1!
1%
#312540000000
0!
0%
#312545000000
1!
1%
#312550000000
0!
0%
#312555000000
1!
1%
#312560000000
0!
0%
#312565000000
1!
1%
#312570000000
0!
0%
#312575000000
1!
1%
#312580000000
0!
0%
#312585000000
1!
1%
#312590000000
0!
0%
#312595000000
1!
1%
#312600000000
0!
0%
#312605000000
1!
1%
#312610000000
0!
0%
#312615000000
1!
1%
#312620000000
0!
0%
#312625000000
1!
1%
#312630000000
0!
0%
#312635000000
1!
1%
#312640000000
0!
0%
#312645000000
1!
1%
#312650000000
0!
0%
#312655000000
1!
1%
#312660000000
0!
0%
#312665000000
1!
1%
#312670000000
0!
0%
#312675000000
1!
1%
#312680000000
0!
0%
#312685000000
1!
1%
#312690000000
0!
0%
#312695000000
1!
1%
#312700000000
0!
0%
#312705000000
1!
1%
#312710000000
0!
0%
#312715000000
1!
1%
#312720000000
0!
0%
#312725000000
1!
1%
#312730000000
0!
0%
#312735000000
1!
1%
#312740000000
0!
0%
#312745000000
1!
1%
#312750000000
0!
0%
#312755000000
1!
1%
#312760000000
0!
0%
#312765000000
1!
1%
#312770000000
0!
0%
#312775000000
1!
1%
#312780000000
0!
0%
#312785000000
1!
1%
#312790000000
0!
0%
#312795000000
1!
1%
#312800000000
0!
0%
#312805000000
1!
1%
#312810000000
0!
0%
#312815000000
1!
1%
#312820000000
0!
0%
#312825000000
1!
1%
#312830000000
0!
0%
#312835000000
1!
1%
#312840000000
0!
0%
#312845000000
1!
1%
#312850000000
0!
0%
#312855000000
1!
1%
#312860000000
0!
0%
#312865000000
1!
1%
#312870000000
0!
0%
#312875000000
1!
1%
#312880000000
0!
0%
#312885000000
1!
1%
#312890000000
0!
0%
#312895000000
1!
1%
#312900000000
0!
0%
#312905000000
1!
1%
#312910000000
0!
0%
#312915000000
1!
1%
#312920000000
0!
0%
#312925000000
1!
1%
#312930000000
0!
0%
#312935000000
1!
1%
#312940000000
0!
0%
#312945000000
1!
1%
#312950000000
0!
0%
#312955000000
1!
1%
#312960000000
0!
0%
#312965000000
1!
1%
#312970000000
0!
0%
#312975000000
1!
1%
#312980000000
0!
0%
#312985000000
1!
1%
#312990000000
0!
0%
#312995000000
1!
1%
#313000000000
0!
0%
#313005000000
1!
1%
#313010000000
0!
0%
#313015000000
1!
1%
#313020000000
0!
0%
#313025000000
1!
1%
#313030000000
0!
0%
#313035000000
1!
1%
#313040000000
0!
0%
#313045000000
1!
1%
#313050000000
0!
0%
#313055000000
1!
1%
#313060000000
0!
0%
#313065000000
1!
1%
#313070000000
0!
0%
#313075000000
1!
1%
#313080000000
0!
0%
#313085000000
1!
1%
#313090000000
0!
0%
#313095000000
1!
1%
#313100000000
0!
0%
#313105000000
1!
1%
#313110000000
0!
0%
#313115000000
1!
1%
#313120000000
0!
0%
#313125000000
1!
1%
#313130000000
0!
0%
#313135000000
1!
1%
#313140000000
0!
0%
#313145000000
1!
1%
#313150000000
0!
0%
#313155000000
1!
1%
#313160000000
0!
0%
#313165000000
1!
1%
#313170000000
0!
0%
#313175000000
1!
1%
#313180000000
0!
0%
#313185000000
1!
1%
#313190000000
0!
0%
#313195000000
1!
1%
#313200000000
0!
0%
#313205000000
1!
1%
#313210000000
0!
0%
#313215000000
1!
1%
#313220000000
0!
0%
#313225000000
1!
1%
#313230000000
0!
0%
#313235000000
1!
1%
#313240000000
0!
0%
#313245000000
1!
1%
#313250000000
0!
0%
#313255000000
1!
1%
#313260000000
0!
0%
#313265000000
1!
1%
#313270000000
0!
0%
#313275000000
1!
1%
#313280000000
0!
0%
#313285000000
1!
1%
#313290000000
0!
0%
#313295000000
1!
1%
#313300000000
0!
0%
#313305000000
1!
1%
#313310000000
0!
0%
#313315000000
1!
1%
#313320000000
0!
0%
#313325000000
1!
1%
#313330000000
0!
0%
#313335000000
1!
1%
#313340000000
0!
0%
#313345000000
1!
1%
#313350000000
0!
0%
#313355000000
1!
1%
#313360000000
0!
0%
#313365000000
1!
1%
#313370000000
0!
0%
#313375000000
1!
1%
#313380000000
0!
0%
#313385000000
1!
1%
#313390000000
0!
0%
#313395000000
1!
1%
#313400000000
0!
0%
#313405000000
1!
1%
#313410000000
0!
0%
#313415000000
1!
1%
#313420000000
0!
0%
#313425000000
1!
1%
#313430000000
0!
0%
#313435000000
1!
1%
#313440000000
0!
0%
#313445000000
1!
1%
#313450000000
0!
0%
#313455000000
1!
1%
#313460000000
0!
0%
#313465000000
1!
1%
#313470000000
0!
0%
#313475000000
1!
1%
#313480000000
0!
0%
#313485000000
1!
1%
#313490000000
0!
0%
#313495000000
1!
1%
#313500000000
0!
0%
#313505000000
1!
1%
#313510000000
0!
0%
#313515000000
1!
1%
#313520000000
0!
0%
#313525000000
1!
1%
#313530000000
0!
0%
#313535000000
1!
1%
#313540000000
0!
0%
#313545000000
1!
1%
#313550000000
0!
0%
#313555000000
1!
1%
#313560000000
0!
0%
#313565000000
1!
1%
#313570000000
0!
0%
#313575000000
1!
1%
#313580000000
0!
0%
#313585000000
1!
1%
#313590000000
0!
0%
#313595000000
1!
1%
#313600000000
0!
0%
#313605000000
1!
1%
#313610000000
0!
0%
#313615000000
1!
1%
#313620000000
0!
0%
#313625000000
1!
1%
#313630000000
0!
0%
#313635000000
1!
1%
#313640000000
0!
0%
#313645000000
1!
1%
#313650000000
0!
0%
#313655000000
1!
1%
#313660000000
0!
0%
#313665000000
1!
1%
#313670000000
0!
0%
#313675000000
1!
1%
#313680000000
0!
0%
#313685000000
1!
1%
#313690000000
0!
0%
#313695000000
1!
1%
#313700000000
0!
0%
#313705000000
1!
1%
#313710000000
0!
0%
#313715000000
1!
1%
#313720000000
0!
0%
#313725000000
1!
1%
#313730000000
0!
0%
#313735000000
1!
1%
#313740000000
0!
0%
#313745000000
1!
1%
#313750000000
0!
0%
#313755000000
1!
1%
#313760000000
0!
0%
#313765000000
1!
1%
#313770000000
0!
0%
#313775000000
1!
1%
#313780000000
0!
0%
#313785000000
1!
1%
#313790000000
0!
0%
#313795000000
1!
1%
#313800000000
0!
0%
#313805000000
1!
1%
#313810000000
0!
0%
#313815000000
1!
1%
#313820000000
0!
0%
#313825000000
1!
1%
#313830000000
0!
0%
#313835000000
1!
1%
#313840000000
0!
0%
#313845000000
1!
1%
#313850000000
0!
0%
#313855000000
1!
1%
#313860000000
0!
0%
#313865000000
1!
1%
#313870000000
0!
0%
#313875000000
1!
1%
#313880000000
0!
0%
#313885000000
1!
1%
#313890000000
0!
0%
#313895000000
1!
1%
#313900000000
0!
0%
#313905000000
1!
1%
#313910000000
0!
0%
#313915000000
1!
1%
#313920000000
0!
0%
#313925000000
1!
1%
#313930000000
0!
0%
#313935000000
1!
1%
#313940000000
0!
0%
#313945000000
1!
1%
#313950000000
0!
0%
#313955000000
1!
1%
#313960000000
0!
0%
#313965000000
1!
1%
#313970000000
0!
0%
#313975000000
1!
1%
#313980000000
0!
0%
#313985000000
1!
1%
#313990000000
0!
0%
#313995000000
1!
1%
#314000000000
0!
0%
#314005000000
1!
1%
#314010000000
0!
0%
#314015000000
1!
1%
#314020000000
0!
0%
#314025000000
1!
1%
#314030000000
0!
0%
#314035000000
1!
1%
#314040000000
0!
0%
#314045000000
1!
1%
#314050000000
0!
0%
#314055000000
1!
1%
#314060000000
0!
0%
#314065000000
1!
1%
#314070000000
0!
0%
#314075000000
1!
1%
#314080000000
0!
0%
#314085000000
1!
1%
#314090000000
0!
0%
#314095000000
1!
1%
#314100000000
0!
0%
#314105000000
1!
1%
#314110000000
0!
0%
#314115000000
1!
1%
#314120000000
0!
0%
#314125000000
1!
1%
#314130000000
0!
0%
#314135000000
1!
1%
#314140000000
0!
0%
#314145000000
1!
1%
#314150000000
0!
0%
#314155000000
1!
1%
#314160000000
0!
0%
#314165000000
1!
1%
#314170000000
0!
0%
#314175000000
1!
1%
#314180000000
0!
0%
#314185000000
1!
1%
#314190000000
0!
0%
#314195000000
1!
1%
#314200000000
0!
0%
#314205000000
1!
1%
#314210000000
0!
0%
#314215000000
1!
1%
#314220000000
0!
0%
#314225000000
1!
1%
#314230000000
0!
0%
#314235000000
1!
1%
#314240000000
0!
0%
#314245000000
1!
1%
#314250000000
0!
0%
#314255000000
1!
1%
#314260000000
0!
0%
#314265000000
1!
1%
#314270000000
0!
0%
#314275000000
1!
1%
#314280000000
0!
0%
#314285000000
1!
1%
#314290000000
0!
0%
#314295000000
1!
1%
#314300000000
0!
0%
#314305000000
1!
1%
#314310000000
0!
0%
#314315000000
1!
1%
#314320000000
0!
0%
#314325000000
1!
1%
#314330000000
0!
0%
#314335000000
1!
1%
#314340000000
0!
0%
#314345000000
1!
1%
#314350000000
0!
0%
#314355000000
1!
1%
#314360000000
0!
0%
#314365000000
1!
1%
#314370000000
0!
0%
#314375000000
1!
1%
#314380000000
0!
0%
#314385000000
1!
1%
#314390000000
0!
0%
#314395000000
1!
1%
#314400000000
0!
0%
#314405000000
1!
1%
#314410000000
0!
0%
#314415000000
1!
1%
#314420000000
0!
0%
#314425000000
1!
1%
#314430000000
0!
0%
#314435000000
1!
1%
#314440000000
0!
0%
#314445000000
1!
1%
#314450000000
0!
0%
#314455000000
1!
1%
#314460000000
0!
0%
#314465000000
1!
1%
#314470000000
0!
0%
#314475000000
1!
1%
#314480000000
0!
0%
#314485000000
1!
1%
#314490000000
0!
0%
#314495000000
1!
1%
#314500000000
0!
0%
#314505000000
1!
1%
#314510000000
0!
0%
#314515000000
1!
1%
#314520000000
0!
0%
#314525000000
1!
1%
#314530000000
0!
0%
#314535000000
1!
1%
#314540000000
0!
0%
#314545000000
1!
1%
#314550000000
0!
0%
#314555000000
1!
1%
#314560000000
0!
0%
#314565000000
1!
1%
#314570000000
0!
0%
#314575000000
1!
1%
#314580000000
0!
0%
#314585000000
1!
1%
#314590000000
0!
0%
#314595000000
1!
1%
#314600000000
0!
0%
#314605000000
1!
1%
#314610000000
0!
0%
#314615000000
1!
1%
#314620000000
0!
0%
#314625000000
1!
1%
#314630000000
0!
0%
#314635000000
1!
1%
#314640000000
0!
0%
#314645000000
1!
1%
#314650000000
0!
0%
#314655000000
1!
1%
#314660000000
0!
0%
#314665000000
1!
1%
#314670000000
0!
0%
#314675000000
1!
1%
#314680000000
0!
0%
#314685000000
1!
1%
#314690000000
0!
0%
#314695000000
1!
1%
#314700000000
0!
0%
#314705000000
1!
1%
#314710000000
0!
0%
#314715000000
1!
1%
#314720000000
0!
0%
#314725000000
1!
1%
#314730000000
0!
0%
#314735000000
1!
1%
#314740000000
0!
0%
#314745000000
1!
1%
#314750000000
0!
0%
#314755000000
1!
1%
#314760000000
0!
0%
#314765000000
1!
1%
#314770000000
0!
0%
#314775000000
1!
1%
#314780000000
0!
0%
#314785000000
1!
1%
#314790000000
0!
0%
#314795000000
1!
1%
#314800000000
0!
0%
#314805000000
1!
1%
#314810000000
0!
0%
#314815000000
1!
1%
#314820000000
0!
0%
#314825000000
1!
1%
#314830000000
0!
0%
#314835000000
1!
1%
#314840000000
0!
0%
#314845000000
1!
1%
#314850000000
0!
0%
#314855000000
1!
1%
#314860000000
0!
0%
#314865000000
1!
1%
#314870000000
0!
0%
#314875000000
1!
1%
#314880000000
0!
0%
#314885000000
1!
1%
#314890000000
0!
0%
#314895000000
1!
1%
#314900000000
0!
0%
#314905000000
1!
1%
#314910000000
0!
0%
#314915000000
1!
1%
#314920000000
0!
0%
#314925000000
1!
1%
#314930000000
0!
0%
#314935000000
1!
1%
#314940000000
0!
0%
#314945000000
1!
1%
#314950000000
0!
0%
#314955000000
1!
1%
#314960000000
0!
0%
#314965000000
1!
1%
#314970000000
0!
0%
#314975000000
1!
1%
#314980000000
0!
0%
#314985000000
1!
1%
#314990000000
0!
0%
#314995000000
1!
1%
#315000000000
0!
0%
#315005000000
1!
1%
#315010000000
0!
0%
#315015000000
1!
1%
#315020000000
0!
0%
#315025000000
1!
1%
#315030000000
0!
0%
#315035000000
1!
1%
#315040000000
0!
0%
#315045000000
1!
1%
#315050000000
0!
0%
#315055000000
1!
1%
#315060000000
0!
0%
#315065000000
1!
1%
#315070000000
0!
0%
#315075000000
1!
1%
#315080000000
0!
0%
#315085000000
1!
1%
#315090000000
0!
0%
#315095000000
1!
1%
#315100000000
0!
0%
#315105000000
1!
1%
#315110000000
0!
0%
#315115000000
1!
1%
#315120000000
0!
0%
#315125000000
1!
1%
#315130000000
0!
0%
#315135000000
1!
1%
#315140000000
0!
0%
#315145000000
1!
1%
#315150000000
0!
0%
#315155000000
1!
1%
#315160000000
0!
0%
#315165000000
1!
1%
#315170000000
0!
0%
#315175000000
1!
1%
#315180000000
0!
0%
#315185000000
1!
1%
#315190000000
0!
0%
#315195000000
1!
1%
#315200000000
0!
0%
#315205000000
1!
1%
#315210000000
0!
0%
#315215000000
1!
1%
#315220000000
0!
0%
#315225000000
1!
1%
#315230000000
0!
0%
#315235000000
1!
1%
#315240000000
0!
0%
#315245000000
1!
1%
#315250000000
0!
0%
#315255000000
1!
1%
#315260000000
0!
0%
#315265000000
1!
1%
#315270000000
0!
0%
#315275000000
1!
1%
#315280000000
0!
0%
#315285000000
1!
1%
#315290000000
0!
0%
#315295000000
1!
1%
#315300000000
0!
0%
#315305000000
1!
1%
#315310000000
0!
0%
#315315000000
1!
1%
#315320000000
0!
0%
#315325000000
1!
1%
#315330000000
0!
0%
#315335000000
1!
1%
#315340000000
0!
0%
#315345000000
1!
1%
#315350000000
0!
0%
#315355000000
1!
1%
#315360000000
0!
0%
#315365000000
1!
1%
#315370000000
0!
0%
#315375000000
1!
1%
#315380000000
0!
0%
#315385000000
1!
1%
#315390000000
0!
0%
#315395000000
1!
1%
#315400000000
0!
0%
#315405000000
1!
1%
#315410000000
0!
0%
#315415000000
1!
1%
#315420000000
0!
0%
#315425000000
1!
1%
#315430000000
0!
0%
#315435000000
1!
1%
#315440000000
0!
0%
#315445000000
1!
1%
#315450000000
0!
0%
#315455000000
1!
1%
#315460000000
0!
0%
#315465000000
1!
1%
#315470000000
0!
0%
#315475000000
1!
1%
#315480000000
0!
0%
#315485000000
1!
1%
#315490000000
0!
0%
#315495000000
1!
1%
#315500000000
0!
0%
#315505000000
1!
1%
#315510000000
0!
0%
#315515000000
1!
1%
#315520000000
0!
0%
#315525000000
1!
1%
#315530000000
0!
0%
#315535000000
1!
1%
#315540000000
0!
0%
#315545000000
1!
1%
#315550000000
0!
0%
#315555000000
1!
1%
#315560000000
0!
0%
#315565000000
1!
1%
#315570000000
0!
0%
#315575000000
1!
1%
#315580000000
0!
0%
#315585000000
1!
1%
#315590000000
0!
0%
#315595000000
1!
1%
#315600000000
0!
0%
#315605000000
1!
1%
#315610000000
0!
0%
#315615000000
1!
1%
#315620000000
0!
0%
#315625000000
1!
1%
#315630000000
0!
0%
#315635000000
1!
1%
#315640000000
0!
0%
#315645000000
1!
1%
#315650000000
0!
0%
#315655000000
1!
1%
#315660000000
0!
0%
#315665000000
1!
1%
#315670000000
0!
0%
#315675000000
1!
1%
#315680000000
0!
0%
#315685000000
1!
1%
#315690000000
0!
0%
#315695000000
1!
1%
#315700000000
0!
0%
#315705000000
1!
1%
#315710000000
0!
0%
#315715000000
1!
1%
#315720000000
0!
0%
#315725000000
1!
1%
#315730000000
0!
0%
#315735000000
1!
1%
#315740000000
0!
0%
#315745000000
1!
1%
#315750000000
0!
0%
#315755000000
1!
1%
#315760000000
0!
0%
#315765000000
1!
1%
#315770000000
0!
0%
#315775000000
1!
1%
#315780000000
0!
0%
#315785000000
1!
1%
#315790000000
0!
0%
#315795000000
1!
1%
#315800000000
0!
0%
#315805000000
1!
1%
#315810000000
0!
0%
#315815000000
1!
1%
#315820000000
0!
0%
#315825000000
1!
1%
#315830000000
0!
0%
#315835000000
1!
1%
#315840000000
0!
0%
#315845000000
1!
1%
#315850000000
0!
0%
#315855000000
1!
1%
#315860000000
0!
0%
#315865000000
1!
1%
#315870000000
0!
0%
#315875000000
1!
1%
#315880000000
0!
0%
#315885000000
1!
1%
#315890000000
0!
0%
#315895000000
1!
1%
#315900000000
0!
0%
#315905000000
1!
1%
#315910000000
0!
0%
#315915000000
1!
1%
#315920000000
0!
0%
#315925000000
1!
1%
#315930000000
0!
0%
#315935000000
1!
1%
#315940000000
0!
0%
#315945000000
1!
1%
#315950000000
0!
0%
#315955000000
1!
1%
#315960000000
0!
0%
#315965000000
1!
1%
#315970000000
0!
0%
#315975000000
1!
1%
#315980000000
0!
0%
#315985000000
1!
1%
#315990000000
0!
0%
#315995000000
1!
1%
#316000000000
0!
0%
#316005000000
1!
1%
#316010000000
0!
0%
#316015000000
1!
1%
#316020000000
0!
0%
#316025000000
1!
1%
#316030000000
0!
0%
#316035000000
1!
1%
#316040000000
0!
0%
#316045000000
1!
1%
#316050000000
0!
0%
#316055000000
1!
1%
#316060000000
0!
0%
#316065000000
1!
1%
#316070000000
0!
0%
#316075000000
1!
1%
#316080000000
0!
0%
#316085000000
1!
1%
#316090000000
0!
0%
#316095000000
1!
1%
#316100000000
0!
0%
#316105000000
1!
1%
#316110000000
0!
0%
#316115000000
1!
1%
#316120000000
0!
0%
#316125000000
1!
1%
#316130000000
0!
0%
#316135000000
1!
1%
#316140000000
0!
0%
#316145000000
1!
1%
#316150000000
0!
0%
#316155000000
1!
1%
#316160000000
0!
0%
#316165000000
1!
1%
#316170000000
0!
0%
#316175000000
1!
1%
#316180000000
0!
0%
#316185000000
1!
1%
#316190000000
0!
0%
#316195000000
1!
1%
#316200000000
0!
0%
#316205000000
1!
1%
#316210000000
0!
0%
#316215000000
1!
1%
#316220000000
0!
0%
#316225000000
1!
1%
#316230000000
0!
0%
#316235000000
1!
1%
#316240000000
0!
0%
#316245000000
1!
1%
#316250000000
0!
0%
#316255000000
1!
1%
#316260000000
0!
0%
#316265000000
1!
1%
#316270000000
0!
0%
#316275000000
1!
1%
#316280000000
0!
0%
#316285000000
1!
1%
#316290000000
0!
0%
#316295000000
1!
1%
#316300000000
0!
0%
#316305000000
1!
1%
#316310000000
0!
0%
#316315000000
1!
1%
#316320000000
0!
0%
#316325000000
1!
1%
#316330000000
0!
0%
#316335000000
1!
1%
#316340000000
0!
0%
#316345000000
1!
1%
#316350000000
0!
0%
#316355000000
1!
1%
#316360000000
0!
0%
#316365000000
1!
1%
#316370000000
0!
0%
#316375000000
1!
1%
#316380000000
0!
0%
#316385000000
1!
1%
#316390000000
0!
0%
#316395000000
1!
1%
#316400000000
0!
0%
#316405000000
1!
1%
#316410000000
0!
0%
#316415000000
1!
1%
#316420000000
0!
0%
#316425000000
1!
1%
#316430000000
0!
0%
#316435000000
1!
1%
#316440000000
0!
0%
#316445000000
1!
1%
#316450000000
0!
0%
#316455000000
1!
1%
#316460000000
0!
0%
#316465000000
1!
1%
#316470000000
0!
0%
#316475000000
1!
1%
#316480000000
0!
0%
#316485000000
1!
1%
#316490000000
0!
0%
#316495000000
1!
1%
#316500000000
0!
0%
#316505000000
1!
1%
#316510000000
0!
0%
#316515000000
1!
1%
#316520000000
0!
0%
#316525000000
1!
1%
#316530000000
0!
0%
#316535000000
1!
1%
#316540000000
0!
0%
#316545000000
1!
1%
#316550000000
0!
0%
#316555000000
1!
1%
#316560000000
0!
0%
#316565000000
1!
1%
#316570000000
0!
0%
#316575000000
1!
1%
#316580000000
0!
0%
#316585000000
1!
1%
#316590000000
0!
0%
#316595000000
1!
1%
#316600000000
0!
0%
#316605000000
1!
1%
#316610000000
0!
0%
#316615000000
1!
1%
#316620000000
0!
0%
#316625000000
1!
1%
#316630000000
0!
0%
#316635000000
1!
1%
#316640000000
0!
0%
#316645000000
1!
1%
#316650000000
0!
0%
#316655000000
1!
1%
#316660000000
0!
0%
#316665000000
1!
1%
#316670000000
0!
0%
#316675000000
1!
1%
#316680000000
0!
0%
#316685000000
1!
1%
#316690000000
0!
0%
#316695000000
1!
1%
#316700000000
0!
0%
#316705000000
1!
1%
#316710000000
0!
0%
#316715000000
1!
1%
#316720000000
0!
0%
#316725000000
1!
1%
#316730000000
0!
0%
#316735000000
1!
1%
#316740000000
0!
0%
#316745000000
1!
1%
#316750000000
0!
0%
#316755000000
1!
1%
#316760000000
0!
0%
#316765000000
1!
1%
#316770000000
0!
0%
#316775000000
1!
1%
#316780000000
0!
0%
#316785000000
1!
1%
#316790000000
0!
0%
#316795000000
1!
1%
#316800000000
0!
0%
#316805000000
1!
1%
#316810000000
0!
0%
#316815000000
1!
1%
#316820000000
0!
0%
#316825000000
1!
1%
#316830000000
0!
0%
#316835000000
1!
1%
#316840000000
0!
0%
#316845000000
1!
1%
#316850000000
0!
0%
#316855000000
1!
1%
#316860000000
0!
0%
#316865000000
1!
1%
#316870000000
0!
0%
#316875000000
1!
1%
#316880000000
0!
0%
#316885000000
1!
1%
#316890000000
0!
0%
#316895000000
1!
1%
#316900000000
0!
0%
#316905000000
1!
1%
#316910000000
0!
0%
#316915000000
1!
1%
#316920000000
0!
0%
#316925000000
1!
1%
#316930000000
0!
0%
#316935000000
1!
1%
#316940000000
0!
0%
#316945000000
1!
1%
#316950000000
0!
0%
#316955000000
1!
1%
#316960000000
0!
0%
#316965000000
1!
1%
#316970000000
0!
0%
#316975000000
1!
1%
#316980000000
0!
0%
#316985000000
1!
1%
#316990000000
0!
0%
#316995000000
1!
1%
#317000000000
0!
0%
#317005000000
1!
1%
#317010000000
0!
0%
#317015000000
1!
1%
#317020000000
0!
0%
#317025000000
1!
1%
#317030000000
0!
0%
#317035000000
1!
1%
#317040000000
0!
0%
#317045000000
1!
1%
#317050000000
0!
0%
#317055000000
1!
1%
#317060000000
0!
0%
#317065000000
1!
1%
#317070000000
0!
0%
#317075000000
1!
1%
#317080000000
0!
0%
#317085000000
1!
1%
#317090000000
0!
0%
#317095000000
1!
1%
#317100000000
0!
0%
#317105000000
1!
1%
#317110000000
0!
0%
#317115000000
1!
1%
#317120000000
0!
0%
#317125000000
1!
1%
#317130000000
0!
0%
#317135000000
1!
1%
#317140000000
0!
0%
#317145000000
1!
1%
#317150000000
0!
0%
#317155000000
1!
1%
#317160000000
0!
0%
#317165000000
1!
1%
#317170000000
0!
0%
#317175000000
1!
1%
#317180000000
0!
0%
#317185000000
1!
1%
#317190000000
0!
0%
#317195000000
1!
1%
#317200000000
0!
0%
#317205000000
1!
1%
#317210000000
0!
0%
#317215000000
1!
1%
#317220000000
0!
0%
#317225000000
1!
1%
#317230000000
0!
0%
#317235000000
1!
1%
#317240000000
0!
0%
#317245000000
1!
1%
#317250000000
0!
0%
#317255000000
1!
1%
#317260000000
0!
0%
#317265000000
1!
1%
#317270000000
0!
0%
#317275000000
1!
1%
#317280000000
0!
0%
#317285000000
1!
1%
#317290000000
0!
0%
#317295000000
1!
1%
#317300000000
0!
0%
#317305000000
1!
1%
#317310000000
0!
0%
#317315000000
1!
1%
#317320000000
0!
0%
#317325000000
1!
1%
#317330000000
0!
0%
#317335000000
1!
1%
#317340000000
0!
0%
#317345000000
1!
1%
#317350000000
0!
0%
#317355000000
1!
1%
#317360000000
0!
0%
#317365000000
1!
1%
#317370000000
0!
0%
#317375000000
1!
1%
#317380000000
0!
0%
#317385000000
1!
1%
#317390000000
0!
0%
#317395000000
1!
1%
#317400000000
0!
0%
#317405000000
1!
1%
#317410000000
0!
0%
#317415000000
1!
1%
#317420000000
0!
0%
#317425000000
1!
1%
#317430000000
0!
0%
#317435000000
1!
1%
#317440000000
0!
0%
#317445000000
1!
1%
#317450000000
0!
0%
#317455000000
1!
1%
#317460000000
0!
0%
#317465000000
1!
1%
#317470000000
0!
0%
#317475000000
1!
1%
#317480000000
0!
0%
#317485000000
1!
1%
#317490000000
0!
0%
#317495000000
1!
1%
#317500000000
0!
0%
#317505000000
1!
1%
#317510000000
0!
0%
#317515000000
1!
1%
#317520000000
0!
0%
#317525000000
1!
1%
#317530000000
0!
0%
#317535000000
1!
1%
#317540000000
0!
0%
#317545000000
1!
1%
#317550000000
0!
0%
#317555000000
1!
1%
#317560000000
0!
0%
#317565000000
1!
1%
#317570000000
0!
0%
#317575000000
1!
1%
#317580000000
0!
0%
#317585000000
1!
1%
#317590000000
0!
0%
#317595000000
1!
1%
#317600000000
0!
0%
#317605000000
1!
1%
#317610000000
0!
0%
#317615000000
1!
1%
#317620000000
0!
0%
#317625000000
1!
1%
#317630000000
0!
0%
#317635000000
1!
1%
#317640000000
0!
0%
#317645000000
1!
1%
#317650000000
0!
0%
#317655000000
1!
1%
#317660000000
0!
0%
#317665000000
1!
1%
#317670000000
0!
0%
#317675000000
1!
1%
#317680000000
0!
0%
#317685000000
1!
1%
#317690000000
0!
0%
#317695000000
1!
1%
#317700000000
0!
0%
#317705000000
1!
1%
#317710000000
0!
0%
#317715000000
1!
1%
#317720000000
0!
0%
#317725000000
1!
1%
#317730000000
0!
0%
#317735000000
1!
1%
#317740000000
0!
0%
#317745000000
1!
1%
#317750000000
0!
0%
#317755000000
1!
1%
#317760000000
0!
0%
#317765000000
1!
1%
#317770000000
0!
0%
#317775000000
1!
1%
#317780000000
0!
0%
#317785000000
1!
1%
#317790000000
0!
0%
#317795000000
1!
1%
#317800000000
0!
0%
#317805000000
1!
1%
#317810000000
0!
0%
#317815000000
1!
1%
#317820000000
0!
0%
#317825000000
1!
1%
#317830000000
0!
0%
#317835000000
1!
1%
#317840000000
0!
0%
#317845000000
1!
1%
#317850000000
0!
0%
#317855000000
1!
1%
#317860000000
0!
0%
#317865000000
1!
1%
#317870000000
0!
0%
#317875000000
1!
1%
#317880000000
0!
0%
#317885000000
1!
1%
#317890000000
0!
0%
#317895000000
1!
1%
#317900000000
0!
0%
#317905000000
1!
1%
#317910000000
0!
0%
#317915000000
1!
1%
#317920000000
0!
0%
#317925000000
1!
1%
#317930000000
0!
0%
#317935000000
1!
1%
#317940000000
0!
0%
#317945000000
1!
1%
#317950000000
0!
0%
#317955000000
1!
1%
#317960000000
0!
0%
#317965000000
1!
1%
#317970000000
0!
0%
#317975000000
1!
1%
#317980000000
0!
0%
#317985000000
1!
1%
#317990000000
0!
0%
#317995000000
1!
1%
#318000000000
0!
0%
#318005000000
1!
1%
#318010000000
0!
0%
#318015000000
1!
1%
#318020000000
0!
0%
#318025000000
1!
1%
#318030000000
0!
0%
#318035000000
1!
1%
#318040000000
0!
0%
#318045000000
1!
1%
#318050000000
0!
0%
#318055000000
1!
1%
#318060000000
0!
0%
#318065000000
1!
1%
#318070000000
0!
0%
#318075000000
1!
1%
#318080000000
0!
0%
#318085000000
1!
1%
#318090000000
0!
0%
#318095000000
1!
1%
#318100000000
0!
0%
#318105000000
1!
1%
#318110000000
0!
0%
#318115000000
1!
1%
#318120000000
0!
0%
#318125000000
1!
1%
#318130000000
0!
0%
#318135000000
1!
1%
#318140000000
0!
0%
#318145000000
1!
1%
#318150000000
0!
0%
#318155000000
1!
1%
#318160000000
0!
0%
#318165000000
1!
1%
#318170000000
0!
0%
#318175000000
1!
1%
#318180000000
0!
0%
#318185000000
1!
1%
#318190000000
0!
0%
#318195000000
1!
1%
#318200000000
0!
0%
#318205000000
1!
1%
#318210000000
0!
0%
#318215000000
1!
1%
#318220000000
0!
0%
#318225000000
1!
1%
#318230000000
0!
0%
#318235000000
1!
1%
#318240000000
0!
0%
#318245000000
1!
1%
#318250000000
0!
0%
#318255000000
1!
1%
#318260000000
0!
0%
#318265000000
1!
1%
#318270000000
0!
0%
#318275000000
1!
1%
#318280000000
0!
0%
#318285000000
1!
1%
#318290000000
0!
0%
#318295000000
1!
1%
#318300000000
0!
0%
#318305000000
1!
1%
#318310000000
0!
0%
#318315000000
1!
1%
#318320000000
0!
0%
#318325000000
1!
1%
#318330000000
0!
0%
#318335000000
1!
1%
#318340000000
0!
0%
#318345000000
1!
1%
#318350000000
0!
0%
#318355000000
1!
1%
#318360000000
0!
0%
#318365000000
1!
1%
#318370000000
0!
0%
#318375000000
1!
1%
#318380000000
0!
0%
#318385000000
1!
1%
#318390000000
0!
0%
#318395000000
1!
1%
#318400000000
0!
0%
#318405000000
1!
1%
#318410000000
0!
0%
#318415000000
1!
1%
#318420000000
0!
0%
#318425000000
1!
1%
#318430000000
0!
0%
#318435000000
1!
1%
#318440000000
0!
0%
#318445000000
1!
1%
#318450000000
0!
0%
#318455000000
1!
1%
#318460000000
0!
0%
#318465000000
1!
1%
#318470000000
0!
0%
#318475000000
1!
1%
#318480000000
0!
0%
#318485000000
1!
1%
#318490000000
0!
0%
#318495000000
1!
1%
#318500000000
0!
0%
#318505000000
1!
1%
#318510000000
0!
0%
#318515000000
1!
1%
#318520000000
0!
0%
#318525000000
1!
1%
#318530000000
0!
0%
#318535000000
1!
1%
#318540000000
0!
0%
#318545000000
1!
1%
#318550000000
0!
0%
#318555000000
1!
1%
#318560000000
0!
0%
#318565000000
1!
1%
#318570000000
0!
0%
#318575000000
1!
1%
#318580000000
0!
0%
#318585000000
1!
1%
#318590000000
0!
0%
#318595000000
1!
1%
#318600000000
0!
0%
#318605000000
1!
1%
#318610000000
0!
0%
#318615000000
1!
1%
#318620000000
0!
0%
#318625000000
1!
1%
#318630000000
0!
0%
#318635000000
1!
1%
#318640000000
0!
0%
#318645000000
1!
1%
#318650000000
0!
0%
#318655000000
1!
1%
#318660000000
0!
0%
#318665000000
1!
1%
#318670000000
0!
0%
#318675000000
1!
1%
#318680000000
0!
0%
#318685000000
1!
1%
#318690000000
0!
0%
#318695000000
1!
1%
#318700000000
0!
0%
#318705000000
1!
1%
#318710000000
0!
0%
#318715000000
1!
1%
#318720000000
0!
0%
#318725000000
1!
1%
#318730000000
0!
0%
#318735000000
1!
1%
#318740000000
0!
0%
#318745000000
1!
1%
#318750000000
0!
0%
#318755000000
1!
1%
#318760000000
0!
0%
#318765000000
1!
1%
#318770000000
0!
0%
#318775000000
1!
1%
#318780000000
0!
0%
#318785000000
1!
1%
#318790000000
0!
0%
#318795000000
1!
1%
#318800000000
0!
0%
#318805000000
1!
1%
#318810000000
0!
0%
#318815000000
1!
1%
#318820000000
0!
0%
#318825000000
1!
1%
#318830000000
0!
0%
#318835000000
1!
1%
#318840000000
0!
0%
#318845000000
1!
1%
#318850000000
0!
0%
#318855000000
1!
1%
#318860000000
0!
0%
#318865000000
1!
1%
#318870000000
0!
0%
#318875000000
1!
1%
#318880000000
0!
0%
#318885000000
1!
1%
#318890000000
0!
0%
#318895000000
1!
1%
#318900000000
0!
0%
#318905000000
1!
1%
#318910000000
0!
0%
#318915000000
1!
1%
#318920000000
0!
0%
#318925000000
1!
1%
#318930000000
0!
0%
#318935000000
1!
1%
#318940000000
0!
0%
#318945000000
1!
1%
#318950000000
0!
0%
#318955000000
1!
1%
#318960000000
0!
0%
#318965000000
1!
1%
#318970000000
0!
0%
#318975000000
1!
1%
#318980000000
0!
0%
#318985000000
1!
1%
#318990000000
0!
0%
#318995000000
1!
1%
#319000000000
0!
0%
#319005000000
1!
1%
#319010000000
0!
0%
#319015000000
1!
1%
#319020000000
0!
0%
#319025000000
1!
1%
#319030000000
0!
0%
#319035000000
1!
1%
#319040000000
0!
0%
#319045000000
1!
1%
#319050000000
0!
0%
#319055000000
1!
1%
#319060000000
0!
0%
#319065000000
1!
1%
#319070000000
0!
0%
#319075000000
1!
1%
#319080000000
0!
0%
#319085000000
1!
1%
#319090000000
0!
0%
#319095000000
1!
1%
#319100000000
0!
0%
#319105000000
1!
1%
#319110000000
0!
0%
#319115000000
1!
1%
#319120000000
0!
0%
#319125000000
1!
1%
#319130000000
0!
0%
#319135000000
1!
1%
#319140000000
0!
0%
#319145000000
1!
1%
#319150000000
0!
0%
#319155000000
1!
1%
#319160000000
0!
0%
#319165000000
1!
1%
#319170000000
0!
0%
#319175000000
1!
1%
#319180000000
0!
0%
#319185000000
1!
1%
#319190000000
0!
0%
#319195000000
1!
1%
#319200000000
0!
0%
#319205000000
1!
1%
#319210000000
0!
0%
#319215000000
1!
1%
#319220000000
0!
0%
#319225000000
1!
1%
#319230000000
0!
0%
#319235000000
1!
1%
#319240000000
0!
0%
#319245000000
1!
1%
#319250000000
0!
0%
#319255000000
1!
1%
#319260000000
0!
0%
#319265000000
1!
1%
#319270000000
0!
0%
#319275000000
1!
1%
#319280000000
0!
0%
#319285000000
1!
1%
#319290000000
0!
0%
#319295000000
1!
1%
#319300000000
0!
0%
#319305000000
1!
1%
#319310000000
0!
0%
#319315000000
1!
1%
#319320000000
0!
0%
#319325000000
1!
1%
#319330000000
0!
0%
#319335000000
1!
1%
#319340000000
0!
0%
#319345000000
1!
1%
#319350000000
0!
0%
#319355000000
1!
1%
#319360000000
0!
0%
#319365000000
1!
1%
#319370000000
0!
0%
#319375000000
1!
1%
#319380000000
0!
0%
#319385000000
1!
1%
#319390000000
0!
0%
#319395000000
1!
1%
#319400000000
0!
0%
#319405000000
1!
1%
#319410000000
0!
0%
#319415000000
1!
1%
#319420000000
0!
0%
#319425000000
1!
1%
#319430000000
0!
0%
#319435000000
1!
1%
#319440000000
0!
0%
#319445000000
1!
1%
#319450000000
0!
0%
#319455000000
1!
1%
#319460000000
0!
0%
#319465000000
1!
1%
#319470000000
0!
0%
#319475000000
1!
1%
#319480000000
0!
0%
#319485000000
1!
1%
#319490000000
0!
0%
#319495000000
1!
1%
#319500000000
0!
0%
#319505000000
1!
1%
#319510000000
0!
0%
#319515000000
1!
1%
#319520000000
0!
0%
#319525000000
1!
1%
#319530000000
0!
0%
#319535000000
1!
1%
#319540000000
0!
0%
#319545000000
1!
1%
#319550000000
0!
0%
#319555000000
1!
1%
#319560000000
0!
0%
#319565000000
1!
1%
#319570000000
0!
0%
#319575000000
1!
1%
#319580000000
0!
0%
#319585000000
1!
1%
#319590000000
0!
0%
#319595000000
1!
1%
#319600000000
0!
0%
#319605000000
1!
1%
#319610000000
0!
0%
#319615000000
1!
1%
#319620000000
0!
0%
#319625000000
1!
1%
#319630000000
0!
0%
#319635000000
1!
1%
#319640000000
0!
0%
#319645000000
1!
1%
#319650000000
0!
0%
#319655000000
1!
1%
#319660000000
0!
0%
#319665000000
1!
1%
#319670000000
0!
0%
#319675000000
1!
1%
#319680000000
0!
0%
#319685000000
1!
1%
#319690000000
0!
0%
#319695000000
1!
1%
#319700000000
0!
0%
#319705000000
1!
1%
#319710000000
0!
0%
#319715000000
1!
1%
#319720000000
0!
0%
#319725000000
1!
1%
#319730000000
0!
0%
#319735000000
1!
1%
#319740000000
0!
0%
#319745000000
1!
1%
#319750000000
0!
0%
#319755000000
1!
1%
#319760000000
0!
0%
#319765000000
1!
1%
#319770000000
0!
0%
#319775000000
1!
1%
#319780000000
0!
0%
#319785000000
1!
1%
#319790000000
0!
0%
#319795000000
1!
1%
#319800000000
0!
0%
#319805000000
1!
1%
#319810000000
0!
0%
#319815000000
1!
1%
#319820000000
0!
0%
#319825000000
1!
1%
#319830000000
0!
0%
#319835000000
1!
1%
#319840000000
0!
0%
#319845000000
1!
1%
#319850000000
0!
0%
#319855000000
1!
1%
#319860000000
0!
0%
#319865000000
1!
1%
#319870000000
0!
0%
#319875000000
1!
1%
#319880000000
0!
0%
#319885000000
1!
1%
#319890000000
0!
0%
#319895000000
1!
1%
#319900000000
0!
0%
#319905000000
1!
1%
#319910000000
0!
0%
#319915000000
1!
1%
#319920000000
0!
0%
#319925000000
1!
1%
#319930000000
0!
0%
#319935000000
1!
1%
#319940000000
0!
0%
#319945000000
1!
1%
#319950000000
0!
0%
#319955000000
1!
1%
#319960000000
0!
0%
#319965000000
1!
1%
#319970000000
0!
0%
#319975000000
1!
1%
#319980000000
0!
0%
#319985000000
1!
1%
#319990000000
0!
0%
#319995000000
1!
1%
#320000000000
0!
0%
#320005000000
1!
1%
#320010000000
0!
0%
#320015000000
1!
1%
#320020000000
0!
0%
#320025000000
1!
1%
#320030000000
0!
0%
#320035000000
1!
1%
#320040000000
0!
0%
#320045000000
1!
1%
#320050000000
0!
0%
#320055000000
1!
1%
#320060000000
0!
0%
#320065000000
1!
1%
#320070000000
0!
0%
#320075000000
1!
1%
#320080000000
0!
0%
#320085000000
1!
1%
#320090000000
0!
0%
#320095000000
1!
1%
#320100000000
0!
0%
#320105000000
1!
1%
#320110000000
0!
0%
#320115000000
1!
1%
#320120000000
0!
0%
#320125000000
1!
1%
#320130000000
0!
0%
#320135000000
1!
1%
#320140000000
0!
0%
#320145000000
1!
1%
#320150000000
0!
0%
#320155000000
1!
1%
#320160000000
0!
0%
#320165000000
1!
1%
#320170000000
0!
0%
#320175000000
1!
1%
#320180000000
0!
0%
#320185000000
1!
1%
#320190000000
0!
0%
#320195000000
1!
1%
#320200000000
0!
0%
#320205000000
1!
1%
#320210000000
0!
0%
#320215000000
1!
1%
#320220000000
0!
0%
#320225000000
1!
1%
#320230000000
0!
0%
#320235000000
1!
1%
#320240000000
0!
0%
#320245000000
1!
1%
#320250000000
0!
0%
#320255000000
1!
1%
#320260000000
0!
0%
#320265000000
1!
1%
#320270000000
0!
0%
#320275000000
1!
1%
#320280000000
0!
0%
#320285000000
1!
1%
#320290000000
0!
0%
#320295000000
1!
1%
#320300000000
0!
0%
#320305000000
1!
1%
#320310000000
0!
0%
#320315000000
1!
1%
#320320000000
0!
0%
#320325000000
1!
1%
#320330000000
0!
0%
#320335000000
1!
1%
#320340000000
0!
0%
#320345000000
1!
1%
#320350000000
0!
0%
#320355000000
1!
1%
#320360000000
0!
0%
#320365000000
1!
1%
#320370000000
0!
0%
#320375000000
1!
1%
#320380000000
0!
0%
#320385000000
1!
1%
#320390000000
0!
0%
#320395000000
1!
1%
#320400000000
0!
0%
#320405000000
1!
1%
#320410000000
0!
0%
#320415000000
1!
1%
#320420000000
0!
0%
#320425000000
1!
1%
#320430000000
0!
0%
#320435000000
1!
1%
#320440000000
0!
0%
#320445000000
1!
1%
#320450000000
0!
0%
#320455000000
1!
1%
#320460000000
0!
0%
#320465000000
1!
1%
#320470000000
0!
0%
#320475000000
1!
1%
#320480000000
0!
0%
#320485000000
1!
1%
#320490000000
0!
0%
#320495000000
1!
1%
#320500000000
0!
0%
#320505000000
1!
1%
#320510000000
0!
0%
#320515000000
1!
1%
#320520000000
0!
0%
#320525000000
1!
1%
#320530000000
0!
0%
#320535000000
1!
1%
#320540000000
0!
0%
#320545000000
1!
1%
#320550000000
0!
0%
#320555000000
1!
1%
#320560000000
0!
0%
#320565000000
1!
1%
#320570000000
0!
0%
#320575000000
1!
1%
#320580000000
0!
0%
#320585000000
1!
1%
#320590000000
0!
0%
#320595000000
1!
1%
#320600000000
0!
0%
#320605000000
1!
1%
#320610000000
0!
0%
#320615000000
1!
1%
#320620000000
0!
0%
#320625000000
1!
1%
#320630000000
0!
0%
#320635000000
1!
1%
#320640000000
0!
0%
#320645000000
1!
1%
#320650000000
0!
0%
#320655000000
1!
1%
#320660000000
0!
0%
#320665000000
1!
1%
#320670000000
0!
0%
#320675000000
1!
1%
#320680000000
0!
0%
#320685000000
1!
1%
#320690000000
0!
0%
#320695000000
1!
1%
#320700000000
0!
0%
#320705000000
1!
1%
#320710000000
0!
0%
#320715000000
1!
1%
#320720000000
0!
0%
#320725000000
1!
1%
#320730000000
0!
0%
#320735000000
1!
1%
#320740000000
0!
0%
#320745000000
1!
1%
#320750000000
0!
0%
#320755000000
1!
1%
#320760000000
0!
0%
#320765000000
1!
1%
#320770000000
0!
0%
#320775000000
1!
1%
#320780000000
0!
0%
#320785000000
1!
1%
#320790000000
0!
0%
#320795000000
1!
1%
#320800000000
0!
0%
#320805000000
1!
1%
#320810000000
0!
0%
#320815000000
1!
1%
#320820000000
0!
0%
#320825000000
1!
1%
#320830000000
0!
0%
#320835000000
1!
1%
#320840000000
0!
0%
#320845000000
1!
1%
#320850000000
0!
0%
#320855000000
1!
1%
#320860000000
0!
0%
#320865000000
1!
1%
#320870000000
0!
0%
#320875000000
1!
1%
#320880000000
0!
0%
#320885000000
1!
1%
#320890000000
0!
0%
#320895000000
1!
1%
#320900000000
0!
0%
#320905000000
1!
1%
#320910000000
0!
0%
#320915000000
1!
1%
#320920000000
0!
0%
#320925000000
1!
1%
#320930000000
0!
0%
#320935000000
1!
1%
#320940000000
0!
0%
#320945000000
1!
1%
#320950000000
0!
0%
#320955000000
1!
1%
#320960000000
0!
0%
#320965000000
1!
1%
#320970000000
0!
0%
#320975000000
1!
1%
#320980000000
0!
0%
#320985000000
1!
1%
#320990000000
0!
0%
#320995000000
1!
1%
#321000000000
0!
0%
#321005000000
1!
1%
#321010000000
0!
0%
#321015000000
1!
1%
#321020000000
0!
0%
#321025000000
1!
1%
#321030000000
0!
0%
#321035000000
1!
1%
#321040000000
0!
0%
#321045000000
1!
1%
#321050000000
0!
0%
#321055000000
1!
1%
#321060000000
0!
0%
#321065000000
1!
1%
#321070000000
0!
0%
#321075000000
1!
1%
#321080000000
0!
0%
#321085000000
1!
1%
#321090000000
0!
0%
#321095000000
1!
1%
#321100000000
0!
0%
#321105000000
1!
1%
#321110000000
0!
0%
#321115000000
1!
1%
#321120000000
0!
0%
#321125000000
1!
1%
#321130000000
0!
0%
#321135000000
1!
1%
#321140000000
0!
0%
#321145000000
1!
1%
#321150000000
0!
0%
#321155000000
1!
1%
#321160000000
0!
0%
#321165000000
1!
1%
#321170000000
0!
0%
#321175000000
1!
1%
#321180000000
0!
0%
#321185000000
1!
1%
#321190000000
0!
0%
#321195000000
1!
1%
#321200000000
0!
0%
#321205000000
1!
1%
#321210000000
0!
0%
#321215000000
1!
1%
#321220000000
0!
0%
#321225000000
1!
1%
#321230000000
0!
0%
#321235000000
1!
1%
#321240000000
0!
0%
#321245000000
1!
1%
#321250000000
0!
0%
#321255000000
1!
1%
#321260000000
0!
0%
#321265000000
1!
1%
#321270000000
0!
0%
#321275000000
1!
1%
#321280000000
0!
0%
#321285000000
1!
1%
#321290000000
0!
0%
#321295000000
1!
1%
#321300000000
0!
0%
#321305000000
1!
1%
#321310000000
0!
0%
#321315000000
1!
1%
#321320000000
0!
0%
#321325000000
1!
1%
#321330000000
0!
0%
#321335000000
1!
1%
#321340000000
0!
0%
#321345000000
1!
1%
#321350000000
0!
0%
#321355000000
1!
1%
#321360000000
0!
0%
#321365000000
1!
1%
#321370000000
0!
0%
#321375000000
1!
1%
#321380000000
0!
0%
#321385000000
1!
1%
#321390000000
0!
0%
#321395000000
1!
1%
#321400000000
0!
0%
#321405000000
1!
1%
#321410000000
0!
0%
#321415000000
1!
1%
#321420000000
0!
0%
#321425000000
1!
1%
#321430000000
0!
0%
#321435000000
1!
1%
#321440000000
0!
0%
#321445000000
1!
1%
#321450000000
0!
0%
#321455000000
1!
1%
#321460000000
0!
0%
#321465000000
1!
1%
#321470000000
0!
0%
#321475000000
1!
1%
#321480000000
0!
0%
#321485000000
1!
1%
#321490000000
0!
0%
#321495000000
1!
1%
#321500000000
0!
0%
#321505000000
1!
1%
#321510000000
0!
0%
#321515000000
1!
1%
#321520000000
0!
0%
#321525000000
1!
1%
#321530000000
0!
0%
#321535000000
1!
1%
#321540000000
0!
0%
#321545000000
1!
1%
#321550000000
0!
0%
#321555000000
1!
1%
#321560000000
0!
0%
#321565000000
1!
1%
#321570000000
0!
0%
#321575000000
1!
1%
#321580000000
0!
0%
#321585000000
1!
1%
#321590000000
0!
0%
#321595000000
1!
1%
#321600000000
0!
0%
#321605000000
1!
1%
#321610000000
0!
0%
#321615000000
1!
1%
#321620000000
0!
0%
#321625000000
1!
1%
#321630000000
0!
0%
#321635000000
1!
1%
#321640000000
0!
0%
#321645000000
1!
1%
#321650000000
0!
0%
#321655000000
1!
1%
#321660000000
0!
0%
#321665000000
1!
1%
#321670000000
0!
0%
#321675000000
1!
1%
#321680000000
0!
0%
#321685000000
1!
1%
#321690000000
0!
0%
#321695000000
1!
1%
#321700000000
0!
0%
#321705000000
1!
1%
#321710000000
0!
0%
#321715000000
1!
1%
#321720000000
0!
0%
#321725000000
1!
1%
#321730000000
0!
0%
#321735000000
1!
1%
#321740000000
0!
0%
#321745000000
1!
1%
#321750000000
0!
0%
#321755000000
1!
1%
#321760000000
0!
0%
#321765000000
1!
1%
#321770000000
0!
0%
#321775000000
1!
1%
#321780000000
0!
0%
#321785000000
1!
1%
#321790000000
0!
0%
#321795000000
1!
1%
#321800000000
0!
0%
#321805000000
1!
1%
#321810000000
0!
0%
#321815000000
1!
1%
#321820000000
0!
0%
#321825000000
1!
1%
#321830000000
0!
0%
#321835000000
1!
1%
#321840000000
0!
0%
#321845000000
1!
1%
#321850000000
0!
0%
#321855000000
1!
1%
#321860000000
0!
0%
#321865000000
1!
1%
#321870000000
0!
0%
#321875000000
1!
1%
#321880000000
0!
0%
#321885000000
1!
1%
#321890000000
0!
0%
#321895000000
1!
1%
#321900000000
0!
0%
#321905000000
1!
1%
#321910000000
0!
0%
#321915000000
1!
1%
#321920000000
0!
0%
#321925000000
1!
1%
#321930000000
0!
0%
#321935000000
1!
1%
#321940000000
0!
0%
#321945000000
1!
1%
#321950000000
0!
0%
#321955000000
1!
1%
#321960000000
0!
0%
#321965000000
1!
1%
#321970000000
0!
0%
#321975000000
1!
1%
#321980000000
0!
0%
#321985000000
1!
1%
#321990000000
0!
0%
#321995000000
1!
1%
#322000000000
0!
0%
#322005000000
1!
1%
#322010000000
0!
0%
#322015000000
1!
1%
#322020000000
0!
0%
#322025000000
1!
1%
#322030000000
0!
0%
#322035000000
1!
1%
#322040000000
0!
0%
#322045000000
1!
1%
#322050000000
0!
0%
#322055000000
1!
1%
#322060000000
0!
0%
#322065000000
1!
1%
#322070000000
0!
0%
#322075000000
1!
1%
#322080000000
0!
0%
#322085000000
1!
1%
#322090000000
0!
0%
#322095000000
1!
1%
#322100000000
0!
0%
#322105000000
1!
1%
#322110000000
0!
0%
#322115000000
1!
1%
#322120000000
0!
0%
#322125000000
1!
1%
#322130000000
0!
0%
#322135000000
1!
1%
#322140000000
0!
0%
#322145000000
1!
1%
#322150000000
0!
0%
#322155000000
1!
1%
#322160000000
0!
0%
#322165000000
1!
1%
#322170000000
0!
0%
#322175000000
1!
1%
#322180000000
0!
0%
#322185000000
1!
1%
#322190000000
0!
0%
#322195000000
1!
1%
#322200000000
0!
0%
#322205000000
1!
1%
#322210000000
0!
0%
#322215000000
1!
1%
#322220000000
0!
0%
#322225000000
1!
1%
#322230000000
0!
0%
#322235000000
1!
1%
#322240000000
0!
0%
#322245000000
1!
1%
#322250000000
0!
0%
#322255000000
1!
1%
#322260000000
0!
0%
#322265000000
1!
1%
#322270000000
0!
0%
#322275000000
1!
1%
#322280000000
0!
0%
#322285000000
1!
1%
#322290000000
0!
0%
#322295000000
1!
1%
#322300000000
0!
0%
#322305000000
1!
1%
#322310000000
0!
0%
#322315000000
1!
1%
#322320000000
0!
0%
#322325000000
1!
1%
#322330000000
0!
0%
#322335000000
1!
1%
#322340000000
0!
0%
#322345000000
1!
1%
#322350000000
0!
0%
#322355000000
1!
1%
#322360000000
0!
0%
#322365000000
1!
1%
#322370000000
0!
0%
#322375000000
1!
1%
#322380000000
0!
0%
#322385000000
1!
1%
#322390000000
0!
0%
#322395000000
1!
1%
#322400000000
0!
0%
#322405000000
1!
1%
#322410000000
0!
0%
#322415000000
1!
1%
#322420000000
0!
0%
#322425000000
1!
1%
#322430000000
0!
0%
#322435000000
1!
1%
#322440000000
0!
0%
#322445000000
1!
1%
#322450000000
0!
0%
#322455000000
1!
1%
#322460000000
0!
0%
#322465000000
1!
1%
#322470000000
0!
0%
#322475000000
1!
1%
#322480000000
0!
0%
#322485000000
1!
1%
#322490000000
0!
0%
#322495000000
1!
1%
#322500000000
0!
0%
#322505000000
1!
1%
#322510000000
0!
0%
#322515000000
1!
1%
#322520000000
0!
0%
#322525000000
1!
1%
#322530000000
0!
0%
#322535000000
1!
1%
#322540000000
0!
0%
#322545000000
1!
1%
#322550000000
0!
0%
#322555000000
1!
1%
#322560000000
0!
0%
#322565000000
1!
1%
#322570000000
0!
0%
#322575000000
1!
1%
#322580000000
0!
0%
#322585000000
1!
1%
#322590000000
0!
0%
#322595000000
1!
1%
#322600000000
0!
0%
#322605000000
1!
1%
#322610000000
0!
0%
#322615000000
1!
1%
#322620000000
0!
0%
#322625000000
1!
1%
#322630000000
0!
0%
#322635000000
1!
1%
#322640000000
0!
0%
#322645000000
1!
1%
#322650000000
0!
0%
#322655000000
1!
1%
#322660000000
0!
0%
#322665000000
1!
1%
#322670000000
0!
0%
#322675000000
1!
1%
#322680000000
0!
0%
#322685000000
1!
1%
#322690000000
0!
0%
#322695000000
1!
1%
#322700000000
0!
0%
#322705000000
1!
1%
#322710000000
0!
0%
#322715000000
1!
1%
#322720000000
0!
0%
#322725000000
1!
1%
#322730000000
0!
0%
#322735000000
1!
1%
#322740000000
0!
0%
#322745000000
1!
1%
#322750000000
0!
0%
#322755000000
1!
1%
#322760000000
0!
0%
#322765000000
1!
1%
#322770000000
0!
0%
#322775000000
1!
1%
#322780000000
0!
0%
#322785000000
1!
1%
#322790000000
0!
0%
#322795000000
1!
1%
#322800000000
0!
0%
#322805000000
1!
1%
#322810000000
0!
0%
#322815000000
1!
1%
#322820000000
0!
0%
#322825000000
1!
1%
#322830000000
0!
0%
#322835000000
1!
1%
#322840000000
0!
0%
#322845000000
1!
1%
#322850000000
0!
0%
#322855000000
1!
1%
#322860000000
0!
0%
#322865000000
1!
1%
#322870000000
0!
0%
#322875000000
1!
1%
#322880000000
0!
0%
#322885000000
1!
1%
#322890000000
0!
0%
#322895000000
1!
1%
#322900000000
0!
0%
#322905000000
1!
1%
#322910000000
0!
0%
#322915000000
1!
1%
#322920000000
0!
0%
#322925000000
1!
1%
#322930000000
0!
0%
#322935000000
1!
1%
#322940000000
0!
0%
#322945000000
1!
1%
#322950000000
0!
0%
#322955000000
1!
1%
#322960000000
0!
0%
#322965000000
1!
1%
#322970000000
0!
0%
#322975000000
1!
1%
#322980000000
0!
0%
#322985000000
1!
1%
#322990000000
0!
0%
#322995000000
1!
1%
#323000000000
0!
0%
#323005000000
1!
1%
#323010000000
0!
0%
#323015000000
1!
1%
#323020000000
0!
0%
#323025000000
1!
1%
#323030000000
0!
0%
#323035000000
1!
1%
#323040000000
0!
0%
#323045000000
1!
1%
#323050000000
0!
0%
#323055000000
1!
1%
#323060000000
0!
0%
#323065000000
1!
1%
#323070000000
0!
0%
#323075000000
1!
1%
#323080000000
0!
0%
#323085000000
1!
1%
#323090000000
0!
0%
#323095000000
1!
1%
#323100000000
0!
0%
#323105000000
1!
1%
#323110000000
0!
0%
#323115000000
1!
1%
#323120000000
0!
0%
#323125000000
1!
1%
#323130000000
0!
0%
#323135000000
1!
1%
#323140000000
0!
0%
#323145000000
1!
1%
#323150000000
0!
0%
#323155000000
1!
1%
#323160000000
0!
0%
#323165000000
1!
1%
#323170000000
0!
0%
#323175000000
1!
1%
#323180000000
0!
0%
#323185000000
1!
1%
#323190000000
0!
0%
#323195000000
1!
1%
#323200000000
0!
0%
#323205000000
1!
1%
#323210000000
0!
0%
#323215000000
1!
1%
#323220000000
0!
0%
#323225000000
1!
1%
#323230000000
0!
0%
#323235000000
1!
1%
#323240000000
0!
0%
#323245000000
1!
1%
#323250000000
0!
0%
#323255000000
1!
1%
#323260000000
0!
0%
#323265000000
1!
1%
#323270000000
0!
0%
#323275000000
1!
1%
#323280000000
0!
0%
#323285000000
1!
1%
#323290000000
0!
0%
#323295000000
1!
1%
#323300000000
0!
0%
#323305000000
1!
1%
#323310000000
0!
0%
#323315000000
1!
1%
#323320000000
0!
0%
#323325000000
1!
1%
#323330000000
0!
0%
#323335000000
1!
1%
#323340000000
0!
0%
#323345000000
1!
1%
#323350000000
0!
0%
#323355000000
1!
1%
#323360000000
0!
0%
#323365000000
1!
1%
#323370000000
0!
0%
#323375000000
1!
1%
#323380000000
0!
0%
#323385000000
1!
1%
#323390000000
0!
0%
#323395000000
1!
1%
#323400000000
0!
0%
#323405000000
1!
1%
#323410000000
0!
0%
#323415000000
1!
1%
#323420000000
0!
0%
#323425000000
1!
1%
#323430000000
0!
0%
#323435000000
1!
1%
#323440000000
0!
0%
#323445000000
1!
1%
#323450000000
0!
0%
#323455000000
1!
1%
#323460000000
0!
0%
#323465000000
1!
1%
#323470000000
0!
0%
#323475000000
1!
1%
#323480000000
0!
0%
#323485000000
1!
1%
#323490000000
0!
0%
#323495000000
1!
1%
#323500000000
0!
0%
#323505000000
1!
1%
#323510000000
0!
0%
#323515000000
1!
1%
#323520000000
0!
0%
#323525000000
1!
1%
#323530000000
0!
0%
#323535000000
1!
1%
#323540000000
0!
0%
#323545000000
1!
1%
#323550000000
0!
0%
#323555000000
1!
1%
#323560000000
0!
0%
#323565000000
1!
1%
#323570000000
0!
0%
#323575000000
1!
1%
#323580000000
0!
0%
#323585000000
1!
1%
#323590000000
0!
0%
#323595000000
1!
1%
#323600000000
0!
0%
#323605000000
1!
1%
#323610000000
0!
0%
#323615000000
1!
1%
#323620000000
0!
0%
#323625000000
1!
1%
#323630000000
0!
0%
#323635000000
1!
1%
#323640000000
0!
0%
#323645000000
1!
1%
#323650000000
0!
0%
#323655000000
1!
1%
#323660000000
0!
0%
#323665000000
1!
1%
#323670000000
0!
0%
#323675000000
1!
1%
#323680000000
0!
0%
#323685000000
1!
1%
#323690000000
0!
0%
#323695000000
1!
1%
#323700000000
0!
0%
#323705000000
1!
1%
#323710000000
0!
0%
#323715000000
1!
1%
#323720000000
0!
0%
#323725000000
1!
1%
#323730000000
0!
0%
#323735000000
1!
1%
#323740000000
0!
0%
#323745000000
1!
1%
#323750000000
0!
0%
#323755000000
1!
1%
#323760000000
0!
0%
#323765000000
1!
1%
#323770000000
0!
0%
#323775000000
1!
1%
#323780000000
0!
0%
#323785000000
1!
1%
#323790000000
0!
0%
#323795000000
1!
1%
#323800000000
0!
0%
#323805000000
1!
1%
#323810000000
0!
0%
#323815000000
1!
1%
#323820000000
0!
0%
#323825000000
1!
1%
#323830000000
0!
0%
#323835000000
1!
1%
#323840000000
0!
0%
#323845000000
1!
1%
#323850000000
0!
0%
#323855000000
1!
1%
#323860000000
0!
0%
#323865000000
1!
1%
#323870000000
0!
0%
#323875000000
1!
1%
#323880000000
0!
0%
#323885000000
1!
1%
#323890000000
0!
0%
#323895000000
1!
1%
#323900000000
0!
0%
#323905000000
1!
1%
#323910000000
0!
0%
#323915000000
1!
1%
#323920000000
0!
0%
#323925000000
1!
1%
#323930000000
0!
0%
#323935000000
1!
1%
#323940000000
0!
0%
#323945000000
1!
1%
#323950000000
0!
0%
#323955000000
1!
1%
#323960000000
0!
0%
#323965000000
1!
1%
#323970000000
0!
0%
#323975000000
1!
1%
#323980000000
0!
0%
#323985000000
1!
1%
#323990000000
0!
0%
#323995000000
1!
1%
#324000000000
0!
0%
#324005000000
1!
1%
#324010000000
0!
0%
#324015000000
1!
1%
#324020000000
0!
0%
#324025000000
1!
1%
#324030000000
0!
0%
#324035000000
1!
1%
#324040000000
0!
0%
#324045000000
1!
1%
#324050000000
0!
0%
#324055000000
1!
1%
#324060000000
0!
0%
#324065000000
1!
1%
#324070000000
0!
0%
#324075000000
1!
1%
#324080000000
0!
0%
#324085000000
1!
1%
#324090000000
0!
0%
#324095000000
1!
1%
#324100000000
0!
0%
#324105000000
1!
1%
#324110000000
0!
0%
#324115000000
1!
1%
#324120000000
0!
0%
#324125000000
1!
1%
#324130000000
0!
0%
#324135000000
1!
1%
#324140000000
0!
0%
#324145000000
1!
1%
#324150000000
0!
0%
#324155000000
1!
1%
#324160000000
0!
0%
#324165000000
1!
1%
#324170000000
0!
0%
#324175000000
1!
1%
#324180000000
0!
0%
#324185000000
1!
1%
#324190000000
0!
0%
#324195000000
1!
1%
#324200000000
0!
0%
#324205000000
1!
1%
#324210000000
0!
0%
#324215000000
1!
1%
#324220000000
0!
0%
#324225000000
1!
1%
#324230000000
0!
0%
#324235000000
1!
1%
#324240000000
0!
0%
#324245000000
1!
1%
#324250000000
0!
0%
#324255000000
1!
1%
#324260000000
0!
0%
#324265000000
1!
1%
#324270000000
0!
0%
#324275000000
1!
1%
#324280000000
0!
0%
#324285000000
1!
1%
#324290000000
0!
0%
#324295000000
1!
1%
#324300000000
0!
0%
#324305000000
1!
1%
#324310000000
0!
0%
#324315000000
1!
1%
#324320000000
0!
0%
#324325000000
1!
1%
#324330000000
0!
0%
#324335000000
1!
1%
#324340000000
0!
0%
#324345000000
1!
1%
#324350000000
0!
0%
#324355000000
1!
1%
#324360000000
0!
0%
#324365000000
1!
1%
#324370000000
0!
0%
#324375000000
1!
1%
#324380000000
0!
0%
#324385000000
1!
1%
#324390000000
0!
0%
#324395000000
1!
1%
#324400000000
0!
0%
#324405000000
1!
1%
#324410000000
0!
0%
#324415000000
1!
1%
#324420000000
0!
0%
#324425000000
1!
1%
#324430000000
0!
0%
#324435000000
1!
1%
#324440000000
0!
0%
#324445000000
1!
1%
#324450000000
0!
0%
#324455000000
1!
1%
#324460000000
0!
0%
#324465000000
1!
1%
#324470000000
0!
0%
#324475000000
1!
1%
#324480000000
0!
0%
#324485000000
1!
1%
#324490000000
0!
0%
#324495000000
1!
1%
#324500000000
0!
0%
#324505000000
1!
1%
#324510000000
0!
0%
#324515000000
1!
1%
#324520000000
0!
0%
#324525000000
1!
1%
#324530000000
0!
0%
#324535000000
1!
1%
#324540000000
0!
0%
#324545000000
1!
1%
#324550000000
0!
0%
#324555000000
1!
1%
#324560000000
0!
0%
#324565000000
1!
1%
#324570000000
0!
0%
#324575000000
1!
1%
#324580000000
0!
0%
#324585000000
1!
1%
#324590000000
0!
0%
#324595000000
1!
1%
#324600000000
0!
0%
#324605000000
1!
1%
#324610000000
0!
0%
#324615000000
1!
1%
#324620000000
0!
0%
#324625000000
1!
1%
#324630000000
0!
0%
#324635000000
1!
1%
#324640000000
0!
0%
#324645000000
1!
1%
#324650000000
0!
0%
#324655000000
1!
1%
#324660000000
0!
0%
#324665000000
1!
1%
#324670000000
0!
0%
#324675000000
1!
1%
#324680000000
0!
0%
#324685000000
1!
1%
#324690000000
0!
0%
#324695000000
1!
1%
#324700000000
0!
0%
#324705000000
1!
1%
#324710000000
0!
0%
#324715000000
1!
1%
#324720000000
0!
0%
#324725000000
1!
1%
#324730000000
0!
0%
#324735000000
1!
1%
#324740000000
0!
0%
#324745000000
1!
1%
#324750000000
0!
0%
#324755000000
1!
1%
#324760000000
0!
0%
#324765000000
1!
1%
#324770000000
0!
0%
#324775000000
1!
1%
#324780000000
0!
0%
#324785000000
1!
1%
#324790000000
0!
0%
#324795000000
1!
1%
#324800000000
0!
0%
#324805000000
1!
1%
#324810000000
0!
0%
#324815000000
1!
1%
#324820000000
0!
0%
#324825000000
1!
1%
#324830000000
0!
0%
#324835000000
1!
1%
#324840000000
0!
0%
#324845000000
1!
1%
#324850000000
0!
0%
#324855000000
1!
1%
#324860000000
0!
0%
#324865000000
1!
1%
#324870000000
0!
0%
#324875000000
1!
1%
#324880000000
0!
0%
#324885000000
1!
1%
#324890000000
0!
0%
#324895000000
1!
1%
#324900000000
0!
0%
#324905000000
1!
1%
#324910000000
0!
0%
#324915000000
1!
1%
#324920000000
0!
0%
#324925000000
1!
1%
#324930000000
0!
0%
#324935000000
1!
1%
#324940000000
0!
0%
#324945000000
1!
1%
#324950000000
0!
0%
#324955000000
1!
1%
#324960000000
0!
0%
#324965000000
1!
1%
#324970000000
0!
0%
#324975000000
1!
1%
#324980000000
0!
0%
#324985000000
1!
1%
#324990000000
0!
0%
#324995000000
1!
1%
#325000000000
0!
0%
#325005000000
1!
1%
#325010000000
0!
0%
#325015000000
1!
1%
#325020000000
0!
0%
#325025000000
1!
1%
#325030000000
0!
0%
#325035000000
1!
1%
#325040000000
0!
0%
#325045000000
1!
1%
#325050000000
0!
0%
#325055000000
1!
1%
#325060000000
0!
0%
#325065000000
1!
1%
#325070000000
0!
0%
#325075000000
1!
1%
#325080000000
0!
0%
#325085000000
1!
1%
#325090000000
0!
0%
#325095000000
1!
1%
#325100000000
0!
0%
#325105000000
1!
1%
#325110000000
0!
0%
#325115000000
1!
1%
#325120000000
0!
0%
#325125000000
1!
1%
#325130000000
0!
0%
#325135000000
1!
1%
#325140000000
0!
0%
#325145000000
1!
1%
#325150000000
0!
0%
#325155000000
1!
1%
#325160000000
0!
0%
#325165000000
1!
1%
#325170000000
0!
0%
#325175000000
1!
1%
#325180000000
0!
0%
#325185000000
1!
1%
#325190000000
0!
0%
#325195000000
1!
1%
#325200000000
0!
0%
#325205000000
1!
1%
#325210000000
0!
0%
#325215000000
1!
1%
#325220000000
0!
0%
#325225000000
1!
1%
#325230000000
0!
0%
#325235000000
1!
1%
#325240000000
0!
0%
#325245000000
1!
1%
#325250000000
0!
0%
#325255000000
1!
1%
#325260000000
0!
0%
#325265000000
1!
1%
#325270000000
0!
0%
#325275000000
1!
1%
#325280000000
0!
0%
#325285000000
1!
1%
#325290000000
0!
0%
#325295000000
1!
1%
#325300000000
0!
0%
#325305000000
1!
1%
#325310000000
0!
0%
#325315000000
1!
1%
#325320000000
0!
0%
#325325000000
1!
1%
#325330000000
0!
0%
#325335000000
1!
1%
#325340000000
0!
0%
#325345000000
1!
1%
#325350000000
0!
0%
#325355000000
1!
1%
#325360000000
0!
0%
#325365000000
1!
1%
#325370000000
0!
0%
#325375000000
1!
1%
#325380000000
0!
0%
#325385000000
1!
1%
#325390000000
0!
0%
#325395000000
1!
1%
#325400000000
0!
0%
#325405000000
1!
1%
#325410000000
0!
0%
#325415000000
1!
1%
#325420000000
0!
0%
#325425000000
1!
1%
#325430000000
0!
0%
#325435000000
1!
1%
#325440000000
0!
0%
#325445000000
1!
1%
#325450000000
0!
0%
#325455000000
1!
1%
#325460000000
0!
0%
#325465000000
1!
1%
#325470000000
0!
0%
#325475000000
1!
1%
#325480000000
0!
0%
#325485000000
1!
1%
#325490000000
0!
0%
#325495000000
1!
1%
#325500000000
0!
0%
#325505000000
1!
1%
#325510000000
0!
0%
#325515000000
1!
1%
#325520000000
0!
0%
#325525000000
1!
1%
#325530000000
0!
0%
#325535000000
1!
1%
#325540000000
0!
0%
#325545000000
1!
1%
#325550000000
0!
0%
#325555000000
1!
1%
#325560000000
0!
0%
#325565000000
1!
1%
#325570000000
0!
0%
#325575000000
1!
1%
#325580000000
0!
0%
#325585000000
1!
1%
#325590000000
0!
0%
#325595000000
1!
1%
#325600000000
0!
0%
#325605000000
1!
1%
#325610000000
0!
0%
#325615000000
1!
1%
#325620000000
0!
0%
#325625000000
1!
1%
#325630000000
0!
0%
#325635000000
1!
1%
#325640000000
0!
0%
#325645000000
1!
1%
#325650000000
0!
0%
#325655000000
1!
1%
#325660000000
0!
0%
#325665000000
1!
1%
#325670000000
0!
0%
#325675000000
1!
1%
#325680000000
0!
0%
#325685000000
1!
1%
#325690000000
0!
0%
#325695000000
1!
1%
#325700000000
0!
0%
#325705000000
1!
1%
#325710000000
0!
0%
#325715000000
1!
1%
#325720000000
0!
0%
#325725000000
1!
1%
#325730000000
0!
0%
#325735000000
1!
1%
#325740000000
0!
0%
#325745000000
1!
1%
#325750000000
0!
0%
#325755000000
1!
1%
#325760000000
0!
0%
#325765000000
1!
1%
#325770000000
0!
0%
#325775000000
1!
1%
#325780000000
0!
0%
#325785000000
1!
1%
#325790000000
0!
0%
#325795000000
1!
1%
#325800000000
0!
0%
#325805000000
1!
1%
#325810000000
0!
0%
#325815000000
1!
1%
#325820000000
0!
0%
#325825000000
1!
1%
#325830000000
0!
0%
#325835000000
1!
1%
#325840000000
0!
0%
#325845000000
1!
1%
#325850000000
0!
0%
#325855000000
1!
1%
#325860000000
0!
0%
#325865000000
1!
1%
#325870000000
0!
0%
#325875000000
1!
1%
#325880000000
0!
0%
#325885000000
1!
1%
#325890000000
0!
0%
#325895000000
1!
1%
#325900000000
0!
0%
#325905000000
1!
1%
#325910000000
0!
0%
#325915000000
1!
1%
#325920000000
0!
0%
#325925000000
1!
1%
#325930000000
0!
0%
#325935000000
1!
1%
#325940000000
0!
0%
#325945000000
1!
1%
#325950000000
0!
0%
#325955000000
1!
1%
#325960000000
0!
0%
#325965000000
1!
1%
#325970000000
0!
0%
#325975000000
1!
1%
#325980000000
0!
0%
#325985000000
1!
1%
#325990000000
0!
0%
#325995000000
1!
1%
#326000000000
0!
0%
#326005000000
1!
1%
#326010000000
0!
0%
#326015000000
1!
1%
#326020000000
0!
0%
#326025000000
1!
1%
#326030000000
0!
0%
#326035000000
1!
1%
#326040000000
0!
0%
#326045000000
1!
1%
#326050000000
0!
0%
#326055000000
1!
1%
#326060000000
0!
0%
#326065000000
1!
1%
#326070000000
0!
0%
#326075000000
1!
1%
#326080000000
0!
0%
#326085000000
1!
1%
#326090000000
0!
0%
#326095000000
1!
1%
#326100000000
0!
0%
#326105000000
1!
1%
#326110000000
0!
0%
#326115000000
1!
1%
#326120000000
0!
0%
#326125000000
1!
1%
#326130000000
0!
0%
#326135000000
1!
1%
#326140000000
0!
0%
#326145000000
1!
1%
#326150000000
0!
0%
#326155000000
1!
1%
#326160000000
0!
0%
#326165000000
1!
1%
#326170000000
0!
0%
#326175000000
1!
1%
#326180000000
0!
0%
#326185000000
1!
1%
#326190000000
0!
0%
#326195000000
1!
1%
#326200000000
0!
0%
#326205000000
1!
1%
#326210000000
0!
0%
#326215000000
1!
1%
#326220000000
0!
0%
#326225000000
1!
1%
#326230000000
0!
0%
#326235000000
1!
1%
#326240000000
0!
0%
#326245000000
1!
1%
#326250000000
0!
0%
#326255000000
1!
1%
#326260000000
0!
0%
#326265000000
1!
1%
#326270000000
0!
0%
#326275000000
1!
1%
#326280000000
0!
0%
#326285000000
1!
1%
#326290000000
0!
0%
#326295000000
1!
1%
#326300000000
0!
0%
#326305000000
1!
1%
#326310000000
0!
0%
#326315000000
1!
1%
#326320000000
0!
0%
#326325000000
1!
1%
#326330000000
0!
0%
#326335000000
1!
1%
#326340000000
0!
0%
#326345000000
1!
1%
#326350000000
0!
0%
#326355000000
1!
1%
#326360000000
0!
0%
#326365000000
1!
1%
#326370000000
0!
0%
#326375000000
1!
1%
#326380000000
0!
0%
#326385000000
1!
1%
#326390000000
0!
0%
#326395000000
1!
1%
#326400000000
0!
0%
#326405000000
1!
1%
#326410000000
0!
0%
#326415000000
1!
1%
#326420000000
0!
0%
#326425000000
1!
1%
#326430000000
0!
0%
#326435000000
1!
1%
#326440000000
0!
0%
#326445000000
1!
1%
#326450000000
0!
0%
#326455000000
1!
1%
#326460000000
0!
0%
#326465000000
1!
1%
#326470000000
0!
0%
#326475000000
1!
1%
#326480000000
0!
0%
#326485000000
1!
1%
#326490000000
0!
0%
#326495000000
1!
1%
#326500000000
0!
0%
#326505000000
1!
1%
#326510000000
0!
0%
#326515000000
1!
1%
#326520000000
0!
0%
#326525000000
1!
1%
#326530000000
0!
0%
#326535000000
1!
1%
#326540000000
0!
0%
#326545000000
1!
1%
#326550000000
0!
0%
#326555000000
1!
1%
#326560000000
0!
0%
#326565000000
1!
1%
#326570000000
0!
0%
#326575000000
1!
1%
#326580000000
0!
0%
#326585000000
1!
1%
#326590000000
0!
0%
#326595000000
1!
1%
#326600000000
0!
0%
#326605000000
1!
1%
#326610000000
0!
0%
#326615000000
1!
1%
#326620000000
0!
0%
#326625000000
1!
1%
#326630000000
0!
0%
#326635000000
1!
1%
#326640000000
0!
0%
#326645000000
1!
1%
#326650000000
0!
0%
#326655000000
1!
1%
#326660000000
0!
0%
#326665000000
1!
1%
#326670000000
0!
0%
#326675000000
1!
1%
#326680000000
0!
0%
#326685000000
1!
1%
#326690000000
0!
0%
#326695000000
1!
1%
#326700000000
0!
0%
#326705000000
1!
1%
#326710000000
0!
0%
#326715000000
1!
1%
#326720000000
0!
0%
#326725000000
1!
1%
#326730000000
0!
0%
#326735000000
1!
1%
#326740000000
0!
0%
#326745000000
1!
1%
#326750000000
0!
0%
#326755000000
1!
1%
#326760000000
0!
0%
#326765000000
1!
1%
#326770000000
0!
0%
#326775000000
1!
1%
#326780000000
0!
0%
#326785000000
1!
1%
#326790000000
0!
0%
#326795000000
1!
1%
#326800000000
0!
0%
#326805000000
1!
1%
#326810000000
0!
0%
#326815000000
1!
1%
#326820000000
0!
0%
#326825000000
1!
1%
#326830000000
0!
0%
#326835000000
1!
1%
#326840000000
0!
0%
#326845000000
1!
1%
#326850000000
0!
0%
#326855000000
1!
1%
#326860000000
0!
0%
#326865000000
1!
1%
#326870000000
0!
0%
#326875000000
1!
1%
#326880000000
0!
0%
#326885000000
1!
1%
#326890000000
0!
0%
#326895000000
1!
1%
#326900000000
0!
0%
#326905000000
1!
1%
#326910000000
0!
0%
#326915000000
1!
1%
#326920000000
0!
0%
#326925000000
1!
1%
#326930000000
0!
0%
#326935000000
1!
1%
#326940000000
0!
0%
#326945000000
1!
1%
#326950000000
0!
0%
#326955000000
1!
1%
#326960000000
0!
0%
#326965000000
1!
1%
#326970000000
0!
0%
#326975000000
1!
1%
#326980000000
0!
0%
#326985000000
1!
1%
#326990000000
0!
0%
#326995000000
1!
1%
#327000000000
0!
0%
#327005000000
1!
1%
#327010000000
0!
0%
#327015000000
1!
1%
#327020000000
0!
0%
#327025000000
1!
1%
#327030000000
0!
0%
#327035000000
1!
1%
#327040000000
0!
0%
#327045000000
1!
1%
#327050000000
0!
0%
#327055000000
1!
1%
#327060000000
0!
0%
#327065000000
1!
1%
#327070000000
0!
0%
#327075000000
1!
1%
#327080000000
0!
0%
#327085000000
1!
1%
#327090000000
0!
0%
#327095000000
1!
1%
#327100000000
0!
0%
#327105000000
1!
1%
#327110000000
0!
0%
#327115000000
1!
1%
#327120000000
0!
0%
#327125000000
1!
1%
#327130000000
0!
0%
#327135000000
1!
1%
#327140000000
0!
0%
#327145000000
1!
1%
#327150000000
0!
0%
#327155000000
1!
1%
#327160000000
0!
0%
#327165000000
1!
1%
#327170000000
0!
0%
#327175000000
1!
1%
#327180000000
0!
0%
#327185000000
1!
1%
#327190000000
0!
0%
#327195000000
1!
1%
#327200000000
0!
0%
#327205000000
1!
1%
#327210000000
0!
0%
#327215000000
1!
1%
#327220000000
0!
0%
#327225000000
1!
1%
#327230000000
0!
0%
#327235000000
1!
1%
#327240000000
0!
0%
#327245000000
1!
1%
#327250000000
0!
0%
#327255000000
1!
1%
#327260000000
0!
0%
#327265000000
1!
1%
#327270000000
0!
0%
#327275000000
1!
1%
#327280000000
0!
0%
#327285000000
1!
1%
#327290000000
0!
0%
#327295000000
1!
1%
#327300000000
0!
0%
#327305000000
1!
1%
#327310000000
0!
0%
#327315000000
1!
1%
#327320000000
0!
0%
#327325000000
1!
1%
#327330000000
0!
0%
#327335000000
1!
1%
#327340000000
0!
0%
#327345000000
1!
1%
#327350000000
0!
0%
#327355000000
1!
1%
#327360000000
0!
0%
#327365000000
1!
1%
#327370000000
0!
0%
#327375000000
1!
1%
#327380000000
0!
0%
#327385000000
1!
1%
#327390000000
0!
0%
#327395000000
1!
1%
#327400000000
0!
0%
#327405000000
1!
1%
#327410000000
0!
0%
#327415000000
1!
1%
#327420000000
0!
0%
#327425000000
1!
1%
#327430000000
0!
0%
#327435000000
1!
1%
#327440000000
0!
0%
#327445000000
1!
1%
#327450000000
0!
0%
#327455000000
1!
1%
#327460000000
0!
0%
#327465000000
1!
1%
#327470000000
0!
0%
#327475000000
1!
1%
#327480000000
0!
0%
#327485000000
1!
1%
#327490000000
0!
0%
#327495000000
1!
1%
#327500000000
0!
0%
#327505000000
1!
1%
#327510000000
0!
0%
#327515000000
1!
1%
#327520000000
0!
0%
#327525000000
1!
1%
#327530000000
0!
0%
#327535000000
1!
1%
#327540000000
0!
0%
#327545000000
1!
1%
#327550000000
0!
0%
#327555000000
1!
1%
#327560000000
0!
0%
#327565000000
1!
1%
#327570000000
0!
0%
#327575000000
1!
1%
#327580000000
0!
0%
#327585000000
1!
1%
#327590000000
0!
0%
#327595000000
1!
1%
#327600000000
0!
0%
#327605000000
1!
1%
#327610000000
0!
0%
#327615000000
1!
1%
#327620000000
0!
0%
#327625000000
1!
1%
#327630000000
0!
0%
#327635000000
1!
1%
#327640000000
0!
0%
#327645000000
1!
1%
#327650000000
0!
0%
#327655000000
1!
1%
#327660000000
0!
0%
#327665000000
1!
1%
#327670000000
0!
0%
#327675000000
1!
1%
#327680000000
0!
0%
#327685000000
1!
1%
#327690000000
0!
0%
#327695000000
1!
1%
#327700000000
0!
0%
#327705000000
1!
1%
#327710000000
0!
0%
#327715000000
1!
1%
#327720000000
0!
0%
#327725000000
1!
1%
#327730000000
0!
0%
#327735000000
1!
1%
#327740000000
0!
0%
#327745000000
1!
1%
#327750000000
0!
0%
#327755000000
1!
1%
#327760000000
0!
0%
#327765000000
1!
1%
#327770000000
0!
0%
#327775000000
1!
1%
#327780000000
0!
0%
#327785000000
1!
1%
#327790000000
0!
0%
#327795000000
1!
1%
#327800000000
0!
0%
#327805000000
1!
1%
#327810000000
0!
0%
#327815000000
1!
1%
#327820000000
0!
0%
#327825000000
1!
1%
#327830000000
0!
0%
#327835000000
1!
1%
#327840000000
0!
0%
#327845000000
1!
1%
#327850000000
0!
0%
#327855000000
1!
1%
#327860000000
0!
0%
#327865000000
1!
1%
#327870000000
0!
0%
#327875000000
1!
1%
#327880000000
0!
0%
#327885000000
1!
1%
#327890000000
0!
0%
#327895000000
1!
1%
#327900000000
0!
0%
#327905000000
1!
1%
#327910000000
0!
0%
#327915000000
1!
1%
#327920000000
0!
0%
#327925000000
1!
1%
#327930000000
0!
0%
#327935000000
1!
1%
#327940000000
0!
0%
#327945000000
1!
1%
#327950000000
0!
0%
#327955000000
1!
1%
#327960000000
0!
0%
#327965000000
1!
1%
#327970000000
0!
0%
#327975000000
1!
1%
#327980000000
0!
0%
#327985000000
1!
1%
#327990000000
0!
0%
#327995000000
1!
1%
#328000000000
0!
0%
#328005000000
1!
1%
#328010000000
0!
0%
#328015000000
1!
1%
#328020000000
0!
0%
#328025000000
1!
1%
#328030000000
0!
0%
#328035000000
1!
1%
#328040000000
0!
0%
#328045000000
1!
1%
#328050000000
0!
0%
#328055000000
1!
1%
#328060000000
0!
0%
#328065000000
1!
1%
#328070000000
0!
0%
#328075000000
1!
1%
#328080000000
0!
0%
#328085000000
1!
1%
#328090000000
0!
0%
#328095000000
1!
1%
#328100000000
0!
0%
#328105000000
1!
1%
#328110000000
0!
0%
#328115000000
1!
1%
#328120000000
0!
0%
#328125000000
1!
1%
#328130000000
0!
0%
#328135000000
1!
1%
#328140000000
0!
0%
#328145000000
1!
1%
#328150000000
0!
0%
#328155000000
1!
1%
#328160000000
0!
0%
#328165000000
1!
1%
#328170000000
0!
0%
#328175000000
1!
1%
#328180000000
0!
0%
#328185000000
1!
1%
#328190000000
0!
0%
#328195000000
1!
1%
#328200000000
0!
0%
#328205000000
1!
1%
#328210000000
0!
0%
#328215000000
1!
1%
#328220000000
0!
0%
#328225000000
1!
1%
#328230000000
0!
0%
#328235000000
1!
1%
#328240000000
0!
0%
#328245000000
1!
1%
#328250000000
0!
0%
#328255000000
1!
1%
#328260000000
0!
0%
#328265000000
1!
1%
#328270000000
0!
0%
#328275000000
1!
1%
#328280000000
0!
0%
#328285000000
1!
1%
#328290000000
0!
0%
#328295000000
1!
1%
#328300000000
0!
0%
#328305000000
1!
1%
#328310000000
0!
0%
#328315000000
1!
1%
#328320000000
0!
0%
#328325000000
1!
1%
#328330000000
0!
0%
#328335000000
1!
1%
#328340000000
0!
0%
#328345000000
1!
1%
#328350000000
0!
0%
#328355000000
1!
1%
#328360000000
0!
0%
#328365000000
1!
1%
#328370000000
0!
0%
#328375000000
1!
1%
#328380000000
0!
0%
#328385000000
1!
1%
#328390000000
0!
0%
#328395000000
1!
1%
#328400000000
0!
0%
#328405000000
1!
1%
#328410000000
0!
0%
#328415000000
1!
1%
#328420000000
0!
0%
#328425000000
1!
1%
#328430000000
0!
0%
#328435000000
1!
1%
#328440000000
0!
0%
#328445000000
1!
1%
#328450000000
0!
0%
#328455000000
1!
1%
#328460000000
0!
0%
#328465000000
1!
1%
#328470000000
0!
0%
#328475000000
1!
1%
#328480000000
0!
0%
#328485000000
1!
1%
#328490000000
0!
0%
#328495000000
1!
1%
#328500000000
0!
0%
#328505000000
1!
1%
#328510000000
0!
0%
#328515000000
1!
1%
#328520000000
0!
0%
#328525000000
1!
1%
#328530000000
0!
0%
#328535000000
1!
1%
#328540000000
0!
0%
#328545000000
1!
1%
#328550000000
0!
0%
#328555000000
1!
1%
#328560000000
0!
0%
#328565000000
1!
1%
#328570000000
0!
0%
#328575000000
1!
1%
#328580000000
0!
0%
#328585000000
1!
1%
#328590000000
0!
0%
#328595000000
1!
1%
#328600000000
0!
0%
#328605000000
1!
1%
#328610000000
0!
0%
#328615000000
1!
1%
#328620000000
0!
0%
#328625000000
1!
1%
#328630000000
0!
0%
#328635000000
1!
1%
#328640000000
0!
0%
#328645000000
1!
1%
#328650000000
0!
0%
#328655000000
1!
1%
#328660000000
0!
0%
#328665000000
1!
1%
#328670000000
0!
0%
#328675000000
1!
1%
#328680000000
0!
0%
#328685000000
1!
1%
#328690000000
0!
0%
#328695000000
1!
1%
#328700000000
0!
0%
#328705000000
1!
1%
#328710000000
0!
0%
#328715000000
1!
1%
#328720000000
0!
0%
#328725000000
1!
1%
#328730000000
0!
0%
#328735000000
1!
1%
#328740000000
0!
0%
#328745000000
1!
1%
#328750000000
0!
0%
#328755000000
1!
1%
#328760000000
0!
0%
#328765000000
1!
1%
#328770000000
0!
0%
#328775000000
1!
1%
#328780000000
0!
0%
#328785000000
1!
1%
#328790000000
0!
0%
#328795000000
1!
1%
#328800000000
0!
0%
#328805000000
1!
1%
#328810000000
0!
0%
#328815000000
1!
1%
#328820000000
0!
0%
#328825000000
1!
1%
#328830000000
0!
0%
#328835000000
1!
1%
#328840000000
0!
0%
#328845000000
1!
1%
#328850000000
0!
0%
#328855000000
1!
1%
#328860000000
0!
0%
#328865000000
1!
1%
#328870000000
0!
0%
#328875000000
1!
1%
#328880000000
0!
0%
#328885000000
1!
1%
#328890000000
0!
0%
#328895000000
1!
1%
#328900000000
0!
0%
#328905000000
1!
1%
#328910000000
0!
0%
#328915000000
1!
1%
#328920000000
0!
0%
#328925000000
1!
1%
#328930000000
0!
0%
#328935000000
1!
1%
#328940000000
0!
0%
#328945000000
1!
1%
#328950000000
0!
0%
#328955000000
1!
1%
#328960000000
0!
0%
#328965000000
1!
1%
#328970000000
0!
0%
#328975000000
1!
1%
#328980000000
0!
0%
#328985000000
1!
1%
#328990000000
0!
0%
#328995000000
1!
1%
#329000000000
0!
0%
#329005000000
1!
1%
#329010000000
0!
0%
#329015000000
1!
1%
#329020000000
0!
0%
#329025000000
1!
1%
#329030000000
0!
0%
#329035000000
1!
1%
#329040000000
0!
0%
#329045000000
1!
1%
#329050000000
0!
0%
#329055000000
1!
1%
#329060000000
0!
0%
#329065000000
1!
1%
#329070000000
0!
0%
#329075000000
1!
1%
#329080000000
0!
0%
#329085000000
1!
1%
#329090000000
0!
0%
#329095000000
1!
1%
#329100000000
0!
0%
#329105000000
1!
1%
#329110000000
0!
0%
#329115000000
1!
1%
#329120000000
0!
0%
#329125000000
1!
1%
#329130000000
0!
0%
#329135000000
1!
1%
#329140000000
0!
0%
#329145000000
1!
1%
#329150000000
0!
0%
#329155000000
1!
1%
#329160000000
0!
0%
#329165000000
1!
1%
#329170000000
0!
0%
#329175000000
1!
1%
#329180000000
0!
0%
#329185000000
1!
1%
#329190000000
0!
0%
#329195000000
1!
1%
#329200000000
0!
0%
#329205000000
1!
1%
#329210000000
0!
0%
#329215000000
1!
1%
#329220000000
0!
0%
#329225000000
1!
1%
#329230000000
0!
0%
#329235000000
1!
1%
#329240000000
0!
0%
#329245000000
1!
1%
#329250000000
0!
0%
#329255000000
1!
1%
#329260000000
0!
0%
#329265000000
1!
1%
#329270000000
0!
0%
#329275000000
1!
1%
#329280000000
0!
0%
#329285000000
1!
1%
#329290000000
0!
0%
#329295000000
1!
1%
#329300000000
0!
0%
#329305000000
1!
1%
#329310000000
0!
0%
#329315000000
1!
1%
#329320000000
0!
0%
#329325000000
1!
1%
#329330000000
0!
0%
#329335000000
1!
1%
#329340000000
0!
0%
#329345000000
1!
1%
#329350000000
0!
0%
#329355000000
1!
1%
#329360000000
0!
0%
#329365000000
1!
1%
#329370000000
0!
0%
#329375000000
1!
1%
#329380000000
0!
0%
#329385000000
1!
1%
#329390000000
0!
0%
#329395000000
1!
1%
#329400000000
0!
0%
#329405000000
1!
1%
#329410000000
0!
0%
#329415000000
1!
1%
#329420000000
0!
0%
#329425000000
1!
1%
#329430000000
0!
0%
#329435000000
1!
1%
#329440000000
0!
0%
#329445000000
1!
1%
#329450000000
0!
0%
#329455000000
1!
1%
#329460000000
0!
0%
#329465000000
1!
1%
#329470000000
0!
0%
#329475000000
1!
1%
#329480000000
0!
0%
#329485000000
1!
1%
#329490000000
0!
0%
#329495000000
1!
1%
#329500000000
0!
0%
#329505000000
1!
1%
#329510000000
0!
0%
#329515000000
1!
1%
#329520000000
0!
0%
#329525000000
1!
1%
#329530000000
0!
0%
#329535000000
1!
1%
#329540000000
0!
0%
#329545000000
1!
1%
#329550000000
0!
0%
#329555000000
1!
1%
#329560000000
0!
0%
#329565000000
1!
1%
#329570000000
0!
0%
#329575000000
1!
1%
#329580000000
0!
0%
#329585000000
1!
1%
#329590000000
0!
0%
#329595000000
1!
1%
#329600000000
0!
0%
#329605000000
1!
1%
#329610000000
0!
0%
#329615000000
1!
1%
#329620000000
0!
0%
#329625000000
1!
1%
#329630000000
0!
0%
#329635000000
1!
1%
#329640000000
0!
0%
#329645000000
1!
1%
#329650000000
0!
0%
#329655000000
1!
1%
#329660000000
0!
0%
#329665000000
1!
1%
#329670000000
0!
0%
#329675000000
1!
1%
#329680000000
0!
0%
#329685000000
1!
1%
#329690000000
0!
0%
#329695000000
1!
1%
#329700000000
0!
0%
#329705000000
1!
1%
#329710000000
0!
0%
#329715000000
1!
1%
#329720000000
0!
0%
#329725000000
1!
1%
#329730000000
0!
0%
#329735000000
1!
1%
#329740000000
0!
0%
#329745000000
1!
1%
#329750000000
0!
0%
#329755000000
1!
1%
#329760000000
0!
0%
#329765000000
1!
1%
#329770000000
0!
0%
#329775000000
1!
1%
#329780000000
0!
0%
#329785000000
1!
1%
#329790000000
0!
0%
#329795000000
1!
1%
#329800000000
0!
0%
#329805000000
1!
1%
#329810000000
0!
0%
#329815000000
1!
1%
#329820000000
0!
0%
#329825000000
1!
1%
#329830000000
0!
0%
#329835000000
1!
1%
#329840000000
0!
0%
#329845000000
1!
1%
#329850000000
0!
0%
#329855000000
1!
1%
#329860000000
0!
0%
#329865000000
1!
1%
#329870000000
0!
0%
#329875000000
1!
1%
#329880000000
0!
0%
#329885000000
1!
1%
#329890000000
0!
0%
#329895000000
1!
1%
#329900000000
0!
0%
#329905000000
1!
1%
#329910000000
0!
0%
#329915000000
1!
1%
#329920000000
0!
0%
#329925000000
1!
1%
#329930000000
0!
0%
#329935000000
1!
1%
#329940000000
0!
0%
#329945000000
1!
1%
#329950000000
0!
0%
#329955000000
1!
1%
#329960000000
0!
0%
#329965000000
1!
1%
#329970000000
0!
0%
#329975000000
1!
1%
#329980000000
0!
0%
#329985000000
1!
1%
#329990000000
0!
0%
#329995000000
1!
1%
#330000000000
0!
0%
#330005000000
1!
1%
#330010000000
0!
0%
#330015000000
1!
1%
#330020000000
0!
0%
#330025000000
1!
1%
#330030000000
0!
0%
#330035000000
1!
1%
#330040000000
0!
0%
#330045000000
1!
1%
#330050000000
0!
0%
#330055000000
1!
1%
#330060000000
0!
0%
#330065000000
1!
1%
#330070000000
0!
0%
#330075000000
1!
1%
#330080000000
0!
0%
#330085000000
1!
1%
#330090000000
0!
0%
#330095000000
1!
1%
#330100000000
0!
0%
#330105000000
1!
1%
#330110000000
0!
0%
#330115000000
1!
1%
#330120000000
0!
0%
#330125000000
1!
1%
#330130000000
0!
0%
#330135000000
1!
1%
#330140000000
0!
0%
#330145000000
1!
1%
#330150000000
0!
0%
#330155000000
1!
1%
#330160000000
0!
0%
#330165000000
1!
1%
#330170000000
0!
0%
#330175000000
1!
1%
#330180000000
0!
0%
#330185000000
1!
1%
#330190000000
0!
0%
#330195000000
1!
1%
#330200000000
0!
0%
#330205000000
1!
1%
#330210000000
0!
0%
#330215000000
1!
1%
#330220000000
0!
0%
#330225000000
1!
1%
#330230000000
0!
0%
#330235000000
1!
1%
#330240000000
0!
0%
#330245000000
1!
1%
#330250000000
0!
0%
#330255000000
1!
1%
#330260000000
0!
0%
#330265000000
1!
1%
#330270000000
0!
0%
#330275000000
1!
1%
#330280000000
0!
0%
#330285000000
1!
1%
#330290000000
0!
0%
#330295000000
1!
1%
#330300000000
0!
0%
#330305000000
1!
1%
#330310000000
0!
0%
#330315000000
1!
1%
#330320000000
0!
0%
#330325000000
1!
1%
#330330000000
0!
0%
#330335000000
1!
1%
#330340000000
0!
0%
#330345000000
1!
1%
#330350000000
0!
0%
#330355000000
1!
1%
#330360000000
0!
0%
#330365000000
1!
1%
#330370000000
0!
0%
#330375000000
1!
1%
#330380000000
0!
0%
#330385000000
1!
1%
#330390000000
0!
0%
#330395000000
1!
1%
#330400000000
0!
0%
#330405000000
1!
1%
#330410000000
0!
0%
#330415000000
1!
1%
#330420000000
0!
0%
#330425000000
1!
1%
#330430000000
0!
0%
#330435000000
1!
1%
#330440000000
0!
0%
#330445000000
1!
1%
#330450000000
0!
0%
#330455000000
1!
1%
#330460000000
0!
0%
#330465000000
1!
1%
#330470000000
0!
0%
#330475000000
1!
1%
#330480000000
0!
0%
#330485000000
1!
1%
#330490000000
0!
0%
#330495000000
1!
1%
#330500000000
0!
0%
#330505000000
1!
1%
#330510000000
0!
0%
#330515000000
1!
1%
#330520000000
0!
0%
#330525000000
1!
1%
#330530000000
0!
0%
#330535000000
1!
1%
#330540000000
0!
0%
#330545000000
1!
1%
#330550000000
0!
0%
#330555000000
1!
1%
#330560000000
0!
0%
#330565000000
1!
1%
#330570000000
0!
0%
#330575000000
1!
1%
#330580000000
0!
0%
#330585000000
1!
1%
#330590000000
0!
0%
#330595000000
1!
1%
#330600000000
0!
0%
#330605000000
1!
1%
#330610000000
0!
0%
#330615000000
1!
1%
#330620000000
0!
0%
#330625000000
1!
1%
#330630000000
0!
0%
#330635000000
1!
1%
#330640000000
0!
0%
#330645000000
1!
1%
#330650000000
0!
0%
#330655000000
1!
1%
#330660000000
0!
0%
#330665000000
1!
1%
#330670000000
0!
0%
#330675000000
1!
1%
#330680000000
0!
0%
#330685000000
1!
1%
#330690000000
0!
0%
#330695000000
1!
1%
#330700000000
0!
0%
#330705000000
1!
1%
#330710000000
0!
0%
#330715000000
1!
1%
#330720000000
0!
0%
#330725000000
1!
1%
#330730000000
0!
0%
#330735000000
1!
1%
#330740000000
0!
0%
#330745000000
1!
1%
#330750000000
0!
0%
#330755000000
1!
1%
#330760000000
0!
0%
#330765000000
1!
1%
#330770000000
0!
0%
#330775000000
1!
1%
#330780000000
0!
0%
#330785000000
1!
1%
#330790000000
0!
0%
#330795000000
1!
1%
#330800000000
0!
0%
#330805000000
1!
1%
#330810000000
0!
0%
#330815000000
1!
1%
#330820000000
0!
0%
#330825000000
1!
1%
#330830000000
0!
0%
#330835000000
1!
1%
#330840000000
0!
0%
#330845000000
1!
1%
#330850000000
0!
0%
#330855000000
1!
1%
#330860000000
0!
0%
#330865000000
1!
1%
#330870000000
0!
0%
#330875000000
1!
1%
#330880000000
0!
0%
#330885000000
1!
1%
#330890000000
0!
0%
#330895000000
1!
1%
#330900000000
0!
0%
#330905000000
1!
1%
#330910000000
0!
0%
#330915000000
1!
1%
#330920000000
0!
0%
#330925000000
1!
1%
#330930000000
0!
0%
#330935000000
1!
1%
#330940000000
0!
0%
#330945000000
1!
1%
#330950000000
0!
0%
#330955000000
1!
1%
#330960000000
0!
0%
#330965000000
1!
1%
#330970000000
0!
0%
#330975000000
1!
1%
#330980000000
0!
0%
#330985000000
1!
1%
#330990000000
0!
0%
#330995000000
1!
1%
#331000000000
0!
0%
#331005000000
1!
1%
#331010000000
0!
0%
#331015000000
1!
1%
#331020000000
0!
0%
#331025000000
1!
1%
#331030000000
0!
0%
#331035000000
1!
1%
#331040000000
0!
0%
#331045000000
1!
1%
#331050000000
0!
0%
#331055000000
1!
1%
#331060000000
0!
0%
#331065000000
1!
1%
#331070000000
0!
0%
#331075000000
1!
1%
#331080000000
0!
0%
#331085000000
1!
1%
#331090000000
0!
0%
#331095000000
1!
1%
#331100000000
0!
0%
#331105000000
1!
1%
#331110000000
0!
0%
#331115000000
1!
1%
#331120000000
0!
0%
#331125000000
1!
1%
#331130000000
0!
0%
#331135000000
1!
1%
#331140000000
0!
0%
#331145000000
1!
1%
#331150000000
0!
0%
#331155000000
1!
1%
#331160000000
0!
0%
#331165000000
1!
1%
#331170000000
0!
0%
#331175000000
1!
1%
#331180000000
0!
0%
#331185000000
1!
1%
#331190000000
0!
0%
#331195000000
1!
1%
#331200000000
0!
0%
#331205000000
1!
1%
#331210000000
0!
0%
#331215000000
1!
1%
#331220000000
0!
0%
#331225000000
1!
1%
#331230000000
0!
0%
#331235000000
1!
1%
#331240000000
0!
0%
#331245000000
1!
1%
#331250000000
0!
0%
#331255000000
1!
1%
#331260000000
0!
0%
#331265000000
1!
1%
#331270000000
0!
0%
#331275000000
1!
1%
#331280000000
0!
0%
#331285000000
1!
1%
#331290000000
0!
0%
#331295000000
1!
1%
#331300000000
0!
0%
#331305000000
1!
1%
#331310000000
0!
0%
#331315000000
1!
1%
#331320000000
0!
0%
#331325000000
1!
1%
#331330000000
0!
0%
#331335000000
1!
1%
#331340000000
0!
0%
#331345000000
1!
1%
#331350000000
0!
0%
#331355000000
1!
1%
#331360000000
0!
0%
#331365000000
1!
1%
#331370000000
0!
0%
#331375000000
1!
1%
#331380000000
0!
0%
#331385000000
1!
1%
#331390000000
0!
0%
#331395000000
1!
1%
#331400000000
0!
0%
#331405000000
1!
1%
#331410000000
0!
0%
#331415000000
1!
1%
#331420000000
0!
0%
#331425000000
1!
1%
#331430000000
0!
0%
#331435000000
1!
1%
#331440000000
0!
0%
#331445000000
1!
1%
#331450000000
0!
0%
#331455000000
1!
1%
#331460000000
0!
0%
#331465000000
1!
1%
#331470000000
0!
0%
#331475000000
1!
1%
#331480000000
0!
0%
#331485000000
1!
1%
#331490000000
0!
0%
#331495000000
1!
1%
#331500000000
0!
0%
#331505000000
1!
1%
#331510000000
0!
0%
#331515000000
1!
1%
#331520000000
0!
0%
#331525000000
1!
1%
#331530000000
0!
0%
#331535000000
1!
1%
#331540000000
0!
0%
#331545000000
1!
1%
#331550000000
0!
0%
#331555000000
1!
1%
#331560000000
0!
0%
#331565000000
1!
1%
#331570000000
0!
0%
#331575000000
1!
1%
#331580000000
0!
0%
#331585000000
1!
1%
#331590000000
0!
0%
#331595000000
1!
1%
#331600000000
0!
0%
#331605000000
1!
1%
#331610000000
0!
0%
#331615000000
1!
1%
#331620000000
0!
0%
#331625000000
1!
1%
#331630000000
0!
0%
#331635000000
1!
1%
#331640000000
0!
0%
#331645000000
1!
1%
#331650000000
0!
0%
#331655000000
1!
1%
#331660000000
0!
0%
#331665000000
1!
1%
#331670000000
0!
0%
#331675000000
1!
1%
#331680000000
0!
0%
#331685000000
1!
1%
#331690000000
0!
0%
#331695000000
1!
1%
#331700000000
0!
0%
#331705000000
1!
1%
#331710000000
0!
0%
#331715000000
1!
1%
#331720000000
0!
0%
#331725000000
1!
1%
#331730000000
0!
0%
#331735000000
1!
1%
#331740000000
0!
0%
#331745000000
1!
1%
#331750000000
0!
0%
#331755000000
1!
1%
#331760000000
0!
0%
#331765000000
1!
1%
#331770000000
0!
0%
#331775000000
1!
1%
#331780000000
0!
0%
#331785000000
1!
1%
#331790000000
0!
0%
#331795000000
1!
1%
#331800000000
0!
0%
#331805000000
1!
1%
#331810000000
0!
0%
#331815000000
1!
1%
#331820000000
0!
0%
#331825000000
1!
1%
#331830000000
0!
0%
#331835000000
1!
1%
#331840000000
0!
0%
#331845000000
1!
1%
#331850000000
0!
0%
#331855000000
1!
1%
#331860000000
0!
0%
#331865000000
1!
1%
#331870000000
0!
0%
#331875000000
1!
1%
#331880000000
0!
0%
#331885000000
1!
1%
#331890000000
0!
0%
#331895000000
1!
1%
#331900000000
0!
0%
#331905000000
1!
1%
#331910000000
0!
0%
#331915000000
1!
1%
#331920000000
0!
0%
#331925000000
1!
1%
#331930000000
0!
0%
#331935000000
1!
1%
#331940000000
0!
0%
#331945000000
1!
1%
#331950000000
0!
0%
#331955000000
1!
1%
#331960000000
0!
0%
#331965000000
1!
1%
#331970000000
0!
0%
#331975000000
1!
1%
#331980000000
0!
0%
#331985000000
1!
1%
#331990000000
0!
0%
#331995000000
1!
1%
#332000000000
0!
0%
#332005000000
1!
1%
#332010000000
0!
0%
#332015000000
1!
1%
#332020000000
0!
0%
#332025000000
1!
1%
#332030000000
0!
0%
#332035000000
1!
1%
#332040000000
0!
0%
#332045000000
1!
1%
#332050000000
0!
0%
#332055000000
1!
1%
#332060000000
0!
0%
#332065000000
1!
1%
#332070000000
0!
0%
#332075000000
1!
1%
#332080000000
0!
0%
#332085000000
1!
1%
#332090000000
0!
0%
#332095000000
1!
1%
#332100000000
0!
0%
#332105000000
1!
1%
#332110000000
0!
0%
#332115000000
1!
1%
#332120000000
0!
0%
#332125000000
1!
1%
#332130000000
0!
0%
#332135000000
1!
1%
#332140000000
0!
0%
#332145000000
1!
1%
#332150000000
0!
0%
#332155000000
1!
1%
#332160000000
0!
0%
#332165000000
1!
1%
#332170000000
0!
0%
#332175000000
1!
1%
#332180000000
0!
0%
#332185000000
1!
1%
#332190000000
0!
0%
#332195000000
1!
1%
#332200000000
0!
0%
#332205000000
1!
1%
#332210000000
0!
0%
#332215000000
1!
1%
#332220000000
0!
0%
#332225000000
1!
1%
#332230000000
0!
0%
#332235000000
1!
1%
#332240000000
0!
0%
#332245000000
1!
1%
#332250000000
0!
0%
#332255000000
1!
1%
#332260000000
0!
0%
#332265000000
1!
1%
#332270000000
0!
0%
#332275000000
1!
1%
#332280000000
0!
0%
#332285000000
1!
1%
#332290000000
0!
0%
#332295000000
1!
1%
#332300000000
0!
0%
#332305000000
1!
1%
#332310000000
0!
0%
#332315000000
1!
1%
#332320000000
0!
0%
#332325000000
1!
1%
#332330000000
0!
0%
#332335000000
1!
1%
#332340000000
0!
0%
#332345000000
1!
1%
#332350000000
0!
0%
#332355000000
1!
1%
#332360000000
0!
0%
#332365000000
1!
1%
#332370000000
0!
0%
#332375000000
1!
1%
#332380000000
0!
0%
#332385000000
1!
1%
#332390000000
0!
0%
#332395000000
1!
1%
#332400000000
0!
0%
#332405000000
1!
1%
#332410000000
0!
0%
#332415000000
1!
1%
#332420000000
0!
0%
#332425000000
1!
1%
#332430000000
0!
0%
#332435000000
1!
1%
#332440000000
0!
0%
#332445000000
1!
1%
#332450000000
0!
0%
#332455000000
1!
1%
#332460000000
0!
0%
#332465000000
1!
1%
#332470000000
0!
0%
#332475000000
1!
1%
#332480000000
0!
0%
#332485000000
1!
1%
#332490000000
0!
0%
#332495000000
1!
1%
#332500000000
0!
0%
#332505000000
1!
1%
#332510000000
0!
0%
#332515000000
1!
1%
#332520000000
0!
0%
#332525000000
1!
1%
#332530000000
0!
0%
#332535000000
1!
1%
#332540000000
0!
0%
#332545000000
1!
1%
#332550000000
0!
0%
#332555000000
1!
1%
#332560000000
0!
0%
#332565000000
1!
1%
#332570000000
0!
0%
#332575000000
1!
1%
#332580000000
0!
0%
#332585000000
1!
1%
#332590000000
0!
0%
#332595000000
1!
1%
#332600000000
0!
0%
#332605000000
1!
1%
#332610000000
0!
0%
#332615000000
1!
1%
#332620000000
0!
0%
#332625000000
1!
1%
#332630000000
0!
0%
#332635000000
1!
1%
#332640000000
0!
0%
#332645000000
1!
1%
#332650000000
0!
0%
#332655000000
1!
1%
#332660000000
0!
0%
#332665000000
1!
1%
#332670000000
0!
0%
#332675000000
1!
1%
#332680000000
0!
0%
#332685000000
1!
1%
#332690000000
0!
0%
#332695000000
1!
1%
#332700000000
0!
0%
#332705000000
1!
1%
#332710000000
0!
0%
#332715000000
1!
1%
#332720000000
0!
0%
#332725000000
1!
1%
#332730000000
0!
0%
#332735000000
1!
1%
#332740000000
0!
0%
#332745000000
1!
1%
#332750000000
0!
0%
#332755000000
1!
1%
#332760000000
0!
0%
#332765000000
1!
1%
#332770000000
0!
0%
#332775000000
1!
1%
#332780000000
0!
0%
#332785000000
1!
1%
#332790000000
0!
0%
#332795000000
1!
1%
#332800000000
0!
0%
#332805000000
1!
1%
#332810000000
0!
0%
#332815000000
1!
1%
#332820000000
0!
0%
#332825000000
1!
1%
#332830000000
0!
0%
#332835000000
1!
1%
#332840000000
0!
0%
#332845000000
1!
1%
#332850000000
0!
0%
#332855000000
1!
1%
#332860000000
0!
0%
#332865000000
1!
1%
#332870000000
0!
0%
#332875000000
1!
1%
#332880000000
0!
0%
#332885000000
1!
1%
#332890000000
0!
0%
#332895000000
1!
1%
#332900000000
0!
0%
#332905000000
1!
1%
#332910000000
0!
0%
#332915000000
1!
1%
#332920000000
0!
0%
#332925000000
1!
1%
#332930000000
0!
0%
#332935000000
1!
1%
#332940000000
0!
0%
#332945000000
1!
1%
#332950000000
0!
0%
#332955000000
1!
1%
#332960000000
0!
0%
#332965000000
1!
1%
#332970000000
0!
0%
#332975000000
1!
1%
#332980000000
0!
0%
#332985000000
1!
1%
#332990000000
0!
0%
#332995000000
1!
1%
#333000000000
0!
0%
#333005000000
1!
1%
#333010000000
0!
0%
#333015000000
1!
1%
#333020000000
0!
0%
#333025000000
1!
1%
#333030000000
0!
0%
#333035000000
1!
1%
#333040000000
0!
0%
#333045000000
1!
1%
#333050000000
0!
0%
#333055000000
1!
1%
#333060000000
0!
0%
#333065000000
1!
1%
#333070000000
0!
0%
#333075000000
1!
1%
#333080000000
0!
0%
#333085000000
1!
1%
#333090000000
0!
0%
#333095000000
1!
1%
#333100000000
0!
0%
#333105000000
1!
1%
#333110000000
0!
0%
#333115000000
1!
1%
#333120000000
0!
0%
#333125000000
1!
1%
#333130000000
0!
0%
#333135000000
1!
1%
#333140000000
0!
0%
#333145000000
1!
1%
#333150000000
0!
0%
#333155000000
1!
1%
#333160000000
0!
0%
#333165000000
1!
1%
#333170000000
0!
0%
#333175000000
1!
1%
#333180000000
0!
0%
#333185000000
1!
1%
#333190000000
0!
0%
#333195000000
1!
1%
#333200000000
0!
0%
#333205000000
1!
1%
#333210000000
0!
0%
#333215000000
1!
1%
#333220000000
0!
0%
#333225000000
1!
1%
#333230000000
0!
0%
#333235000000
1!
1%
#333240000000
0!
0%
#333245000000
1!
1%
#333250000000
0!
0%
#333255000000
1!
1%
#333260000000
0!
0%
#333265000000
1!
1%
#333270000000
0!
0%
#333275000000
1!
1%
#333280000000
0!
0%
#333285000000
1!
1%
#333290000000
0!
0%
#333295000000
1!
1%
#333300000000
0!
0%
#333305000000
1!
1%
#333310000000
0!
0%
#333315000000
1!
1%
#333320000000
0!
0%
#333325000000
1!
1%
#333330000000
0!
0%
#333335000000
1!
1%
#333340000000
0!
0%
#333345000000
1!
1%
#333350000000
0!
0%
#333355000000
1!
1%
#333360000000
0!
0%
#333365000000
1!
1%
#333370000000
0!
0%
#333375000000
1!
1%
#333380000000
0!
0%
#333385000000
1!
1%
#333390000000
0!
0%
#333395000000
1!
1%
#333400000000
0!
0%
#333405000000
1!
1%
#333410000000
0!
0%
#333415000000
1!
1%
#333420000000
0!
0%
#333425000000
1!
1%
#333430000000
0!
0%
#333435000000
1!
1%
#333440000000
0!
0%
#333445000000
1!
1%
#333450000000
0!
0%
#333455000000
1!
1%
#333460000000
0!
0%
#333465000000
1!
1%
#333470000000
0!
0%
#333475000000
1!
1%
#333480000000
0!
0%
#333485000000
1!
1%
#333490000000
0!
0%
#333495000000
1!
1%
#333500000000
0!
0%
#333505000000
1!
1%
#333510000000
0!
0%
#333515000000
1!
1%
#333520000000
0!
0%
#333525000000
1!
1%
#333530000000
0!
0%
#333535000000
1!
1%
#333540000000
0!
0%
#333545000000
1!
1%
#333550000000
0!
0%
#333555000000
1!
1%
#333560000000
0!
0%
#333565000000
1!
1%
#333570000000
0!
0%
#333575000000
1!
1%
#333580000000
0!
0%
#333585000000
1!
1%
#333590000000
0!
0%
#333595000000
1!
1%
#333600000000
0!
0%
#333605000000
1!
1%
#333610000000
0!
0%
#333615000000
1!
1%
#333620000000
0!
0%
#333625000000
1!
1%
#333630000000
0!
0%
#333635000000
1!
1%
#333640000000
0!
0%
#333645000000
1!
1%
#333650000000
0!
0%
#333655000000
1!
1%
#333660000000
0!
0%
#333665000000
1!
1%
#333670000000
0!
0%
#333675000000
1!
1%
#333680000000
0!
0%
#333685000000
1!
1%
#333690000000
0!
0%
#333695000000
1!
1%
#333700000000
0!
0%
#333705000000
1!
1%
#333710000000
0!
0%
#333715000000
1!
1%
#333720000000
0!
0%
#333725000000
1!
1%
#333730000000
0!
0%
#333735000000
1!
1%
#333740000000
0!
0%
#333745000000
1!
1%
#333750000000
0!
0%
#333755000000
1!
1%
#333760000000
0!
0%
#333765000000
1!
1%
#333770000000
0!
0%
#333775000000
1!
1%
#333780000000
0!
0%
#333785000000
1!
1%
#333790000000
0!
0%
#333795000000
1!
1%
#333800000000
0!
0%
#333805000000
1!
1%
#333810000000
0!
0%
#333815000000
1!
1%
#333820000000
0!
0%
#333825000000
1!
1%
#333830000000
0!
0%
#333835000000
1!
1%
#333840000000
0!
0%
#333845000000
1!
1%
#333850000000
0!
0%
#333855000000
1!
1%
#333860000000
0!
0%
#333865000000
1!
1%
#333870000000
0!
0%
#333875000000
1!
1%
#333880000000
0!
0%
#333885000000
1!
1%
#333890000000
0!
0%
#333895000000
1!
1%
#333900000000
0!
0%
#333905000000
1!
1%
#333910000000
0!
0%
#333915000000
1!
1%
#333920000000
0!
0%
#333925000000
1!
1%
#333930000000
0!
0%
#333935000000
1!
1%
#333940000000
0!
0%
#333945000000
1!
1%
#333950000000
0!
0%
#333955000000
1!
1%
#333960000000
0!
0%
#333965000000
1!
1%
#333970000000
0!
0%
#333975000000
1!
1%
#333980000000
0!
0%
#333985000000
1!
1%
#333990000000
0!
0%
#333995000000
1!
1%
#334000000000
0!
0%
#334005000000
1!
1%
#334010000000
0!
0%
#334015000000
1!
1%
#334020000000
0!
0%
#334025000000
1!
1%
#334030000000
0!
0%
#334035000000
1!
1%
#334040000000
0!
0%
#334045000000
1!
1%
#334050000000
0!
0%
#334055000000
1!
1%
#334060000000
0!
0%
#334065000000
1!
1%
#334070000000
0!
0%
#334075000000
1!
1%
#334080000000
0!
0%
#334085000000
1!
1%
#334090000000
0!
0%
#334095000000
1!
1%
#334100000000
0!
0%
#334105000000
1!
1%
#334110000000
0!
0%
#334115000000
1!
1%
#334120000000
0!
0%
#334125000000
1!
1%
#334130000000
0!
0%
#334135000000
1!
1%
#334140000000
0!
0%
#334145000000
1!
1%
#334150000000
0!
0%
#334155000000
1!
1%
#334160000000
0!
0%
#334165000000
1!
1%
#334170000000
0!
0%
#334175000000
1!
1%
#334180000000
0!
0%
#334185000000
1!
1%
#334190000000
0!
0%
#334195000000
1!
1%
#334200000000
0!
0%
#334205000000
1!
1%
#334210000000
0!
0%
#334215000000
1!
1%
#334220000000
0!
0%
#334225000000
1!
1%
#334230000000
0!
0%
#334235000000
1!
1%
#334240000000
0!
0%
#334245000000
1!
1%
#334250000000
0!
0%
#334255000000
1!
1%
#334260000000
0!
0%
#334265000000
1!
1%
#334270000000
0!
0%
#334275000000
1!
1%
#334280000000
0!
0%
#334285000000
1!
1%
#334290000000
0!
0%
#334295000000
1!
1%
#334300000000
0!
0%
#334305000000
1!
1%
#334310000000
0!
0%
#334315000000
1!
1%
#334320000000
0!
0%
#334325000000
1!
1%
#334330000000
0!
0%
#334335000000
1!
1%
#334340000000
0!
0%
#334345000000
1!
1%
#334350000000
0!
0%
#334355000000
1!
1%
#334360000000
0!
0%
#334365000000
1!
1%
#334370000000
0!
0%
#334375000000
1!
1%
#334380000000
0!
0%
#334385000000
1!
1%
#334390000000
0!
0%
#334395000000
1!
1%
#334400000000
0!
0%
#334405000000
1!
1%
#334410000000
0!
0%
#334415000000
1!
1%
#334420000000
0!
0%
#334425000000
1!
1%
#334430000000
0!
0%
#334435000000
1!
1%
#334440000000
0!
0%
#334445000000
1!
1%
#334450000000
0!
0%
#334455000000
1!
1%
#334460000000
0!
0%
#334465000000
1!
1%
#334470000000
0!
0%
#334475000000
1!
1%
#334480000000
0!
0%
#334485000000
1!
1%
#334490000000
0!
0%
#334495000000
1!
1%
#334500000000
0!
0%
#334505000000
1!
1%
#334510000000
0!
0%
#334515000000
1!
1%
#334520000000
0!
0%
#334525000000
1!
1%
#334530000000
0!
0%
#334535000000
1!
1%
#334540000000
0!
0%
#334545000000
1!
1%
#334550000000
0!
0%
#334555000000
1!
1%
#334560000000
0!
0%
#334565000000
1!
1%
#334570000000
0!
0%
#334575000000
1!
1%
#334580000000
0!
0%
#334585000000
1!
1%
#334590000000
0!
0%
#334595000000
1!
1%
#334600000000
0!
0%
#334605000000
1!
1%
#334610000000
0!
0%
#334615000000
1!
1%
#334620000000
0!
0%
#334625000000
1!
1%
#334630000000
0!
0%
#334635000000
1!
1%
#334640000000
0!
0%
#334645000000
1!
1%
#334650000000
0!
0%
#334655000000
1!
1%
#334660000000
0!
0%
#334665000000
1!
1%
#334670000000
0!
0%
#334675000000
1!
1%
#334680000000
0!
0%
#334685000000
1!
1%
#334690000000
0!
0%
#334695000000
1!
1%
#334700000000
0!
0%
#334705000000
1!
1%
#334710000000
0!
0%
#334715000000
1!
1%
#334720000000
0!
0%
#334725000000
1!
1%
#334730000000
0!
0%
#334735000000
1!
1%
#334740000000
0!
0%
#334745000000
1!
1%
#334750000000
0!
0%
#334755000000
1!
1%
#334760000000
0!
0%
#334765000000
1!
1%
#334770000000
0!
0%
#334775000000
1!
1%
#334780000000
0!
0%
#334785000000
1!
1%
#334790000000
0!
0%
#334795000000
1!
1%
#334800000000
0!
0%
#334805000000
1!
1%
#334810000000
0!
0%
#334815000000
1!
1%
#334820000000
0!
0%
#334825000000
1!
1%
#334830000000
0!
0%
#334835000000
1!
1%
#334840000000
0!
0%
#334845000000
1!
1%
#334850000000
0!
0%
#334855000000
1!
1%
#334860000000
0!
0%
#334865000000
1!
1%
#334870000000
0!
0%
#334875000000
1!
1%
#334880000000
0!
0%
#334885000000
1!
1%
#334890000000
0!
0%
#334895000000
1!
1%
#334900000000
0!
0%
#334905000000
1!
1%
#334910000000
0!
0%
#334915000000
1!
1%
#334920000000
0!
0%
#334925000000
1!
1%
#334930000000
0!
0%
#334935000000
1!
1%
#334940000000
0!
0%
#334945000000
1!
1%
#334950000000
0!
0%
#334955000000
1!
1%
#334960000000
0!
0%
#334965000000
1!
1%
#334970000000
0!
0%
#334975000000
1!
1%
#334980000000
0!
0%
#334985000000
1!
1%
#334990000000
0!
0%
#334995000000
1!
1%
#335000000000
0!
0%
#335005000000
1!
1%
#335010000000
0!
0%
#335015000000
1!
1%
#335020000000
0!
0%
#335025000000
1!
1%
#335030000000
0!
0%
#335035000000
1!
1%
#335040000000
0!
0%
#335045000000
1!
1%
#335050000000
0!
0%
#335055000000
1!
1%
#335060000000
0!
0%
#335065000000
1!
1%
#335070000000
0!
0%
#335075000000
1!
1%
#335080000000
0!
0%
#335085000000
1!
1%
#335090000000
0!
0%
#335095000000
1!
1%
#335100000000
0!
0%
#335105000000
1!
1%
#335110000000
0!
0%
#335115000000
1!
1%
#335120000000
0!
0%
#335125000000
1!
1%
#335130000000
0!
0%
#335135000000
1!
1%
#335140000000
0!
0%
#335145000000
1!
1%
#335150000000
0!
0%
#335155000000
1!
1%
#335160000000
0!
0%
#335165000000
1!
1%
#335170000000
0!
0%
#335175000000
1!
1%
#335180000000
0!
0%
#335185000000
1!
1%
#335190000000
0!
0%
#335195000000
1!
1%
#335200000000
0!
0%
#335205000000
1!
1%
#335210000000
0!
0%
#335215000000
1!
1%
#335220000000
0!
0%
#335225000000
1!
1%
#335230000000
0!
0%
#335235000000
1!
1%
#335240000000
0!
0%
#335245000000
1!
1%
#335250000000
0!
0%
#335255000000
1!
1%
#335260000000
0!
0%
#335265000000
1!
1%
#335270000000
0!
0%
#335275000000
1!
1%
#335280000000
0!
0%
#335285000000
1!
1%
#335290000000
0!
0%
#335295000000
1!
1%
#335300000000
0!
0%
#335305000000
1!
1%
#335310000000
0!
0%
#335315000000
1!
1%
#335320000000
0!
0%
#335325000000
1!
1%
#335330000000
0!
0%
#335335000000
1!
1%
#335340000000
0!
0%
#335345000000
1!
1%
#335350000000
0!
0%
#335355000000
1!
1%
#335360000000
0!
0%
#335365000000
1!
1%
#335370000000
0!
0%
#335375000000
1!
1%
#335380000000
0!
0%
#335385000000
1!
1%
#335390000000
0!
0%
#335395000000
1!
1%
#335400000000
0!
0%
#335405000000
1!
1%
#335410000000
0!
0%
#335415000000
1!
1%
#335420000000
0!
0%
#335425000000
1!
1%
#335430000000
0!
0%
#335435000000
1!
1%
#335440000000
0!
0%
#335445000000
1!
1%
#335450000000
0!
0%
#335455000000
1!
1%
#335460000000
0!
0%
#335465000000
1!
1%
#335470000000
0!
0%
#335475000000
1!
1%
#335480000000
0!
0%
#335485000000
1!
1%
#335490000000
0!
0%
#335495000000
1!
1%
#335500000000
0!
0%
#335505000000
1!
1%
#335510000000
0!
0%
#335515000000
1!
1%
#335520000000
0!
0%
#335525000000
1!
1%
#335530000000
0!
0%
#335535000000
1!
1%
#335540000000
0!
0%
#335545000000
1!
1%
#335550000000
0!
0%
#335555000000
1!
1%
#335560000000
0!
0%
#335565000000
1!
1%
#335570000000
0!
0%
#335575000000
1!
1%
#335580000000
0!
0%
#335585000000
1!
1%
#335590000000
0!
0%
#335595000000
1!
1%
#335600000000
0!
0%
#335605000000
1!
1%
#335610000000
0!
0%
#335615000000
1!
1%
#335620000000
0!
0%
#335625000000
1!
1%
#335630000000
0!
0%
#335635000000
1!
1%
#335640000000
0!
0%
#335645000000
1!
1%
#335650000000
0!
0%
#335655000000
1!
1%
#335660000000
0!
0%
#335665000000
1!
1%
#335670000000
0!
0%
#335675000000
1!
1%
#335680000000
0!
0%
#335685000000
1!
1%
#335690000000
0!
0%
#335695000000
1!
1%
#335700000000
0!
0%
#335705000000
1!
1%
#335710000000
0!
0%
#335715000000
1!
1%
#335720000000
0!
0%
#335725000000
1!
1%
#335730000000
0!
0%
#335735000000
1!
1%
#335740000000
0!
0%
#335745000000
1!
1%
#335750000000
0!
0%
#335755000000
1!
1%
#335760000000
0!
0%
#335765000000
1!
1%
#335770000000
0!
0%
#335775000000
1!
1%
#335780000000
0!
0%
#335785000000
1!
1%
#335790000000
0!
0%
#335795000000
1!
1%
#335800000000
0!
0%
#335805000000
1!
1%
#335810000000
0!
0%
#335815000000
1!
1%
#335820000000
0!
0%
#335825000000
1!
1%
#335830000000
0!
0%
#335835000000
1!
1%
#335840000000
0!
0%
#335845000000
1!
1%
#335850000000
0!
0%
#335855000000
1!
1%
#335860000000
0!
0%
#335865000000
1!
1%
#335870000000
0!
0%
#335875000000
1!
1%
#335880000000
0!
0%
#335885000000
1!
1%
#335890000000
0!
0%
#335895000000
1!
1%
#335900000000
0!
0%
#335905000000
1!
1%
#335910000000
0!
0%
#335915000000
1!
1%
#335920000000
0!
0%
#335925000000
1!
1%
#335930000000
0!
0%
#335935000000
1!
1%
#335940000000
0!
0%
#335945000000
1!
1%
#335950000000
0!
0%
#335955000000
1!
1%
#335960000000
0!
0%
#335965000000
1!
1%
#335970000000
0!
0%
#335975000000
1!
1%
#335980000000
0!
0%
#335985000000
1!
1%
#335990000000
0!
0%
#335995000000
1!
1%
#336000000000
0!
0%
#336005000000
1!
1%
#336010000000
0!
0%
#336015000000
1!
1%
#336020000000
0!
0%
#336025000000
1!
1%
#336030000000
0!
0%
#336035000000
1!
1%
#336040000000
0!
0%
#336045000000
1!
1%
#336050000000
0!
0%
#336055000000
1!
1%
#336060000000
0!
0%
#336065000000
1!
1%
#336070000000
0!
0%
#336075000000
1!
1%
#336080000000
0!
0%
#336085000000
1!
1%
#336090000000
0!
0%
#336095000000
1!
1%
#336100000000
0!
0%
#336105000000
1!
1%
#336110000000
0!
0%
#336115000000
1!
1%
#336120000000
0!
0%
#336125000000
1!
1%
#336130000000
0!
0%
#336135000000
1!
1%
#336140000000
0!
0%
#336145000000
1!
1%
#336150000000
0!
0%
#336155000000
1!
1%
#336160000000
0!
0%
#336165000000
1!
1%
#336170000000
0!
0%
#336175000000
1!
1%
#336180000000
0!
0%
#336185000000
1!
1%
#336190000000
0!
0%
#336195000000
1!
1%
#336200000000
0!
0%
#336205000000
1!
1%
#336210000000
0!
0%
#336215000000
1!
1%
#336220000000
0!
0%
#336225000000
1!
1%
#336230000000
0!
0%
#336235000000
1!
1%
#336240000000
0!
0%
#336245000000
1!
1%
#336250000000
0!
0%
#336255000000
1!
1%
#336260000000
0!
0%
#336265000000
1!
1%
#336270000000
0!
0%
#336275000000
1!
1%
#336280000000
0!
0%
#336285000000
1!
1%
#336290000000
0!
0%
#336295000000
1!
1%
#336300000000
0!
0%
#336305000000
1!
1%
#336310000000
0!
0%
#336315000000
1!
1%
#336320000000
0!
0%
#336325000000
1!
1%
#336330000000
0!
0%
#336335000000
1!
1%
#336340000000
0!
0%
#336345000000
1!
1%
#336350000000
0!
0%
#336355000000
1!
1%
#336360000000
0!
0%
#336365000000
1!
1%
#336370000000
0!
0%
#336375000000
1!
1%
#336380000000
0!
0%
#336385000000
1!
1%
#336390000000
0!
0%
#336395000000
1!
1%
#336400000000
0!
0%
#336405000000
1!
1%
#336410000000
0!
0%
#336415000000
1!
1%
#336420000000
0!
0%
#336425000000
1!
1%
#336430000000
0!
0%
#336435000000
1!
1%
#336440000000
0!
0%
#336445000000
1!
1%
#336450000000
0!
0%
#336455000000
1!
1%
#336460000000
0!
0%
#336465000000
1!
1%
#336470000000
0!
0%
#336475000000
1!
1%
#336480000000
0!
0%
#336485000000
1!
1%
#336490000000
0!
0%
#336495000000
1!
1%
#336500000000
0!
0%
#336505000000
1!
1%
#336510000000
0!
0%
#336515000000
1!
1%
#336520000000
0!
0%
#336525000000
1!
1%
#336530000000
0!
0%
#336535000000
1!
1%
#336540000000
0!
0%
#336545000000
1!
1%
#336550000000
0!
0%
#336555000000
1!
1%
#336560000000
0!
0%
#336565000000
1!
1%
#336570000000
0!
0%
#336575000000
1!
1%
#336580000000
0!
0%
#336585000000
1!
1%
#336590000000
0!
0%
#336595000000
1!
1%
#336600000000
0!
0%
#336605000000
1!
1%
#336610000000
0!
0%
#336615000000
1!
1%
#336620000000
0!
0%
#336625000000
1!
1%
#336630000000
0!
0%
#336635000000
1!
1%
#336640000000
0!
0%
#336645000000
1!
1%
#336650000000
0!
0%
#336655000000
1!
1%
#336660000000
0!
0%
#336665000000
1!
1%
#336670000000
0!
0%
#336675000000
1!
1%
#336680000000
0!
0%
#336685000000
1!
1%
#336690000000
0!
0%
#336695000000
1!
1%
#336700000000
0!
0%
#336705000000
1!
1%
#336710000000
0!
0%
#336715000000
1!
1%
#336720000000
0!
0%
#336725000000
1!
1%
#336730000000
0!
0%
#336735000000
1!
1%
#336740000000
0!
0%
#336745000000
1!
1%
#336750000000
0!
0%
#336755000000
1!
1%
#336760000000
0!
0%
#336765000000
1!
1%
#336770000000
0!
0%
#336775000000
1!
1%
#336780000000
0!
0%
#336785000000
1!
1%
#336790000000
0!
0%
#336795000000
1!
1%
#336800000000
0!
0%
#336805000000
1!
1%
#336810000000
0!
0%
#336815000000
1!
1%
#336820000000
0!
0%
#336825000000
1!
1%
#336830000000
0!
0%
#336835000000
1!
1%
#336840000000
0!
0%
#336845000000
1!
1%
#336850000000
0!
0%
#336855000000
1!
1%
#336860000000
0!
0%
#336865000000
1!
1%
#336870000000
0!
0%
#336875000000
1!
1%
#336880000000
0!
0%
#336885000000
1!
1%
#336890000000
0!
0%
#336895000000
1!
1%
#336900000000
0!
0%
#336905000000
1!
1%
#336910000000
0!
0%
#336915000000
1!
1%
#336920000000
0!
0%
#336925000000
1!
1%
#336930000000
0!
0%
#336935000000
1!
1%
#336940000000
0!
0%
#336945000000
1!
1%
#336950000000
0!
0%
#336955000000
1!
1%
#336960000000
0!
0%
#336965000000
1!
1%
#336970000000
0!
0%
#336975000000
1!
1%
#336980000000
0!
0%
#336985000000
1!
1%
#336990000000
0!
0%
#336995000000
1!
1%
#337000000000
0!
0%
#337005000000
1!
1%
#337010000000
0!
0%
#337015000000
1!
1%
#337020000000
0!
0%
#337025000000
1!
1%
#337030000000
0!
0%
#337035000000
1!
1%
#337040000000
0!
0%
#337045000000
1!
1%
#337050000000
0!
0%
#337055000000
1!
1%
#337060000000
0!
0%
#337065000000
1!
1%
#337070000000
0!
0%
#337075000000
1!
1%
#337080000000
0!
0%
#337085000000
1!
1%
#337090000000
0!
0%
#337095000000
1!
1%
#337100000000
0!
0%
#337105000000
1!
1%
#337110000000
0!
0%
#337115000000
1!
1%
#337120000000
0!
0%
#337125000000
1!
1%
#337130000000
0!
0%
#337135000000
1!
1%
#337140000000
0!
0%
#337145000000
1!
1%
#337150000000
0!
0%
#337155000000
1!
1%
#337160000000
0!
0%
#337165000000
1!
1%
#337170000000
0!
0%
#337175000000
1!
1%
#337180000000
0!
0%
#337185000000
1!
1%
#337190000000
0!
0%
#337195000000
1!
1%
#337200000000
0!
0%
#337205000000
1!
1%
#337210000000
0!
0%
#337215000000
1!
1%
#337220000000
0!
0%
#337225000000
1!
1%
#337230000000
0!
0%
#337235000000
1!
1%
#337240000000
0!
0%
#337245000000
1!
1%
#337250000000
0!
0%
#337255000000
1!
1%
#337260000000
0!
0%
#337265000000
1!
1%
#337270000000
0!
0%
#337275000000
1!
1%
#337280000000
0!
0%
#337285000000
1!
1%
#337290000000
0!
0%
#337295000000
1!
1%
#337300000000
0!
0%
#337305000000
1!
1%
#337310000000
0!
0%
#337315000000
1!
1%
#337320000000
0!
0%
#337325000000
1!
1%
#337330000000
0!
0%
#337335000000
1!
1%
#337340000000
0!
0%
#337345000000
1!
1%
#337350000000
0!
0%
#337355000000
1!
1%
#337360000000
0!
0%
#337365000000
1!
1%
#337370000000
0!
0%
#337375000000
1!
1%
#337380000000
0!
0%
#337385000000
1!
1%
#337390000000
0!
0%
#337395000000
1!
1%
#337400000000
0!
0%
#337405000000
1!
1%
#337410000000
0!
0%
#337415000000
1!
1%
#337420000000
0!
0%
#337425000000
1!
1%
#337430000000
0!
0%
#337435000000
1!
1%
#337440000000
0!
0%
#337445000000
1!
1%
#337450000000
0!
0%
#337455000000
1!
1%
#337460000000
0!
0%
#337465000000
1!
1%
#337470000000
0!
0%
#337475000000
1!
1%
#337480000000
0!
0%
#337485000000
1!
1%
#337490000000
0!
0%
#337495000000
1!
1%
#337500000000
0!
0%
#337505000000
1!
1%
#337510000000
0!
0%
#337515000000
1!
1%
#337520000000
0!
0%
#337525000000
1!
1%
#337530000000
0!
0%
#337535000000
1!
1%
#337540000000
0!
0%
#337545000000
1!
1%
#337550000000
0!
0%
#337555000000
1!
1%
#337560000000
0!
0%
#337565000000
1!
1%
#337570000000
0!
0%
#337575000000
1!
1%
#337580000000
0!
0%
#337585000000
1!
1%
#337590000000
0!
0%
#337595000000
1!
1%
#337600000000
0!
0%
#337605000000
1!
1%
#337610000000
0!
0%
#337615000000
1!
1%
#337620000000
0!
0%
#337625000000
1!
1%
#337630000000
0!
0%
#337635000000
1!
1%
#337640000000
0!
0%
#337645000000
1!
1%
#337650000000
0!
0%
#337655000000
1!
1%
#337660000000
0!
0%
#337665000000
1!
1%
#337670000000
0!
0%
#337675000000
1!
1%
#337680000000
0!
0%
#337685000000
1!
1%
#337690000000
0!
0%
#337695000000
1!
1%
#337700000000
0!
0%
#337705000000
1!
1%
#337710000000
0!
0%
#337715000000
1!
1%
#337720000000
0!
0%
#337725000000
1!
1%
#337730000000
0!
0%
#337735000000
1!
1%
#337740000000
0!
0%
#337745000000
1!
1%
#337750000000
0!
0%
#337755000000
1!
1%
#337760000000
0!
0%
#337765000000
1!
1%
#337770000000
0!
0%
#337775000000
1!
1%
#337780000000
0!
0%
#337785000000
1!
1%
#337790000000
0!
0%
#337795000000
1!
1%
#337800000000
0!
0%
#337805000000
1!
1%
#337810000000
0!
0%
#337815000000
1!
1%
#337820000000
0!
0%
#337825000000
1!
1%
#337830000000
0!
0%
#337835000000
1!
1%
#337840000000
0!
0%
#337845000000
1!
1%
#337850000000
0!
0%
#337855000000
1!
1%
#337860000000
0!
0%
#337865000000
1!
1%
#337870000000
0!
0%
#337875000000
1!
1%
#337880000000
0!
0%
#337885000000
1!
1%
#337890000000
0!
0%
#337895000000
1!
1%
#337900000000
0!
0%
#337905000000
1!
1%
#337910000000
0!
0%
#337915000000
1!
1%
#337920000000
0!
0%
#337925000000
1!
1%
#337930000000
0!
0%
#337935000000
1!
1%
#337940000000
0!
0%
#337945000000
1!
1%
#337950000000
0!
0%
#337955000000
1!
1%
#337960000000
0!
0%
#337965000000
1!
1%
#337970000000
0!
0%
#337975000000
1!
1%
#337980000000
0!
0%
#337985000000
1!
1%
#337990000000
0!
0%
#337995000000
1!
1%
#338000000000
0!
0%
#338005000000
1!
1%
#338010000000
0!
0%
#338015000000
1!
1%
#338020000000
0!
0%
#338025000000
1!
1%
#338030000000
0!
0%
#338035000000
1!
1%
#338040000000
0!
0%
#338045000000
1!
1%
#338050000000
0!
0%
#338055000000
1!
1%
#338060000000
0!
0%
#338065000000
1!
1%
#338070000000
0!
0%
#338075000000
1!
1%
#338080000000
0!
0%
#338085000000
1!
1%
#338090000000
0!
0%
#338095000000
1!
1%
#338100000000
0!
0%
#338105000000
1!
1%
#338110000000
0!
0%
#338115000000
1!
1%
#338120000000
0!
0%
#338125000000
1!
1%
#338130000000
0!
0%
#338135000000
1!
1%
#338140000000
0!
0%
#338145000000
1!
1%
#338150000000
0!
0%
#338155000000
1!
1%
#338160000000
0!
0%
#338165000000
1!
1%
#338170000000
0!
0%
#338175000000
1!
1%
#338180000000
0!
0%
#338185000000
1!
1%
#338190000000
0!
0%
#338195000000
1!
1%
#338200000000
0!
0%
#338205000000
1!
1%
#338210000000
0!
0%
#338215000000
1!
1%
#338220000000
0!
0%
#338225000000
1!
1%
#338230000000
0!
0%
#338235000000
1!
1%
#338240000000
0!
0%
#338245000000
1!
1%
#338250000000
0!
0%
#338255000000
1!
1%
#338260000000
0!
0%
#338265000000
1!
1%
#338270000000
0!
0%
#338275000000
1!
1%
#338280000000
0!
0%
#338285000000
1!
1%
#338290000000
0!
0%
#338295000000
1!
1%
#338300000000
0!
0%
#338305000000
1!
1%
#338310000000
0!
0%
#338315000000
1!
1%
#338320000000
0!
0%
#338325000000
1!
1%
#338330000000
0!
0%
#338335000000
1!
1%
#338340000000
0!
0%
#338345000000
1!
1%
#338350000000
0!
0%
#338355000000
1!
1%
#338360000000
0!
0%
#338365000000
1!
1%
#338370000000
0!
0%
#338375000000
1!
1%
#338380000000
0!
0%
#338385000000
1!
1%
#338390000000
0!
0%
#338395000000
1!
1%
#338400000000
0!
0%
#338405000000
1!
1%
#338410000000
0!
0%
#338415000000
1!
1%
#338420000000
0!
0%
#338425000000
1!
1%
#338430000000
0!
0%
#338435000000
1!
1%
#338440000000
0!
0%
#338445000000
1!
1%
#338450000000
0!
0%
#338455000000
1!
1%
#338460000000
0!
0%
#338465000000
1!
1%
#338470000000
0!
0%
#338475000000
1!
1%
#338480000000
0!
0%
#338485000000
1!
1%
#338490000000
0!
0%
#338495000000
1!
1%
#338500000000
0!
0%
#338505000000
1!
1%
#338510000000
0!
0%
#338515000000
1!
1%
#338520000000
0!
0%
#338525000000
1!
1%
#338530000000
0!
0%
#338535000000
1!
1%
#338540000000
0!
0%
#338545000000
1!
1%
#338550000000
0!
0%
#338555000000
1!
1%
#338560000000
0!
0%
#338565000000
1!
1%
#338570000000
0!
0%
#338575000000
1!
1%
#338580000000
0!
0%
#338585000000
1!
1%
#338590000000
0!
0%
#338595000000
1!
1%
#338600000000
0!
0%
#338605000000
1!
1%
#338610000000
0!
0%
#338615000000
1!
1%
#338620000000
0!
0%
#338625000000
1!
1%
#338630000000
0!
0%
#338635000000
1!
1%
#338640000000
0!
0%
#338645000000
1!
1%
#338650000000
0!
0%
#338655000000
1!
1%
#338660000000
0!
0%
#338665000000
1!
1%
#338670000000
0!
0%
#338675000000
1!
1%
#338680000000
0!
0%
#338685000000
1!
1%
#338690000000
0!
0%
#338695000000
1!
1%
#338700000000
0!
0%
#338705000000
1!
1%
#338710000000
0!
0%
#338715000000
1!
1%
#338720000000
0!
0%
#338725000000
1!
1%
#338730000000
0!
0%
#338735000000
1!
1%
#338740000000
0!
0%
#338745000000
1!
1%
#338750000000
0!
0%
#338755000000
1!
1%
#338760000000
0!
0%
#338765000000
1!
1%
#338770000000
0!
0%
#338775000000
1!
1%
#338780000000
0!
0%
#338785000000
1!
1%
#338790000000
0!
0%
#338795000000
1!
1%
#338800000000
0!
0%
#338805000000
1!
1%
#338810000000
0!
0%
#338815000000
1!
1%
#338820000000
0!
0%
#338825000000
1!
1%
#338830000000
0!
0%
#338835000000
1!
1%
#338840000000
0!
0%
#338845000000
1!
1%
#338850000000
0!
0%
#338855000000
1!
1%
#338860000000
0!
0%
#338865000000
1!
1%
#338870000000
0!
0%
#338875000000
1!
1%
#338880000000
0!
0%
#338885000000
1!
1%
#338890000000
0!
0%
#338895000000
1!
1%
#338900000000
0!
0%
#338905000000
1!
1%
#338910000000
0!
0%
#338915000000
1!
1%
#338920000000
0!
0%
#338925000000
1!
1%
#338930000000
0!
0%
#338935000000
1!
1%
#338940000000
0!
0%
#338945000000
1!
1%
#338950000000
0!
0%
#338955000000
1!
1%
#338960000000
0!
0%
#338965000000
1!
1%
#338970000000
0!
0%
#338975000000
1!
1%
#338980000000
0!
0%
#338985000000
1!
1%
#338990000000
0!
0%
#338995000000
1!
1%
#339000000000
0!
0%
#339005000000
1!
1%
#339010000000
0!
0%
#339015000000
1!
1%
#339020000000
0!
0%
#339025000000
1!
1%
#339030000000
0!
0%
#339035000000
1!
1%
#339040000000
0!
0%
#339045000000
1!
1%
#339050000000
0!
0%
#339055000000
1!
1%
#339060000000
0!
0%
#339065000000
1!
1%
#339070000000
0!
0%
#339075000000
1!
1%
#339080000000
0!
0%
#339085000000
1!
1%
#339090000000
0!
0%
#339095000000
1!
1%
#339100000000
0!
0%
#339105000000
1!
1%
#339110000000
0!
0%
#339115000000
1!
1%
#339120000000
0!
0%
#339125000000
1!
1%
#339130000000
0!
0%
#339135000000
1!
1%
#339140000000
0!
0%
#339145000000
1!
1%
#339150000000
0!
0%
#339155000000
1!
1%
#339160000000
0!
0%
#339165000000
1!
1%
#339170000000
0!
0%
#339175000000
1!
1%
#339180000000
0!
0%
#339185000000
1!
1%
#339190000000
0!
0%
#339195000000
1!
1%
#339200000000
0!
0%
#339205000000
1!
1%
#339210000000
0!
0%
#339215000000
1!
1%
#339220000000
0!
0%
#339225000000
1!
1%
#339230000000
0!
0%
#339235000000
1!
1%
#339240000000
0!
0%
#339245000000
1!
1%
#339250000000
0!
0%
#339255000000
1!
1%
#339260000000
0!
0%
#339265000000
1!
1%
#339270000000
0!
0%
#339275000000
1!
1%
#339280000000
0!
0%
#339285000000
1!
1%
#339290000000
0!
0%
#339295000000
1!
1%
#339300000000
0!
0%
#339305000000
1!
1%
#339310000000
0!
0%
#339315000000
1!
1%
#339320000000
0!
0%
#339325000000
1!
1%
#339330000000
0!
0%
#339335000000
1!
1%
#339340000000
0!
0%
#339345000000
1!
1%
#339350000000
0!
0%
#339355000000
1!
1%
#339360000000
0!
0%
#339365000000
1!
1%
#339370000000
0!
0%
#339375000000
1!
1%
#339380000000
0!
0%
#339385000000
1!
1%
#339390000000
0!
0%
#339395000000
1!
1%
#339400000000
0!
0%
#339405000000
1!
1%
#339410000000
0!
0%
#339415000000
1!
1%
#339420000000
0!
0%
#339425000000
1!
1%
#339430000000
0!
0%
#339435000000
1!
1%
#339440000000
0!
0%
#339445000000
1!
1%
#339450000000
0!
0%
#339455000000
1!
1%
#339460000000
0!
0%
#339465000000
1!
1%
#339470000000
0!
0%
#339475000000
1!
1%
#339480000000
0!
0%
#339485000000
1!
1%
#339490000000
0!
0%
#339495000000
1!
1%
#339500000000
0!
0%
#339505000000
1!
1%
#339510000000
0!
0%
#339515000000
1!
1%
#339520000000
0!
0%
#339525000000
1!
1%
#339530000000
0!
0%
#339535000000
1!
1%
#339540000000
0!
0%
#339545000000
1!
1%
#339550000000
0!
0%
#339555000000
1!
1%
#339560000000
0!
0%
#339565000000
1!
1%
#339570000000
0!
0%
#339575000000
1!
1%
#339580000000
0!
0%
#339585000000
1!
1%
#339590000000
0!
0%
#339595000000
1!
1%
#339600000000
0!
0%
#339605000000
1!
1%
#339610000000
0!
0%
#339615000000
1!
1%
#339620000000
0!
0%
#339625000000
1!
1%
#339630000000
0!
0%
#339635000000
1!
1%
#339640000000
0!
0%
#339645000000
1!
1%
#339650000000
0!
0%
#339655000000
1!
1%
#339660000000
0!
0%
#339665000000
1!
1%
#339670000000
0!
0%
#339675000000
1!
1%
#339680000000
0!
0%
#339685000000
1!
1%
#339690000000
0!
0%
#339695000000
1!
1%
#339700000000
0!
0%
#339705000000
1!
1%
#339710000000
0!
0%
#339715000000
1!
1%
#339720000000
0!
0%
#339725000000
1!
1%
#339730000000
0!
0%
#339735000000
1!
1%
#339740000000
0!
0%
#339745000000
1!
1%
#339750000000
0!
0%
#339755000000
1!
1%
#339760000000
0!
0%
#339765000000
1!
1%
#339770000000
0!
0%
#339775000000
1!
1%
#339780000000
0!
0%
#339785000000
1!
1%
#339790000000
0!
0%
#339795000000
1!
1%
#339800000000
0!
0%
#339805000000
1!
1%
#339810000000
0!
0%
#339815000000
1!
1%
#339820000000
0!
0%
#339825000000
1!
1%
#339830000000
0!
0%
#339835000000
1!
1%
#339840000000
0!
0%
#339845000000
1!
1%
#339850000000
0!
0%
#339855000000
1!
1%
#339860000000
0!
0%
#339865000000
1!
1%
#339870000000
0!
0%
#339875000000
1!
1%
#339880000000
0!
0%
#339885000000
1!
1%
#339890000000
0!
0%
#339895000000
1!
1%
#339900000000
0!
0%
#339905000000
1!
1%
#339910000000
0!
0%
#339915000000
1!
1%
#339920000000
0!
0%
#339925000000
1!
1%
#339930000000
0!
0%
#339935000000
1!
1%
#339940000000
0!
0%
#339945000000
1!
1%
#339950000000
0!
0%
#339955000000
1!
1%
#339960000000
0!
0%
#339965000000
1!
1%
#339970000000
0!
0%
#339975000000
1!
1%
#339980000000
0!
0%
#339985000000
1!
1%
#339990000000
0!
0%
#339995000000
1!
1%
#340000000000
0!
0%
#340005000000
1!
1%
#340010000000
0!
0%
#340015000000
1!
1%
#340020000000
0!
0%
#340025000000
1!
1%
#340030000000
0!
0%
#340035000000
1!
1%
#340040000000
0!
0%
#340045000000
1!
1%
#340050000000
0!
0%
#340055000000
1!
1%
#340060000000
0!
0%
#340065000000
1!
1%
#340070000000
0!
0%
#340075000000
1!
1%
#340080000000
0!
0%
#340085000000
1!
1%
#340090000000
0!
0%
#340095000000
1!
1%
#340100000000
0!
0%
#340105000000
1!
1%
#340110000000
0!
0%
#340115000000
1!
1%
#340120000000
0!
0%
#340125000000
1!
1%
#340130000000
0!
0%
#340135000000
1!
1%
#340140000000
0!
0%
#340145000000
1!
1%
#340150000000
0!
0%
#340155000000
1!
1%
#340160000000
0!
0%
#340165000000
1!
1%
#340170000000
0!
0%
#340175000000
1!
1%
#340180000000
0!
0%
#340185000000
1!
1%
#340190000000
0!
0%
#340195000000
1!
1%
#340200000000
0!
0%
#340205000000
1!
1%
#340210000000
0!
0%
#340215000000
1!
1%
#340220000000
0!
0%
#340225000000
1!
1%
#340230000000
0!
0%
#340235000000
1!
1%
#340240000000
0!
0%
#340245000000
1!
1%
#340250000000
0!
0%
#340255000000
1!
1%
#340260000000
0!
0%
#340265000000
1!
1%
#340270000000
0!
0%
#340275000000
1!
1%
#340280000000
0!
0%
#340285000000
1!
1%
#340290000000
0!
0%
#340295000000
1!
1%
#340300000000
0!
0%
#340305000000
1!
1%
#340310000000
0!
0%
#340315000000
1!
1%
#340320000000
0!
0%
#340325000000
1!
1%
#340330000000
0!
0%
#340335000000
1!
1%
#340340000000
0!
0%
#340345000000
1!
1%
#340350000000
0!
0%
#340355000000
1!
1%
#340360000000
0!
0%
#340365000000
1!
1%
#340370000000
0!
0%
#340375000000
1!
1%
#340380000000
0!
0%
#340385000000
1!
1%
#340390000000
0!
0%
#340395000000
1!
1%
#340400000000
0!
0%
#340405000000
1!
1%
#340410000000
0!
0%
#340415000000
1!
1%
#340420000000
0!
0%
#340425000000
1!
1%
#340430000000
0!
0%
#340435000000
1!
1%
#340440000000
0!
0%
#340445000000
1!
1%
#340450000000
0!
0%
#340455000000
1!
1%
#340460000000
0!
0%
#340465000000
1!
1%
#340470000000
0!
0%
#340475000000
1!
1%
#340480000000
0!
0%
#340485000000
1!
1%
#340490000000
0!
0%
#340495000000
1!
1%
#340500000000
0!
0%
#340505000000
1!
1%
#340510000000
0!
0%
#340515000000
1!
1%
#340520000000
0!
0%
#340525000000
1!
1%
#340530000000
0!
0%
#340535000000
1!
1%
#340540000000
0!
0%
#340545000000
1!
1%
#340550000000
0!
0%
#340555000000
1!
1%
#340560000000
0!
0%
#340565000000
1!
1%
#340570000000
0!
0%
#340575000000
1!
1%
#340580000000
0!
0%
#340585000000
1!
1%
#340590000000
0!
0%
#340595000000
1!
1%
#340600000000
0!
0%
#340605000000
1!
1%
#340610000000
0!
0%
#340615000000
1!
1%
#340620000000
0!
0%
#340625000000
1!
1%
#340630000000
0!
0%
#340635000000
1!
1%
#340640000000
0!
0%
#340645000000
1!
1%
#340650000000
0!
0%
#340655000000
1!
1%
#340660000000
0!
0%
#340665000000
1!
1%
#340670000000
0!
0%
#340675000000
1!
1%
#340680000000
0!
0%
#340685000000
1!
1%
#340690000000
0!
0%
#340695000000
1!
1%
#340700000000
0!
0%
#340705000000
1!
1%
#340710000000
0!
0%
#340715000000
1!
1%
#340720000000
0!
0%
#340725000000
1!
1%
#340730000000
0!
0%
#340735000000
1!
1%
#340740000000
0!
0%
#340745000000
1!
1%
#340750000000
0!
0%
#340755000000
1!
1%
#340760000000
0!
0%
#340765000000
1!
1%
#340770000000
0!
0%
#340775000000
1!
1%
#340780000000
0!
0%
#340785000000
1!
1%
#340790000000
0!
0%
#340795000000
1!
1%
#340800000000
0!
0%
#340805000000
1!
1%
#340810000000
0!
0%
#340815000000
1!
1%
#340820000000
0!
0%
#340825000000
1!
1%
#340830000000
0!
0%
#340835000000
1!
1%
#340840000000
0!
0%
#340845000000
1!
1%
#340850000000
0!
0%
#340855000000
1!
1%
#340860000000
0!
0%
#340865000000
1!
1%
#340870000000
0!
0%
#340875000000
1!
1%
#340880000000
0!
0%
#340885000000
1!
1%
#340890000000
0!
0%
#340895000000
1!
1%
#340900000000
0!
0%
#340905000000
1!
1%
#340910000000
0!
0%
#340915000000
1!
1%
#340920000000
0!
0%
#340925000000
1!
1%
#340930000000
0!
0%
#340935000000
1!
1%
#340940000000
0!
0%
#340945000000
1!
1%
#340950000000
0!
0%
#340955000000
1!
1%
#340960000000
0!
0%
#340965000000
1!
1%
#340970000000
0!
0%
#340975000000
1!
1%
#340980000000
0!
0%
#340985000000
1!
1%
#340990000000
0!
0%
#340995000000
1!
1%
#341000000000
0!
0%
#341005000000
1!
1%
#341010000000
0!
0%
#341015000000
1!
1%
#341020000000
0!
0%
#341025000000
1!
1%
#341030000000
0!
0%
#341035000000
1!
1%
#341040000000
0!
0%
#341045000000
1!
1%
#341050000000
0!
0%
#341055000000
1!
1%
#341060000000
0!
0%
#341065000000
1!
1%
#341070000000
0!
0%
#341075000000
1!
1%
#341080000000
0!
0%
#341085000000
1!
1%
#341090000000
0!
0%
#341095000000
1!
1%
#341100000000
0!
0%
#341105000000
1!
1%
#341110000000
0!
0%
#341115000000
1!
1%
#341120000000
0!
0%
#341125000000
1!
1%
#341130000000
0!
0%
#341135000000
1!
1%
#341140000000
0!
0%
#341145000000
1!
1%
#341150000000
0!
0%
#341155000000
1!
1%
#341160000000
0!
0%
#341165000000
1!
1%
#341170000000
0!
0%
#341175000000
1!
1%
#341180000000
0!
0%
#341185000000
1!
1%
#341190000000
0!
0%
#341195000000
1!
1%
#341200000000
0!
0%
#341205000000
1!
1%
#341210000000
0!
0%
#341215000000
1!
1%
#341220000000
0!
0%
#341225000000
1!
1%
#341230000000
0!
0%
#341235000000
1!
1%
#341240000000
0!
0%
#341245000000
1!
1%
#341250000000
0!
0%
#341255000000
1!
1%
#341260000000
0!
0%
#341265000000
1!
1%
#341270000000
0!
0%
#341275000000
1!
1%
#341280000000
0!
0%
#341285000000
1!
1%
#341290000000
0!
0%
#341295000000
1!
1%
#341300000000
0!
0%
#341305000000
1!
1%
#341310000000
0!
0%
#341315000000
1!
1%
#341320000000
0!
0%
#341325000000
1!
1%
#341330000000
0!
0%
#341335000000
1!
1%
#341340000000
0!
0%
#341345000000
1!
1%
#341350000000
0!
0%
#341355000000
1!
1%
#341360000000
0!
0%
#341365000000
1!
1%
#341370000000
0!
0%
#341375000000
1!
1%
#341380000000
0!
0%
#341385000000
1!
1%
#341390000000
0!
0%
#341395000000
1!
1%
#341400000000
0!
0%
#341405000000
1!
1%
#341410000000
0!
0%
#341415000000
1!
1%
#341420000000
0!
0%
#341425000000
1!
1%
#341430000000
0!
0%
#341435000000
1!
1%
#341440000000
0!
0%
#341445000000
1!
1%
#341450000000
0!
0%
#341455000000
1!
1%
#341460000000
0!
0%
#341465000000
1!
1%
#341470000000
0!
0%
#341475000000
1!
1%
#341480000000
0!
0%
#341485000000
1!
1%
#341490000000
0!
0%
#341495000000
1!
1%
#341500000000
0!
0%
#341505000000
1!
1%
#341510000000
0!
0%
#341515000000
1!
1%
#341520000000
0!
0%
#341525000000
1!
1%
#341530000000
0!
0%
#341535000000
1!
1%
#341540000000
0!
0%
#341545000000
1!
1%
#341550000000
0!
0%
#341555000000
1!
1%
#341560000000
0!
0%
#341565000000
1!
1%
#341570000000
0!
0%
#341575000000
1!
1%
#341580000000
0!
0%
#341585000000
1!
1%
#341590000000
0!
0%
#341595000000
1!
1%
#341600000000
0!
0%
#341605000000
1!
1%
#341610000000
0!
0%
#341615000000
1!
1%
#341620000000
0!
0%
#341625000000
1!
1%
#341630000000
0!
0%
#341635000000
1!
1%
#341640000000
0!
0%
#341645000000
1!
1%
#341650000000
0!
0%
#341655000000
1!
1%
#341660000000
0!
0%
#341665000000
1!
1%
#341670000000
0!
0%
#341675000000
1!
1%
#341680000000
0!
0%
#341685000000
1!
1%
#341690000000
0!
0%
#341695000000
1!
1%
#341700000000
0!
0%
#341705000000
1!
1%
#341710000000
0!
0%
#341715000000
1!
1%
#341720000000
0!
0%
#341725000000
1!
1%
#341730000000
0!
0%
#341735000000
1!
1%
#341740000000
0!
0%
#341745000000
1!
1%
#341750000000
0!
0%
#341755000000
1!
1%
#341760000000
0!
0%
#341765000000
1!
1%
#341770000000
0!
0%
#341775000000
1!
1%
#341780000000
0!
0%
#341785000000
1!
1%
#341790000000
0!
0%
#341795000000
1!
1%
#341800000000
0!
0%
#341805000000
1!
1%
#341810000000
0!
0%
#341815000000
1!
1%
#341820000000
0!
0%
#341825000000
1!
1%
#341830000000
0!
0%
#341835000000
1!
1%
#341840000000
0!
0%
#341845000000
1!
1%
#341850000000
0!
0%
#341855000000
1!
1%
#341860000000
0!
0%
#341865000000
1!
1%
#341870000000
0!
0%
#341875000000
1!
1%
#341880000000
0!
0%
#341885000000
1!
1%
#341890000000
0!
0%
#341895000000
1!
1%
#341900000000
0!
0%
#341905000000
1!
1%
#341910000000
0!
0%
#341915000000
1!
1%
#341920000000
0!
0%
#341925000000
1!
1%
#341930000000
0!
0%
#341935000000
1!
1%
#341940000000
0!
0%
#341945000000
1!
1%
#341950000000
0!
0%
#341955000000
1!
1%
#341960000000
0!
0%
#341965000000
1!
1%
#341970000000
0!
0%
#341975000000
1!
1%
#341980000000
0!
0%
#341985000000
1!
1%
#341990000000
0!
0%
#341995000000
1!
1%
#342000000000
0!
0%
#342005000000
1!
1%
#342010000000
0!
0%
#342015000000
1!
1%
#342020000000
0!
0%
#342025000000
1!
1%
#342030000000
0!
0%
#342035000000
1!
1%
#342040000000
0!
0%
#342045000000
1!
1%
#342050000000
0!
0%
#342055000000
1!
1%
#342060000000
0!
0%
#342065000000
1!
1%
#342070000000
0!
0%
#342075000000
1!
1%
#342080000000
0!
0%
#342085000000
1!
1%
#342090000000
0!
0%
#342095000000
1!
1%
#342100000000
0!
0%
#342105000000
1!
1%
#342110000000
0!
0%
#342115000000
1!
1%
#342120000000
0!
0%
#342125000000
1!
1%
#342130000000
0!
0%
#342135000000
1!
1%
#342140000000
0!
0%
#342145000000
1!
1%
#342150000000
0!
0%
#342155000000
1!
1%
#342160000000
0!
0%
#342165000000
1!
1%
#342170000000
0!
0%
#342175000000
1!
1%
#342180000000
0!
0%
#342185000000
1!
1%
#342190000000
0!
0%
#342195000000
1!
1%
#342200000000
0!
0%
#342205000000
1!
1%
#342210000000
0!
0%
#342215000000
1!
1%
#342220000000
0!
0%
#342225000000
1!
1%
#342230000000
0!
0%
#342235000000
1!
1%
#342240000000
0!
0%
#342245000000
1!
1%
#342250000000
0!
0%
#342255000000
1!
1%
#342260000000
0!
0%
#342265000000
1!
1%
#342270000000
0!
0%
#342275000000
1!
1%
#342280000000
0!
0%
#342285000000
1!
1%
#342290000000
0!
0%
#342295000000
1!
1%
#342300000000
0!
0%
#342305000000
1!
1%
#342310000000
0!
0%
#342315000000
1!
1%
#342320000000
0!
0%
#342325000000
1!
1%
#342330000000
0!
0%
#342335000000
1!
1%
#342340000000
0!
0%
#342345000000
1!
1%
#342350000000
0!
0%
#342355000000
1!
1%
#342360000000
0!
0%
#342365000000
1!
1%
#342370000000
0!
0%
#342375000000
1!
1%
#342380000000
0!
0%
#342385000000
1!
1%
#342390000000
0!
0%
#342395000000
1!
1%
#342400000000
0!
0%
#342405000000
1!
1%
#342410000000
0!
0%
#342415000000
1!
1%
#342420000000
0!
0%
#342425000000
1!
1%
#342430000000
0!
0%
#342435000000
1!
1%
#342440000000
0!
0%
#342445000000
1!
1%
#342450000000
0!
0%
#342455000000
1!
1%
#342460000000
0!
0%
#342465000000
1!
1%
#342470000000
0!
0%
#342475000000
1!
1%
#342480000000
0!
0%
#342485000000
1!
1%
#342490000000
0!
0%
#342495000000
1!
1%
#342500000000
0!
0%
#342505000000
1!
1%
#342510000000
0!
0%
#342515000000
1!
1%
#342520000000
0!
0%
#342525000000
1!
1%
#342530000000
0!
0%
#342535000000
1!
1%
#342540000000
0!
0%
#342545000000
1!
1%
#342550000000
0!
0%
#342555000000
1!
1%
#342560000000
0!
0%
#342565000000
1!
1%
#342570000000
0!
0%
#342575000000
1!
1%
#342580000000
0!
0%
#342585000000
1!
1%
#342590000000
0!
0%
#342595000000
1!
1%
#342600000000
0!
0%
#342605000000
1!
1%
#342610000000
0!
0%
#342615000000
1!
1%
#342620000000
0!
0%
#342625000000
1!
1%
#342630000000
0!
0%
#342635000000
1!
1%
#342640000000
0!
0%
#342645000000
1!
1%
#342650000000
0!
0%
#342655000000
1!
1%
#342660000000
0!
0%
#342665000000
1!
1%
#342670000000
0!
0%
#342675000000
1!
1%
#342680000000
0!
0%
#342685000000
1!
1%
#342690000000
0!
0%
#342695000000
1!
1%
#342700000000
0!
0%
#342705000000
1!
1%
#342710000000
0!
0%
#342715000000
1!
1%
#342720000000
0!
0%
#342725000000
1!
1%
#342730000000
0!
0%
#342735000000
1!
1%
#342740000000
0!
0%
#342745000000
1!
1%
#342750000000
0!
0%
#342755000000
1!
1%
#342760000000
0!
0%
#342765000000
1!
1%
#342770000000
0!
0%
#342775000000
1!
1%
#342780000000
0!
0%
#342785000000
1!
1%
#342790000000
0!
0%
#342795000000
1!
1%
#342800000000
0!
0%
#342805000000
1!
1%
#342810000000
0!
0%
#342815000000
1!
1%
#342820000000
0!
0%
#342825000000
1!
1%
#342830000000
0!
0%
#342835000000
1!
1%
#342840000000
0!
0%
#342845000000
1!
1%
#342850000000
0!
0%
#342855000000
1!
1%
#342860000000
0!
0%
#342865000000
1!
1%
#342870000000
0!
0%
#342875000000
1!
1%
#342880000000
0!
0%
#342885000000
1!
1%
#342890000000
0!
0%
#342895000000
1!
1%
#342900000000
0!
0%
#342905000000
1!
1%
#342910000000
0!
0%
#342915000000
1!
1%
#342920000000
0!
0%
#342925000000
1!
1%
#342930000000
0!
0%
#342935000000
1!
1%
#342940000000
0!
0%
#342945000000
1!
1%
#342950000000
0!
0%
#342955000000
1!
1%
#342960000000
0!
0%
#342965000000
1!
1%
#342970000000
0!
0%
#342975000000
1!
1%
#342980000000
0!
0%
#342985000000
1!
1%
#342990000000
0!
0%
#342995000000
1!
1%
#343000000000
0!
0%
#343005000000
1!
1%
#343010000000
0!
0%
#343015000000
1!
1%
#343020000000
0!
0%
#343025000000
1!
1%
#343030000000
0!
0%
#343035000000
1!
1%
#343040000000
0!
0%
#343045000000
1!
1%
#343050000000
0!
0%
#343055000000
1!
1%
#343060000000
0!
0%
#343065000000
1!
1%
#343070000000
0!
0%
#343075000000
1!
1%
#343080000000
0!
0%
#343085000000
1!
1%
#343090000000
0!
0%
#343095000000
1!
1%
#343100000000
0!
0%
#343105000000
1!
1%
#343110000000
0!
0%
#343115000000
1!
1%
#343120000000
0!
0%
#343125000000
1!
1%
#343130000000
0!
0%
#343135000000
1!
1%
#343140000000
0!
0%
#343145000000
1!
1%
#343150000000
0!
0%
#343155000000
1!
1%
#343160000000
0!
0%
#343165000000
1!
1%
#343170000000
0!
0%
#343175000000
1!
1%
#343180000000
0!
0%
#343185000000
1!
1%
#343190000000
0!
0%
#343195000000
1!
1%
#343200000000
0!
0%
#343205000000
1!
1%
#343210000000
0!
0%
#343215000000
1!
1%
#343220000000
0!
0%
#343225000000
1!
1%
#343230000000
0!
0%
#343235000000
1!
1%
#343240000000
0!
0%
#343245000000
1!
1%
#343250000000
0!
0%
#343255000000
1!
1%
#343260000000
0!
0%
#343265000000
1!
1%
#343270000000
0!
0%
#343275000000
1!
1%
#343280000000
0!
0%
#343285000000
1!
1%
#343290000000
0!
0%
#343295000000
1!
1%
#343300000000
0!
0%
#343305000000
1!
1%
#343310000000
0!
0%
#343315000000
1!
1%
#343320000000
0!
0%
#343325000000
1!
1%
#343330000000
0!
0%
#343335000000
1!
1%
#343340000000
0!
0%
#343345000000
1!
1%
#343350000000
0!
0%
#343355000000
1!
1%
#343360000000
0!
0%
#343365000000
1!
1%
#343370000000
0!
0%
#343375000000
1!
1%
#343380000000
0!
0%
#343385000000
1!
1%
#343390000000
0!
0%
#343395000000
1!
1%
#343400000000
0!
0%
#343405000000
1!
1%
#343410000000
0!
0%
#343415000000
1!
1%
#343420000000
0!
0%
#343425000000
1!
1%
#343430000000
0!
0%
#343435000000
1!
1%
#343440000000
0!
0%
#343445000000
1!
1%
#343450000000
0!
0%
#343455000000
1!
1%
#343460000000
0!
0%
#343465000000
1!
1%
#343470000000
0!
0%
#343475000000
1!
1%
#343480000000
0!
0%
#343485000000
1!
1%
#343490000000
0!
0%
#343495000000
1!
1%
#343500000000
0!
0%
#343505000000
1!
1%
#343510000000
0!
0%
#343515000000
1!
1%
#343520000000
0!
0%
#343525000000
1!
1%
#343530000000
0!
0%
#343535000000
1!
1%
#343540000000
0!
0%
#343545000000
1!
1%
#343550000000
0!
0%
#343555000000
1!
1%
#343560000000
0!
0%
#343565000000
1!
1%
#343570000000
0!
0%
#343575000000
1!
1%
#343580000000
0!
0%
#343585000000
1!
1%
#343590000000
0!
0%
#343595000000
1!
1%
#343600000000
0!
0%
#343605000000
1!
1%
#343610000000
0!
0%
#343615000000
1!
1%
#343620000000
0!
0%
#343625000000
1!
1%
#343630000000
0!
0%
#343635000000
1!
1%
#343640000000
0!
0%
#343645000000
1!
1%
#343650000000
0!
0%
#343655000000
1!
1%
#343660000000
0!
0%
#343665000000
1!
1%
#343670000000
0!
0%
#343675000000
1!
1%
#343680000000
0!
0%
#343685000000
1!
1%
#343690000000
0!
0%
#343695000000
1!
1%
#343700000000
0!
0%
#343705000000
1!
1%
#343710000000
0!
0%
#343715000000
1!
1%
#343720000000
0!
0%
#343725000000
1!
1%
#343730000000
0!
0%
#343735000000
1!
1%
#343740000000
0!
0%
#343745000000
1!
1%
#343750000000
0!
0%
#343755000000
1!
1%
#343760000000
0!
0%
#343765000000
1!
1%
#343770000000
0!
0%
#343775000000
1!
1%
#343780000000
0!
0%
#343785000000
1!
1%
#343790000000
0!
0%
#343795000000
1!
1%
#343800000000
0!
0%
#343805000000
1!
1%
#343810000000
0!
0%
#343815000000
1!
1%
#343820000000
0!
0%
#343825000000
1!
1%
#343830000000
0!
0%
#343835000000
1!
1%
#343840000000
0!
0%
#343845000000
1!
1%
#343850000000
0!
0%
#343855000000
1!
1%
#343860000000
0!
0%
#343865000000
1!
1%
#343870000000
0!
0%
#343875000000
1!
1%
#343880000000
0!
0%
#343885000000
1!
1%
#343890000000
0!
0%
#343895000000
1!
1%
#343900000000
0!
0%
#343905000000
1!
1%
#343910000000
0!
0%
#343915000000
1!
1%
#343920000000
0!
0%
#343925000000
1!
1%
#343930000000
0!
0%
#343935000000
1!
1%
#343940000000
0!
0%
#343945000000
1!
1%
#343950000000
0!
0%
#343955000000
1!
1%
#343960000000
0!
0%
#343965000000
1!
1%
#343970000000
0!
0%
#343975000000
1!
1%
#343980000000
0!
0%
#343985000000
1!
1%
#343990000000
0!
0%
#343995000000
1!
1%
#344000000000
0!
0%
#344005000000
1!
1%
#344010000000
0!
0%
#344015000000
1!
1%
#344020000000
0!
0%
#344025000000
1!
1%
#344030000000
0!
0%
#344035000000
1!
1%
#344040000000
0!
0%
#344045000000
1!
1%
#344050000000
0!
0%
#344055000000
1!
1%
#344060000000
0!
0%
#344065000000
1!
1%
#344070000000
0!
0%
#344075000000
1!
1%
#344080000000
0!
0%
#344085000000
1!
1%
#344090000000
0!
0%
#344095000000
1!
1%
#344100000000
0!
0%
#344105000000
1!
1%
#344110000000
0!
0%
#344115000000
1!
1%
#344120000000
0!
0%
#344125000000
1!
1%
#344130000000
0!
0%
#344135000000
1!
1%
#344140000000
0!
0%
#344145000000
1!
1%
#344150000000
0!
0%
#344155000000
1!
1%
#344160000000
0!
0%
#344165000000
1!
1%
#344170000000
0!
0%
#344175000000
1!
1%
#344180000000
0!
0%
#344185000000
1!
1%
#344190000000
0!
0%
#344195000000
1!
1%
#344200000000
0!
0%
#344205000000
1!
1%
#344210000000
0!
0%
#344215000000
1!
1%
#344220000000
0!
0%
#344225000000
1!
1%
#344230000000
0!
0%
#344235000000
1!
1%
#344240000000
0!
0%
#344245000000
1!
1%
#344250000000
0!
0%
#344255000000
1!
1%
#344260000000
0!
0%
#344265000000
1!
1%
#344270000000
0!
0%
#344275000000
1!
1%
#344280000000
0!
0%
#344285000000
1!
1%
#344290000000
0!
0%
#344295000000
1!
1%
#344300000000
0!
0%
#344305000000
1!
1%
#344310000000
0!
0%
#344315000000
1!
1%
#344320000000
0!
0%
#344325000000
1!
1%
#344330000000
0!
0%
#344335000000
1!
1%
#344340000000
0!
0%
#344345000000
1!
1%
#344350000000
0!
0%
#344355000000
1!
1%
#344360000000
0!
0%
#344365000000
1!
1%
#344370000000
0!
0%
#344375000000
1!
1%
#344380000000
0!
0%
#344385000000
1!
1%
#344390000000
0!
0%
#344395000000
1!
1%
#344400000000
0!
0%
#344405000000
1!
1%
#344410000000
0!
0%
#344415000000
1!
1%
#344420000000
0!
0%
#344425000000
1!
1%
#344430000000
0!
0%
#344435000000
1!
1%
#344440000000
0!
0%
#344445000000
1!
1%
#344450000000
0!
0%
#344455000000
1!
1%
#344460000000
0!
0%
#344465000000
1!
1%
#344470000000
0!
0%
#344475000000
1!
1%
#344480000000
0!
0%
#344485000000
1!
1%
#344490000000
0!
0%
#344495000000
1!
1%
#344500000000
0!
0%
#344505000000
1!
1%
#344510000000
0!
0%
#344515000000
1!
1%
#344520000000
0!
0%
#344525000000
1!
1%
#344530000000
0!
0%
#344535000000
1!
1%
#344540000000
0!
0%
#344545000000
1!
1%
#344550000000
0!
0%
#344555000000
1!
1%
#344560000000
0!
0%
#344565000000
1!
1%
#344570000000
0!
0%
#344575000000
1!
1%
#344580000000
0!
0%
#344585000000
1!
1%
#344590000000
0!
0%
#344595000000
1!
1%
#344600000000
0!
0%
#344605000000
1!
1%
#344610000000
0!
0%
#344615000000
1!
1%
#344620000000
0!
0%
#344625000000
1!
1%
#344630000000
0!
0%
#344635000000
1!
1%
#344640000000
0!
0%
#344645000000
1!
1%
#344650000000
0!
0%
#344655000000
1!
1%
#344660000000
0!
0%
#344665000000
1!
1%
#344670000000
0!
0%
#344675000000
1!
1%
#344680000000
0!
0%
#344685000000
1!
1%
#344690000000
0!
0%
#344695000000
1!
1%
#344700000000
0!
0%
#344705000000
1!
1%
#344710000000
0!
0%
#344715000000
1!
1%
#344720000000
0!
0%
#344725000000
1!
1%
#344730000000
0!
0%
#344735000000
1!
1%
#344740000000
0!
0%
#344745000000
1!
1%
#344750000000
0!
0%
#344755000000
1!
1%
#344760000000
0!
0%
#344765000000
1!
1%
#344770000000
0!
0%
#344775000000
1!
1%
#344780000000
0!
0%
#344785000000
1!
1%
#344790000000
0!
0%
#344795000000
1!
1%
#344800000000
0!
0%
#344805000000
1!
1%
#344810000000
0!
0%
#344815000000
1!
1%
#344820000000
0!
0%
#344825000000
1!
1%
#344830000000
0!
0%
#344835000000
1!
1%
#344840000000
0!
0%
#344845000000
1!
1%
#344850000000
0!
0%
#344855000000
1!
1%
#344860000000
0!
0%
#344865000000
1!
1%
#344870000000
0!
0%
#344875000000
1!
1%
#344880000000
0!
0%
#344885000000
1!
1%
#344890000000
0!
0%
#344895000000
1!
1%
#344900000000
0!
0%
#344905000000
1!
1%
#344910000000
0!
0%
#344915000000
1!
1%
#344920000000
0!
0%
#344925000000
1!
1%
#344930000000
0!
0%
#344935000000
1!
1%
#344940000000
0!
0%
#344945000000
1!
1%
#344950000000
0!
0%
#344955000000
1!
1%
#344960000000
0!
0%
#344965000000
1!
1%
#344970000000
0!
0%
#344975000000
1!
1%
#344980000000
0!
0%
#344985000000
1!
1%
#344990000000
0!
0%
#344995000000
1!
1%
#345000000000
0!
0%
#345005000000
1!
1%
#345010000000
0!
0%
#345015000000
1!
1%
#345020000000
0!
0%
#345025000000
1!
1%
#345030000000
0!
0%
#345035000000
1!
1%
#345040000000
0!
0%
#345045000000
1!
1%
#345050000000
0!
0%
#345055000000
1!
1%
#345060000000
0!
0%
#345065000000
1!
1%
#345070000000
0!
0%
#345075000000
1!
1%
#345080000000
0!
0%
#345085000000
1!
1%
#345090000000
0!
0%
#345095000000
1!
1%
#345100000000
0!
0%
#345105000000
1!
1%
#345110000000
0!
0%
#345115000000
1!
1%
#345120000000
0!
0%
#345125000000
1!
1%
#345130000000
0!
0%
#345135000000
1!
1%
#345140000000
0!
0%
#345145000000
1!
1%
#345150000000
0!
0%
#345155000000
1!
1%
#345160000000
0!
0%
#345165000000
1!
1%
#345170000000
0!
0%
#345175000000
1!
1%
#345180000000
0!
0%
#345185000000
1!
1%
#345190000000
0!
0%
#345195000000
1!
1%
#345200000000
0!
0%
#345205000000
1!
1%
#345210000000
0!
0%
#345215000000
1!
1%
#345220000000
0!
0%
#345225000000
1!
1%
#345230000000
0!
0%
#345235000000
1!
1%
#345240000000
0!
0%
#345245000000
1!
1%
#345250000000
0!
0%
#345255000000
1!
1%
#345260000000
0!
0%
#345265000000
1!
1%
#345270000000
0!
0%
#345275000000
1!
1%
#345280000000
0!
0%
#345285000000
1!
1%
#345290000000
0!
0%
#345295000000
1!
1%
#345300000000
0!
0%
#345305000000
1!
1%
#345310000000
0!
0%
#345315000000
1!
1%
#345320000000
0!
0%
#345325000000
1!
1%
#345330000000
0!
0%
#345335000000
1!
1%
#345340000000
0!
0%
#345345000000
1!
1%
#345350000000
0!
0%
#345355000000
1!
1%
#345360000000
0!
0%
#345365000000
1!
1%
#345370000000
0!
0%
#345375000000
1!
1%
#345380000000
0!
0%
#345385000000
1!
1%
#345390000000
0!
0%
#345395000000
1!
1%
#345400000000
0!
0%
#345405000000
1!
1%
#345410000000
0!
0%
#345415000000
1!
1%
#345420000000
0!
0%
#345425000000
1!
1%
#345430000000
0!
0%
#345435000000
1!
1%
#345440000000
0!
0%
#345445000000
1!
1%
#345450000000
0!
0%
#345455000000
1!
1%
#345460000000
0!
0%
#345465000000
1!
1%
#345470000000
0!
0%
#345475000000
1!
1%
#345480000000
0!
0%
#345485000000
1!
1%
#345490000000
0!
0%
#345495000000
1!
1%
#345500000000
0!
0%
#345505000000
1!
1%
#345510000000
0!
0%
#345515000000
1!
1%
#345520000000
0!
0%
#345525000000
1!
1%
#345530000000
0!
0%
#345535000000
1!
1%
#345540000000
0!
0%
#345545000000
1!
1%
#345550000000
0!
0%
#345555000000
1!
1%
#345560000000
0!
0%
#345565000000
1!
1%
#345570000000
0!
0%
#345575000000
1!
1%
#345580000000
0!
0%
#345585000000
1!
1%
#345590000000
0!
0%
#345595000000
1!
1%
#345600000000
0!
0%
#345605000000
1!
1%
#345610000000
0!
0%
#345615000000
1!
1%
#345620000000
0!
0%
#345625000000
1!
1%
#345630000000
0!
0%
#345635000000
1!
1%
#345640000000
0!
0%
#345645000000
1!
1%
#345650000000
0!
0%
#345655000000
1!
1%
#345660000000
0!
0%
#345665000000
1!
1%
#345670000000
0!
0%
#345675000000
1!
1%
#345680000000
0!
0%
#345685000000
1!
1%
#345690000000
0!
0%
#345695000000
1!
1%
#345700000000
0!
0%
#345705000000
1!
1%
#345710000000
0!
0%
#345715000000
1!
1%
#345720000000
0!
0%
#345725000000
1!
1%
#345730000000
0!
0%
#345735000000
1!
1%
#345740000000
0!
0%
#345745000000
1!
1%
#345750000000
0!
0%
#345755000000
1!
1%
#345760000000
0!
0%
#345765000000
1!
1%
#345770000000
0!
0%
#345775000000
1!
1%
#345780000000
0!
0%
#345785000000
1!
1%
#345790000000
0!
0%
#345795000000
1!
1%
#345800000000
0!
0%
#345805000000
1!
1%
#345810000000
0!
0%
#345815000000
1!
1%
#345820000000
0!
0%
#345825000000
1!
1%
#345830000000
0!
0%
#345835000000
1!
1%
#345840000000
0!
0%
#345845000000
1!
1%
#345850000000
0!
0%
#345855000000
1!
1%
#345860000000
0!
0%
#345865000000
1!
1%
#345870000000
0!
0%
#345875000000
1!
1%
#345880000000
0!
0%
#345885000000
1!
1%
#345890000000
0!
0%
#345895000000
1!
1%
#345900000000
0!
0%
#345905000000
1!
1%
#345910000000
0!
0%
#345915000000
1!
1%
#345920000000
0!
0%
#345925000000
1!
1%
#345930000000
0!
0%
#345935000000
1!
1%
#345940000000
0!
0%
#345945000000
1!
1%
#345950000000
0!
0%
#345955000000
1!
1%
#345960000000
0!
0%
#345965000000
1!
1%
#345970000000
0!
0%
#345975000000
1!
1%
#345980000000
0!
0%
#345985000000
1!
1%
#345990000000
0!
0%
#345995000000
1!
1%
#346000000000
0!
0%
#346005000000
1!
1%
#346010000000
0!
0%
#346015000000
1!
1%
#346020000000
0!
0%
#346025000000
1!
1%
#346030000000
0!
0%
#346035000000
1!
1%
#346040000000
0!
0%
#346045000000
1!
1%
#346050000000
0!
0%
#346055000000
1!
1%
#346060000000
0!
0%
#346065000000
1!
1%
#346070000000
0!
0%
#346075000000
1!
1%
#346080000000
0!
0%
#346085000000
1!
1%
#346090000000
0!
0%
#346095000000
1!
1%
#346100000000
0!
0%
#346105000000
1!
1%
#346110000000
0!
0%
#346115000000
1!
1%
#346120000000
0!
0%
#346125000000
1!
1%
#346130000000
0!
0%
#346135000000
1!
1%
#346140000000
0!
0%
#346145000000
1!
1%
#346150000000
0!
0%
#346155000000
1!
1%
#346160000000
0!
0%
#346165000000
1!
1%
#346170000000
0!
0%
#346175000000
1!
1%
#346180000000
0!
0%
#346185000000
1!
1%
#346190000000
0!
0%
#346195000000
1!
1%
#346200000000
0!
0%
#346205000000
1!
1%
#346210000000
0!
0%
#346215000000
1!
1%
#346220000000
0!
0%
#346225000000
1!
1%
#346230000000
0!
0%
#346235000000
1!
1%
#346240000000
0!
0%
#346245000000
1!
1%
#346250000000
0!
0%
#346255000000
1!
1%
#346260000000
0!
0%
#346265000000
1!
1%
#346270000000
0!
0%
#346275000000
1!
1%
#346280000000
0!
0%
#346285000000
1!
1%
#346290000000
0!
0%
#346295000000
1!
1%
#346300000000
0!
0%
#346305000000
1!
1%
#346310000000
0!
0%
#346315000000
1!
1%
#346320000000
0!
0%
#346325000000
1!
1%
#346330000000
0!
0%
#346335000000
1!
1%
#346340000000
0!
0%
#346345000000
1!
1%
#346350000000
0!
0%
#346355000000
1!
1%
#346360000000
0!
0%
#346365000000
1!
1%
#346370000000
0!
0%
#346375000000
1!
1%
#346380000000
0!
0%
#346385000000
1!
1%
#346390000000
0!
0%
#346395000000
1!
1%
#346400000000
0!
0%
#346405000000
1!
1%
#346410000000
0!
0%
#346415000000
1!
1%
#346420000000
0!
0%
#346425000000
1!
1%
#346430000000
0!
0%
#346435000000
1!
1%
#346440000000
0!
0%
#346445000000
1!
1%
#346450000000
0!
0%
#346455000000
1!
1%
#346460000000
0!
0%
#346465000000
1!
1%
#346470000000
0!
0%
#346475000000
1!
1%
#346480000000
0!
0%
#346485000000
1!
1%
#346490000000
0!
0%
#346495000000
1!
1%
#346500000000
0!
0%
#346505000000
1!
1%
#346510000000
0!
0%
#346515000000
1!
1%
#346520000000
0!
0%
#346525000000
1!
1%
#346530000000
0!
0%
#346535000000
1!
1%
#346540000000
0!
0%
#346545000000
1!
1%
#346550000000
0!
0%
#346555000000
1!
1%
#346560000000
0!
0%
#346565000000
1!
1%
#346570000000
0!
0%
#346575000000
1!
1%
#346580000000
0!
0%
#346585000000
1!
1%
#346590000000
0!
0%
#346595000000
1!
1%
#346600000000
0!
0%
#346605000000
1!
1%
#346610000000
0!
0%
#346615000000
1!
1%
#346620000000
0!
0%
#346625000000
1!
1%
#346630000000
0!
0%
#346635000000
1!
1%
#346640000000
0!
0%
#346645000000
1!
1%
#346650000000
0!
0%
#346655000000
1!
1%
#346660000000
0!
0%
#346665000000
1!
1%
#346670000000
0!
0%
#346675000000
1!
1%
#346680000000
0!
0%
#346685000000
1!
1%
#346690000000
0!
0%
#346695000000
1!
1%
#346700000000
0!
0%
#346705000000
1!
1%
#346710000000
0!
0%
#346715000000
1!
1%
#346720000000
0!
0%
#346725000000
1!
1%
#346730000000
0!
0%
#346735000000
1!
1%
#346740000000
0!
0%
#346745000000
1!
1%
#346750000000
0!
0%
#346755000000
1!
1%
#346760000000
0!
0%
#346765000000
1!
1%
#346770000000
0!
0%
#346775000000
1!
1%
#346780000000
0!
0%
#346785000000
1!
1%
#346790000000
0!
0%
#346795000000
1!
1%
#346800000000
0!
0%
#346805000000
1!
1%
#346810000000
0!
0%
#346815000000
1!
1%
#346820000000
0!
0%
#346825000000
1!
1%
#346830000000
0!
0%
#346835000000
1!
1%
#346840000000
0!
0%
#346845000000
1!
1%
#346850000000
0!
0%
#346855000000
1!
1%
#346860000000
0!
0%
#346865000000
1!
1%
#346870000000
0!
0%
#346875000000
1!
1%
#346880000000
0!
0%
#346885000000
1!
1%
#346890000000
0!
0%
#346895000000
1!
1%
#346900000000
0!
0%
#346905000000
1!
1%
#346910000000
0!
0%
#346915000000
1!
1%
#346920000000
0!
0%
#346925000000
1!
1%
#346930000000
0!
0%
#346935000000
1!
1%
#346940000000
0!
0%
#346945000000
1!
1%
#346950000000
0!
0%
#346955000000
1!
1%
#346960000000
0!
0%
#346965000000
1!
1%
#346970000000
0!
0%
#346975000000
1!
1%
#346980000000
0!
0%
#346985000000
1!
1%
#346990000000
0!
0%
#346995000000
1!
1%
#347000000000
0!
0%
#347005000000
1!
1%
#347010000000
0!
0%
#347015000000
1!
1%
#347020000000
0!
0%
#347025000000
1!
1%
#347030000000
0!
0%
#347035000000
1!
1%
#347040000000
0!
0%
#347045000000
1!
1%
#347050000000
0!
0%
#347055000000
1!
1%
#347060000000
0!
0%
#347065000000
1!
1%
#347070000000
0!
0%
#347075000000
1!
1%
#347080000000
0!
0%
#347085000000
1!
1%
#347090000000
0!
0%
#347095000000
1!
1%
#347100000000
0!
0%
#347105000000
1!
1%
#347110000000
0!
0%
#347115000000
1!
1%
#347120000000
0!
0%
#347125000000
1!
1%
#347130000000
0!
0%
#347135000000
1!
1%
#347140000000
0!
0%
#347145000000
1!
1%
#347150000000
0!
0%
#347155000000
1!
1%
#347160000000
0!
0%
#347165000000
1!
1%
#347170000000
0!
0%
#347175000000
1!
1%
#347180000000
0!
0%
#347185000000
1!
1%
#347190000000
0!
0%
#347195000000
1!
1%
#347200000000
0!
0%
#347205000000
1!
1%
#347210000000
0!
0%
#347215000000
1!
1%
#347220000000
0!
0%
#347225000000
1!
1%
#347230000000
0!
0%
#347235000000
1!
1%
#347240000000
0!
0%
#347245000000
1!
1%
#347250000000
0!
0%
#347255000000
1!
1%
#347260000000
0!
0%
#347265000000
1!
1%
#347270000000
0!
0%
#347275000000
1!
1%
#347280000000
0!
0%
#347285000000
1!
1%
#347290000000
0!
0%
#347295000000
1!
1%
#347300000000
0!
0%
#347305000000
1!
1%
#347310000000
0!
0%
#347315000000
1!
1%
#347320000000
0!
0%
#347325000000
1!
1%
#347330000000
0!
0%
#347335000000
1!
1%
#347340000000
0!
0%
#347345000000
1!
1%
#347350000000
0!
0%
#347355000000
1!
1%
#347360000000
0!
0%
#347365000000
1!
1%
#347370000000
0!
0%
#347375000000
1!
1%
#347380000000
0!
0%
#347385000000
1!
1%
#347390000000
0!
0%
#347395000000
1!
1%
#347400000000
0!
0%
#347405000000
1!
1%
#347410000000
0!
0%
#347415000000
1!
1%
#347420000000
0!
0%
#347425000000
1!
1%
#347430000000
0!
0%
#347435000000
1!
1%
#347440000000
0!
0%
#347445000000
1!
1%
#347450000000
0!
0%
#347455000000
1!
1%
#347460000000
0!
0%
#347465000000
1!
1%
#347470000000
0!
0%
#347475000000
1!
1%
#347480000000
0!
0%
#347485000000
1!
1%
#347490000000
0!
0%
#347495000000
1!
1%
#347500000000
0!
0%
#347505000000
1!
1%
#347510000000
0!
0%
#347515000000
1!
1%
#347520000000
0!
0%
#347525000000
1!
1%
#347530000000
0!
0%
#347535000000
1!
1%
#347540000000
0!
0%
#347545000000
1!
1%
#347550000000
0!
0%
#347555000000
1!
1%
#347560000000
0!
0%
#347565000000
1!
1%
#347570000000
0!
0%
#347575000000
1!
1%
#347580000000
0!
0%
#347585000000
1!
1%
#347590000000
0!
0%
#347595000000
1!
1%
#347600000000
0!
0%
#347605000000
1!
1%
#347610000000
0!
0%
#347615000000
1!
1%
#347620000000
0!
0%
#347625000000
1!
1%
#347630000000
0!
0%
#347635000000
1!
1%
#347640000000
0!
0%
#347645000000
1!
1%
#347650000000
0!
0%
#347655000000
1!
1%
#347660000000
0!
0%
#347665000000
1!
1%
#347670000000
0!
0%
#347675000000
1!
1%
#347680000000
0!
0%
#347685000000
1!
1%
#347690000000
0!
0%
#347695000000
1!
1%
#347700000000
0!
0%
#347705000000
1!
1%
#347710000000
0!
0%
#347715000000
1!
1%
#347720000000
0!
0%
#347725000000
1!
1%
#347730000000
0!
0%
#347735000000
1!
1%
#347740000000
0!
0%
#347745000000
1!
1%
#347750000000
0!
0%
#347755000000
1!
1%
#347760000000
0!
0%
#347765000000
1!
1%
#347770000000
0!
0%
#347775000000
1!
1%
#347780000000
0!
0%
#347785000000
1!
1%
#347790000000
0!
0%
#347795000000
1!
1%
#347800000000
0!
0%
#347805000000
1!
1%
#347810000000
0!
0%
#347815000000
1!
1%
#347820000000
0!
0%
#347825000000
1!
1%
#347830000000
0!
0%
#347835000000
1!
1%
#347840000000
0!
0%
#347845000000
1!
1%
#347850000000
0!
0%
#347855000000
1!
1%
#347860000000
0!
0%
#347865000000
1!
1%
#347870000000
0!
0%
#347875000000
1!
1%
#347880000000
0!
0%
#347885000000
1!
1%
#347890000000
0!
0%
#347895000000
1!
1%
#347900000000
0!
0%
#347905000000
1!
1%
#347910000000
0!
0%
#347915000000
1!
1%
#347920000000
0!
0%
#347925000000
1!
1%
#347930000000
0!
0%
#347935000000
1!
1%
#347940000000
0!
0%
#347945000000
1!
1%
#347950000000
0!
0%
#347955000000
1!
1%
#347960000000
0!
0%
#347965000000
1!
1%
#347970000000
0!
0%
#347975000000
1!
1%
#347980000000
0!
0%
#347985000000
1!
1%
#347990000000
0!
0%
#347995000000
1!
1%
#348000000000
0!
0%
#348005000000
1!
1%
#348010000000
0!
0%
#348015000000
1!
1%
#348020000000
0!
0%
#348025000000
1!
1%
#348030000000
0!
0%
#348035000000
1!
1%
#348040000000
0!
0%
#348045000000
1!
1%
#348050000000
0!
0%
#348055000000
1!
1%
#348060000000
0!
0%
#348065000000
1!
1%
#348070000000
0!
0%
#348075000000
1!
1%
#348080000000
0!
0%
#348085000000
1!
1%
#348090000000
0!
0%
#348095000000
1!
1%
#348100000000
0!
0%
#348105000000
1!
1%
#348110000000
0!
0%
#348115000000
1!
1%
#348120000000
0!
0%
#348125000000
1!
1%
#348130000000
0!
0%
#348135000000
1!
1%
#348140000000
0!
0%
#348145000000
1!
1%
#348150000000
0!
0%
#348155000000
1!
1%
#348160000000
0!
0%
#348165000000
1!
1%
#348170000000
0!
0%
#348175000000
1!
1%
#348180000000
0!
0%
#348185000000
1!
1%
#348190000000
0!
0%
#348195000000
1!
1%
#348200000000
0!
0%
#348205000000
1!
1%
#348210000000
0!
0%
#348215000000
1!
1%
#348220000000
0!
0%
#348225000000
1!
1%
#348230000000
0!
0%
#348235000000
1!
1%
#348240000000
0!
0%
#348245000000
1!
1%
#348250000000
0!
0%
#348255000000
1!
1%
#348260000000
0!
0%
#348265000000
1!
1%
#348270000000
0!
0%
#348275000000
1!
1%
#348280000000
0!
0%
#348285000000
1!
1%
#348290000000
0!
0%
#348295000000
1!
1%
#348300000000
0!
0%
#348305000000
1!
1%
#348310000000
0!
0%
#348315000000
1!
1%
#348320000000
0!
0%
#348325000000
1!
1%
#348330000000
0!
0%
#348335000000
1!
1%
#348340000000
0!
0%
#348345000000
1!
1%
#348350000000
0!
0%
#348355000000
1!
1%
#348360000000
0!
0%
#348365000000
1!
1%
#348370000000
0!
0%
#348375000000
1!
1%
#348380000000
0!
0%
#348385000000
1!
1%
#348390000000
0!
0%
#348395000000
1!
1%
#348400000000
0!
0%
#348405000000
1!
1%
#348410000000
0!
0%
#348415000000
1!
1%
#348420000000
0!
0%
#348425000000
1!
1%
#348430000000
0!
0%
#348435000000
1!
1%
#348440000000
0!
0%
#348445000000
1!
1%
#348450000000
0!
0%
#348455000000
1!
1%
#348460000000
0!
0%
#348465000000
1!
1%
#348470000000
0!
0%
#348475000000
1!
1%
#348480000000
0!
0%
#348485000000
1!
1%
#348490000000
0!
0%
#348495000000
1!
1%
#348500000000
0!
0%
#348505000000
1!
1%
#348510000000
0!
0%
#348515000000
1!
1%
#348520000000
0!
0%
#348525000000
1!
1%
#348530000000
0!
0%
#348535000000
1!
1%
#348540000000
0!
0%
#348545000000
1!
1%
#348550000000
0!
0%
#348555000000
1!
1%
#348560000000
0!
0%
#348565000000
1!
1%
#348570000000
0!
0%
#348575000000
1!
1%
#348580000000
0!
0%
#348585000000
1!
1%
#348590000000
0!
0%
#348595000000
1!
1%
#348600000000
0!
0%
#348605000000
1!
1%
#348610000000
0!
0%
#348615000000
1!
1%
#348620000000
0!
0%
#348625000000
1!
1%
#348630000000
0!
0%
#348635000000
1!
1%
#348640000000
0!
0%
#348645000000
1!
1%
#348650000000
0!
0%
#348655000000
1!
1%
#348660000000
0!
0%
#348665000000
1!
1%
#348670000000
0!
0%
#348675000000
1!
1%
#348680000000
0!
0%
#348685000000
1!
1%
#348690000000
0!
0%
#348695000000
1!
1%
#348700000000
0!
0%
#348705000000
1!
1%
#348710000000
0!
0%
#348715000000
1!
1%
#348720000000
0!
0%
#348725000000
1!
1%
#348730000000
0!
0%
#348735000000
1!
1%
#348740000000
0!
0%
#348745000000
1!
1%
#348750000000
0!
0%
#348755000000
1!
1%
#348760000000
0!
0%
#348765000000
1!
1%
#348770000000
0!
0%
#348775000000
1!
1%
#348780000000
0!
0%
#348785000000
1!
1%
#348790000000
0!
0%
#348795000000
1!
1%
#348800000000
0!
0%
#348805000000
1!
1%
#348810000000
0!
0%
#348815000000
1!
1%
#348820000000
0!
0%
#348825000000
1!
1%
#348830000000
0!
0%
#348835000000
1!
1%
#348840000000
0!
0%
#348845000000
1!
1%
#348850000000
0!
0%
#348855000000
1!
1%
#348860000000
0!
0%
#348865000000
1!
1%
#348870000000
0!
0%
#348875000000
1!
1%
#348880000000
0!
0%
#348885000000
1!
1%
#348890000000
0!
0%
#348895000000
1!
1%
#348900000000
0!
0%
#348905000000
1!
1%
#348910000000
0!
0%
#348915000000
1!
1%
#348920000000
0!
0%
#348925000000
1!
1%
#348930000000
0!
0%
#348935000000
1!
1%
#348940000000
0!
0%
#348945000000
1!
1%
#348950000000
0!
0%
#348955000000
1!
1%
#348960000000
0!
0%
#348965000000
1!
1%
#348970000000
0!
0%
#348975000000
1!
1%
#348980000000
0!
0%
#348985000000
1!
1%
#348990000000
0!
0%
#348995000000
1!
1%
#349000000000
0!
0%
#349005000000
1!
1%
#349010000000
0!
0%
#349015000000
1!
1%
#349020000000
0!
0%
#349025000000
1!
1%
#349030000000
0!
0%
#349035000000
1!
1%
#349040000000
0!
0%
#349045000000
1!
1%
#349050000000
0!
0%
#349055000000
1!
1%
#349060000000
0!
0%
#349065000000
1!
1%
#349070000000
0!
0%
#349075000000
1!
1%
#349080000000
0!
0%
#349085000000
1!
1%
#349090000000
0!
0%
#349095000000
1!
1%
#349100000000
0!
0%
#349105000000
1!
1%
#349110000000
0!
0%
#349115000000
1!
1%
#349120000000
0!
0%
#349125000000
1!
1%
#349130000000
0!
0%
#349135000000
1!
1%
#349140000000
0!
0%
#349145000000
1!
1%
#349150000000
0!
0%
#349155000000
1!
1%
#349160000000
0!
0%
#349165000000
1!
1%
#349170000000
0!
0%
#349175000000
1!
1%
#349180000000
0!
0%
#349185000000
1!
1%
#349190000000
0!
0%
#349195000000
1!
1%
#349200000000
0!
0%
#349205000000
1!
1%
#349210000000
0!
0%
#349215000000
1!
1%
#349220000000
0!
0%
#349225000000
1!
1%
#349230000000
0!
0%
#349235000000
1!
1%
#349240000000
0!
0%
#349245000000
1!
1%
#349250000000
0!
0%
#349255000000
1!
1%
#349260000000
0!
0%
#349265000000
1!
1%
#349270000000
0!
0%
#349275000000
1!
1%
#349280000000
0!
0%
#349285000000
1!
1%
#349290000000
0!
0%
#349295000000
1!
1%
#349300000000
0!
0%
#349305000000
1!
1%
#349310000000
0!
0%
#349315000000
1!
1%
#349320000000
0!
0%
#349325000000
1!
1%
#349330000000
0!
0%
#349335000000
1!
1%
#349340000000
0!
0%
#349345000000
1!
1%
#349350000000
0!
0%
#349355000000
1!
1%
#349360000000
0!
0%
#349365000000
1!
1%
#349370000000
0!
0%
#349375000000
1!
1%
#349380000000
0!
0%
#349385000000
1!
1%
#349390000000
0!
0%
#349395000000
1!
1%
#349400000000
0!
0%
#349405000000
1!
1%
#349410000000
0!
0%
#349415000000
1!
1%
#349420000000
0!
0%
#349425000000
1!
1%
#349430000000
0!
0%
#349435000000
1!
1%
#349440000000
0!
0%
#349445000000
1!
1%
#349450000000
0!
0%
#349455000000
1!
1%
#349460000000
0!
0%
#349465000000
1!
1%
#349470000000
0!
0%
#349475000000
1!
1%
#349480000000
0!
0%
#349485000000
1!
1%
#349490000000
0!
0%
#349495000000
1!
1%
#349500000000
0!
0%
#349505000000
1!
1%
#349510000000
0!
0%
#349515000000
1!
1%
#349520000000
0!
0%
#349525000000
1!
1%
#349530000000
0!
0%
#349535000000
1!
1%
#349540000000
0!
0%
#349545000000
1!
1%
#349550000000
0!
0%
#349555000000
1!
1%
#349560000000
0!
0%
#349565000000
1!
1%
#349570000000
0!
0%
#349575000000
1!
1%
#349580000000
0!
0%
#349585000000
1!
1%
#349590000000
0!
0%
#349595000000
1!
1%
#349600000000
0!
0%
#349605000000
1!
1%
#349610000000
0!
0%
#349615000000
1!
1%
#349620000000
0!
0%
#349625000000
1!
1%
#349630000000
0!
0%
#349635000000
1!
1%
#349640000000
0!
0%
#349645000000
1!
1%
#349650000000
0!
0%
#349655000000
1!
1%
#349660000000
0!
0%
#349665000000
1!
1%
#349670000000
0!
0%
#349675000000
1!
1%
#349680000000
0!
0%
#349685000000
1!
1%
#349690000000
0!
0%
#349695000000
1!
1%
#349700000000
0!
0%
#349705000000
1!
1%
#349710000000
0!
0%
#349715000000
1!
1%
#349720000000
0!
0%
#349725000000
1!
1%
#349730000000
0!
0%
#349735000000
1!
1%
#349740000000
0!
0%
#349745000000
1!
1%
#349750000000
0!
0%
#349755000000
1!
1%
#349760000000
0!
0%
#349765000000
1!
1%
#349770000000
0!
0%
#349775000000
1!
1%
#349780000000
0!
0%
#349785000000
1!
1%
#349790000000
0!
0%
#349795000000
1!
1%
#349800000000
0!
0%
#349805000000
1!
1%
#349810000000
0!
0%
#349815000000
1!
1%
#349820000000
0!
0%
#349825000000
1!
1%
#349830000000
0!
0%
#349835000000
1!
1%
#349840000000
0!
0%
#349845000000
1!
1%
#349850000000
0!
0%
#349855000000
1!
1%
#349860000000
0!
0%
#349865000000
1!
1%
#349870000000
0!
0%
#349875000000
1!
1%
#349880000000
0!
0%
#349885000000
1!
1%
#349890000000
0!
0%
#349895000000
1!
1%
#349900000000
0!
0%
#349905000000
1!
1%
#349910000000
0!
0%
#349915000000
1!
1%
#349920000000
0!
0%
#349925000000
1!
1%
#349930000000
0!
0%
#349935000000
1!
1%
#349940000000
0!
0%
#349945000000
1!
1%
#349950000000
0!
0%
#349955000000
1!
1%
#349960000000
0!
0%
#349965000000
1!
1%
#349970000000
0!
0%
#349975000000
1!
1%
#349980000000
0!
0%
#349985000000
1!
1%
#349990000000
0!
0%
#349995000000
1!
1%
#350000000000
0!
0%
#350005000000
1!
1%
#350010000000
0!
0%
#350015000000
1!
1%
#350020000000
0!
0%
#350025000000
1!
1%
#350030000000
0!
0%
#350035000000
1!
1%
#350040000000
0!
0%
#350045000000
1!
1%
#350050000000
0!
0%
#350055000000
1!
1%
#350060000000
0!
0%
#350065000000
1!
1%
#350070000000
0!
0%
#350075000000
1!
1%
#350080000000
0!
0%
#350085000000
1!
1%
#350090000000
0!
0%
#350095000000
1!
1%
#350100000000
0!
0%
#350105000000
1!
1%
#350110000000
0!
0%
#350115000000
1!
1%
#350120000000
0!
0%
#350125000000
1!
1%
#350130000000
0!
0%
#350135000000
1!
1%
#350140000000
0!
0%
#350145000000
1!
1%
#350150000000
0!
0%
#350155000000
1!
1%
#350160000000
0!
0%
#350165000000
1!
1%
#350170000000
0!
0%
#350175000000
1!
1%
#350180000000
0!
0%
#350185000000
1!
1%
#350190000000
0!
0%
#350195000000
1!
1%
#350200000000
0!
0%
#350205000000
1!
1%
#350210000000
0!
0%
#350215000000
1!
1%
#350220000000
0!
0%
#350225000000
1!
1%
#350230000000
0!
0%
#350235000000
1!
1%
#350240000000
0!
0%
#350245000000
1!
1%
#350250000000
0!
0%
#350255000000
1!
1%
#350260000000
0!
0%
#350265000000
1!
1%
#350270000000
0!
0%
#350275000000
1!
1%
#350280000000
0!
0%
#350285000000
1!
1%
#350290000000
0!
0%
#350295000000
1!
1%
#350300000000
0!
0%
#350305000000
1!
1%
#350310000000
0!
0%
#350315000000
1!
1%
#350320000000
0!
0%
#350325000000
1!
1%
#350330000000
0!
0%
#350335000000
1!
1%
#350340000000
0!
0%
#350345000000
1!
1%
#350350000000
0!
0%
#350355000000
1!
1%
#350360000000
0!
0%
#350365000000
1!
1%
#350370000000
0!
0%
#350375000000
1!
1%
#350380000000
0!
0%
#350385000000
1!
1%
#350390000000
0!
0%
#350395000000
1!
1%
#350400000000
0!
0%
#350405000000
1!
1%
#350410000000
0!
0%
#350415000000
1!
1%
#350420000000
0!
0%
#350425000000
1!
1%
#350430000000
0!
0%
#350435000000
1!
1%
#350440000000
0!
0%
#350445000000
1!
1%
#350450000000
0!
0%
#350455000000
1!
1%
#350460000000
0!
0%
#350465000000
1!
1%
#350470000000
0!
0%
#350475000000
1!
1%
#350480000000
0!
0%
#350485000000
1!
1%
#350490000000
0!
0%
#350495000000
1!
1%
#350500000000
0!
0%
#350505000000
1!
1%
#350510000000
0!
0%
#350515000000
1!
1%
#350520000000
0!
0%
#350525000000
1!
1%
#350530000000
0!
0%
#350535000000
1!
1%
#350540000000
0!
0%
#350545000000
1!
1%
#350550000000
0!
0%
#350555000000
1!
1%
#350560000000
0!
0%
#350565000000
1!
1%
#350570000000
0!
0%
#350575000000
1!
1%
#350580000000
0!
0%
#350585000000
1!
1%
#350590000000
0!
0%
#350595000000
1!
1%
#350600000000
0!
0%
#350605000000
1!
1%
#350610000000
0!
0%
#350615000000
1!
1%
#350620000000
0!
0%
#350625000000
1!
1%
#350630000000
0!
0%
#350635000000
1!
1%
#350640000000
0!
0%
#350645000000
1!
1%
#350650000000
0!
0%
#350655000000
1!
1%
#350660000000
0!
0%
#350665000000
1!
1%
#350670000000
0!
0%
#350675000000
1!
1%
#350680000000
0!
0%
#350685000000
1!
1%
#350690000000
0!
0%
#350695000000
1!
1%
#350700000000
0!
0%
#350705000000
1!
1%
#350710000000
0!
0%
#350715000000
1!
1%
#350720000000
0!
0%
#350725000000
1!
1%
#350730000000
0!
0%
#350735000000
1!
1%
#350740000000
0!
0%
#350745000000
1!
1%
#350750000000
0!
0%
#350755000000
1!
1%
#350760000000
0!
0%
#350765000000
1!
1%
#350770000000
0!
0%
#350775000000
1!
1%
#350780000000
0!
0%
#350785000000
1!
1%
#350790000000
0!
0%
#350795000000
1!
1%
#350800000000
0!
0%
#350805000000
1!
1%
#350810000000
0!
0%
#350815000000
1!
1%
#350820000000
0!
0%
#350825000000
1!
1%
#350830000000
0!
0%
#350835000000
1!
1%
#350840000000
0!
0%
#350845000000
1!
1%
#350850000000
0!
0%
#350855000000
1!
1%
#350860000000
0!
0%
#350865000000
1!
1%
#350870000000
0!
0%
#350875000000
1!
1%
#350880000000
0!
0%
#350885000000
1!
1%
#350890000000
0!
0%
#350895000000
1!
1%
#350900000000
0!
0%
#350905000000
1!
1%
#350910000000
0!
0%
#350915000000
1!
1%
#350920000000
0!
0%
#350925000000
1!
1%
#350930000000
0!
0%
#350935000000
1!
1%
#350940000000
0!
0%
#350945000000
1!
1%
#350950000000
0!
0%
#350955000000
1!
1%
#350960000000
0!
0%
#350965000000
1!
1%
#350970000000
0!
0%
#350975000000
1!
1%
#350980000000
0!
0%
#350985000000
1!
1%
#350990000000
0!
0%
#350995000000
1!
1%
#351000000000
0!
0%
#351005000000
1!
1%
#351010000000
0!
0%
#351015000000
1!
1%
#351020000000
0!
0%
#351025000000
1!
1%
#351030000000
0!
0%
#351035000000
1!
1%
#351040000000
0!
0%
#351045000000
1!
1%
#351050000000
0!
0%
#351055000000
1!
1%
#351060000000
0!
0%
#351065000000
1!
1%
#351070000000
0!
0%
#351075000000
1!
1%
#351080000000
0!
0%
#351085000000
1!
1%
#351090000000
0!
0%
#351095000000
1!
1%
#351100000000
0!
0%
#351105000000
1!
1%
#351110000000
0!
0%
#351115000000
1!
1%
#351120000000
0!
0%
#351125000000
1!
1%
#351130000000
0!
0%
#351135000000
1!
1%
#351140000000
0!
0%
#351145000000
1!
1%
#351150000000
0!
0%
#351155000000
1!
1%
#351160000000
0!
0%
#351165000000
1!
1%
#351170000000
0!
0%
#351175000000
1!
1%
#351180000000
0!
0%
#351185000000
1!
1%
#351190000000
0!
0%
#351195000000
1!
1%
#351200000000
0!
0%
#351205000000
1!
1%
#351210000000
0!
0%
#351215000000
1!
1%
#351220000000
0!
0%
#351225000000
1!
1%
#351230000000
0!
0%
#351235000000
1!
1%
#351240000000
0!
0%
#351245000000
1!
1%
#351250000000
0!
0%
#351255000000
1!
1%
#351260000000
0!
0%
#351265000000
1!
1%
#351270000000
0!
0%
#351275000000
1!
1%
#351280000000
0!
0%
#351285000000
1!
1%
#351290000000
0!
0%
#351295000000
1!
1%
#351300000000
0!
0%
#351305000000
1!
1%
#351310000000
0!
0%
#351315000000
1!
1%
#351320000000
0!
0%
#351325000000
1!
1%
#351330000000
0!
0%
#351335000000
1!
1%
#351340000000
0!
0%
#351345000000
1!
1%
#351350000000
0!
0%
#351355000000
1!
1%
#351360000000
0!
0%
#351365000000
1!
1%
#351370000000
0!
0%
#351375000000
1!
1%
#351380000000
0!
0%
#351385000000
1!
1%
#351390000000
0!
0%
#351395000000
1!
1%
#351400000000
0!
0%
#351405000000
1!
1%
#351410000000
0!
0%
#351415000000
1!
1%
#351420000000
0!
0%
#351425000000
1!
1%
#351430000000
0!
0%
#351435000000
1!
1%
#351440000000
0!
0%
#351445000000
1!
1%
#351450000000
0!
0%
#351455000000
1!
1%
#351460000000
0!
0%
#351465000000
1!
1%
#351470000000
0!
0%
#351475000000
1!
1%
#351480000000
0!
0%
#351485000000
1!
1%
#351490000000
0!
0%
#351495000000
1!
1%
#351500000000
0!
0%
#351505000000
1!
1%
#351510000000
0!
0%
#351515000000
1!
1%
#351520000000
0!
0%
#351525000000
1!
1%
#351530000000
0!
0%
#351535000000
1!
1%
#351540000000
0!
0%
#351545000000
1!
1%
#351550000000
0!
0%
#351555000000
1!
1%
#351560000000
0!
0%
#351565000000
1!
1%
#351570000000
0!
0%
#351575000000
1!
1%
#351580000000
0!
0%
#351585000000
1!
1%
#351590000000
0!
0%
#351595000000
1!
1%
#351600000000
0!
0%
#351605000000
1!
1%
#351610000000
0!
0%
#351615000000
1!
1%
#351620000000
0!
0%
#351625000000
1!
1%
#351630000000
0!
0%
#351635000000
1!
1%
#351640000000
0!
0%
#351645000000
1!
1%
#351650000000
0!
0%
#351655000000
1!
1%
#351660000000
0!
0%
#351665000000
1!
1%
#351670000000
0!
0%
#351675000000
1!
1%
#351680000000
0!
0%
#351685000000
1!
1%
#351690000000
0!
0%
#351695000000
1!
1%
#351700000000
0!
0%
#351705000000
1!
1%
#351710000000
0!
0%
#351715000000
1!
1%
#351720000000
0!
0%
#351725000000
1!
1%
#351730000000
0!
0%
#351735000000
1!
1%
#351740000000
0!
0%
#351745000000
1!
1%
#351750000000
0!
0%
#351755000000
1!
1%
#351760000000
0!
0%
#351765000000
1!
1%
#351770000000
0!
0%
#351775000000
1!
1%
#351780000000
0!
0%
#351785000000
1!
1%
#351790000000
0!
0%
#351795000000
1!
1%
#351800000000
0!
0%
#351805000000
1!
1%
#351810000000
0!
0%
#351815000000
1!
1%
#351820000000
0!
0%
#351825000000
1!
1%
#351830000000
0!
0%
#351835000000
1!
1%
#351840000000
0!
0%
#351845000000
1!
1%
#351850000000
0!
0%
#351855000000
1!
1%
#351860000000
0!
0%
#351865000000
1!
1%
#351870000000
0!
0%
#351875000000
1!
1%
#351880000000
0!
0%
#351885000000
1!
1%
#351890000000
0!
0%
#351895000000
1!
1%
#351900000000
0!
0%
#351905000000
1!
1%
#351910000000
0!
0%
#351915000000
1!
1%
#351920000000
0!
0%
#351925000000
1!
1%
#351930000000
0!
0%
#351935000000
1!
1%
#351940000000
0!
0%
#351945000000
1!
1%
#351950000000
0!
0%
#351955000000
1!
1%
#351960000000
0!
0%
#351965000000
1!
1%
#351970000000
0!
0%
#351975000000
1!
1%
#351980000000
0!
0%
#351985000000
1!
1%
#351990000000
0!
0%
#351995000000
1!
1%
#352000000000
0!
0%
#352005000000
1!
1%
#352010000000
0!
0%
#352015000000
1!
1%
#352020000000
0!
0%
#352025000000
1!
1%
#352030000000
0!
0%
#352035000000
1!
1%
#352040000000
0!
0%
#352045000000
1!
1%
#352050000000
0!
0%
#352055000000
1!
1%
#352060000000
0!
0%
#352065000000
1!
1%
#352070000000
0!
0%
#352075000000
1!
1%
#352080000000
0!
0%
#352085000000
1!
1%
#352090000000
0!
0%
#352095000000
1!
1%
#352100000000
0!
0%
#352105000000
1!
1%
#352110000000
0!
0%
#352115000000
1!
1%
#352120000000
0!
0%
#352125000000
1!
1%
#352130000000
0!
0%
#352135000000
1!
1%
#352140000000
0!
0%
#352145000000
1!
1%
#352150000000
0!
0%
#352155000000
1!
1%
#352160000000
0!
0%
#352165000000
1!
1%
#352170000000
0!
0%
#352175000000
1!
1%
#352180000000
0!
0%
#352185000000
1!
1%
#352190000000
0!
0%
#352195000000
1!
1%
#352200000000
0!
0%
#352205000000
1!
1%
#352210000000
0!
0%
#352215000000
1!
1%
#352220000000
0!
0%
#352225000000
1!
1%
#352230000000
0!
0%
#352235000000
1!
1%
#352240000000
0!
0%
#352245000000
1!
1%
#352250000000
0!
0%
#352255000000
1!
1%
#352260000000
0!
0%
#352265000000
1!
1%
#352270000000
0!
0%
#352275000000
1!
1%
#352280000000
0!
0%
#352285000000
1!
1%
#352290000000
0!
0%
#352295000000
1!
1%
#352300000000
0!
0%
#352305000000
1!
1%
#352310000000
0!
0%
#352315000000
1!
1%
#352320000000
0!
0%
#352325000000
1!
1%
#352330000000
0!
0%
#352335000000
1!
1%
#352340000000
0!
0%
#352345000000
1!
1%
#352350000000
0!
0%
#352355000000
1!
1%
#352360000000
0!
0%
#352365000000
1!
1%
#352370000000
0!
0%
#352375000000
1!
1%
#352380000000
0!
0%
#352385000000
1!
1%
#352390000000
0!
0%
#352395000000
1!
1%
#352400000000
0!
0%
#352405000000
1!
1%
#352410000000
0!
0%
#352415000000
1!
1%
#352420000000
0!
0%
#352425000000
1!
1%
#352430000000
0!
0%
#352435000000
1!
1%
#352440000000
0!
0%
#352445000000
1!
1%
#352450000000
0!
0%
#352455000000
1!
1%
#352460000000
0!
0%
#352465000000
1!
1%
#352470000000
0!
0%
#352475000000
1!
1%
#352480000000
0!
0%
#352485000000
1!
1%
#352490000000
0!
0%
#352495000000
1!
1%
#352500000000
0!
0%
#352505000000
1!
1%
#352510000000
0!
0%
#352515000000
1!
1%
#352520000000
0!
0%
#352525000000
1!
1%
#352530000000
0!
0%
#352535000000
1!
1%
#352540000000
0!
0%
#352545000000
1!
1%
#352550000000
0!
0%
#352555000000
1!
1%
#352560000000
0!
0%
#352565000000
1!
1%
#352570000000
0!
0%
#352575000000
1!
1%
#352580000000
0!
0%
#352585000000
1!
1%
#352590000000
0!
0%
#352595000000
1!
1%
#352600000000
0!
0%
#352605000000
1!
1%
#352610000000
0!
0%
#352615000000
1!
1%
#352620000000
0!
0%
#352625000000
1!
1%
#352630000000
0!
0%
#352635000000
1!
1%
#352640000000
0!
0%
#352645000000
1!
1%
#352650000000
0!
0%
#352655000000
1!
1%
#352660000000
0!
0%
#352665000000
1!
1%
#352670000000
0!
0%
#352675000000
1!
1%
#352680000000
0!
0%
#352685000000
1!
1%
#352690000000
0!
0%
#352695000000
1!
1%
#352700000000
0!
0%
#352705000000
1!
1%
#352710000000
0!
0%
#352715000000
1!
1%
#352720000000
0!
0%
#352725000000
1!
1%
#352730000000
0!
0%
#352735000000
1!
1%
#352740000000
0!
0%
#352745000000
1!
1%
#352750000000
0!
0%
#352755000000
1!
1%
#352760000000
0!
0%
#352765000000
1!
1%
#352770000000
0!
0%
#352775000000
1!
1%
#352780000000
0!
0%
#352785000000
1!
1%
#352790000000
0!
0%
#352795000000
1!
1%
#352800000000
0!
0%
#352805000000
1!
1%
#352810000000
0!
0%
#352815000000
1!
1%
#352820000000
0!
0%
#352825000000
1!
1%
#352830000000
0!
0%
#352835000000
1!
1%
#352840000000
0!
0%
#352845000000
1!
1%
#352850000000
0!
0%
#352855000000
1!
1%
#352860000000
0!
0%
#352865000000
1!
1%
#352870000000
0!
0%
#352875000000
1!
1%
#352880000000
0!
0%
#352885000000
1!
1%
#352890000000
0!
0%
#352895000000
1!
1%
#352900000000
0!
0%
#352905000000
1!
1%
#352910000000
0!
0%
#352915000000
1!
1%
#352920000000
0!
0%
#352925000000
1!
1%
#352930000000
0!
0%
#352935000000
1!
1%
#352940000000
0!
0%
#352945000000
1!
1%
#352950000000
0!
0%
#352955000000
1!
1%
#352960000000
0!
0%
#352965000000
1!
1%
#352970000000
0!
0%
#352975000000
1!
1%
#352980000000
0!
0%
#352985000000
1!
1%
#352990000000
0!
0%
#352995000000
1!
1%
#353000000000
0!
0%
#353005000000
1!
1%
#353010000000
0!
0%
#353015000000
1!
1%
#353020000000
0!
0%
#353025000000
1!
1%
#353030000000
0!
0%
#353035000000
1!
1%
#353040000000
0!
0%
#353045000000
1!
1%
#353050000000
0!
0%
#353055000000
1!
1%
#353060000000
0!
0%
#353065000000
1!
1%
#353070000000
0!
0%
#353075000000
1!
1%
#353080000000
0!
0%
#353085000000
1!
1%
#353090000000
0!
0%
#353095000000
1!
1%
#353100000000
0!
0%
#353105000000
1!
1%
#353110000000
0!
0%
#353115000000
1!
1%
#353120000000
0!
0%
#353125000000
1!
1%
#353130000000
0!
0%
#353135000000
1!
1%
#353140000000
0!
0%
#353145000000
1!
1%
#353150000000
0!
0%
#353155000000
1!
1%
#353160000000
0!
0%
#353165000000
1!
1%
#353170000000
0!
0%
#353175000000
1!
1%
#353180000000
0!
0%
#353185000000
1!
1%
#353190000000
0!
0%
#353195000000
1!
1%
#353200000000
0!
0%
#353205000000
1!
1%
#353210000000
0!
0%
#353215000000
1!
1%
#353220000000
0!
0%
#353225000000
1!
1%
#353230000000
0!
0%
#353235000000
1!
1%
#353240000000
0!
0%
#353245000000
1!
1%
#353250000000
0!
0%
#353255000000
1!
1%
#353260000000
0!
0%
#353265000000
1!
1%
#353270000000
0!
0%
#353275000000
1!
1%
#353280000000
0!
0%
#353285000000
1!
1%
#353290000000
0!
0%
#353295000000
1!
1%
#353300000000
0!
0%
#353305000000
1!
1%
#353310000000
0!
0%
#353315000000
1!
1%
#353320000000
0!
0%
#353325000000
1!
1%
#353330000000
0!
0%
#353335000000
1!
1%
#353340000000
0!
0%
#353345000000
1!
1%
#353350000000
0!
0%
#353355000000
1!
1%
#353360000000
0!
0%
#353365000000
1!
1%
#353370000000
0!
0%
#353375000000
1!
1%
#353380000000
0!
0%
#353385000000
1!
1%
#353390000000
0!
0%
#353395000000
1!
1%
#353400000000
0!
0%
#353405000000
1!
1%
#353410000000
0!
0%
#353415000000
1!
1%
#353420000000
0!
0%
#353425000000
1!
1%
#353430000000
0!
0%
#353435000000
1!
1%
#353440000000
0!
0%
#353445000000
1!
1%
#353450000000
0!
0%
#353455000000
1!
1%
#353460000000
0!
0%
#353465000000
1!
1%
#353470000000
0!
0%
#353475000000
1!
1%
#353480000000
0!
0%
#353485000000
1!
1%
#353490000000
0!
0%
#353495000000
1!
1%
#353500000000
0!
0%
#353505000000
1!
1%
#353510000000
0!
0%
#353515000000
1!
1%
#353520000000
0!
0%
#353525000000
1!
1%
#353530000000
0!
0%
#353535000000
1!
1%
#353540000000
0!
0%
#353545000000
1!
1%
#353550000000
0!
0%
#353555000000
1!
1%
#353560000000
0!
0%
#353565000000
1!
1%
#353570000000
0!
0%
#353575000000
1!
1%
#353580000000
0!
0%
#353585000000
1!
1%
#353590000000
0!
0%
#353595000000
1!
1%
#353600000000
0!
0%
#353605000000
1!
1%
#353610000000
0!
0%
#353615000000
1!
1%
#353620000000
0!
0%
#353625000000
1!
1%
#353630000000
0!
0%
#353635000000
1!
1%
#353640000000
0!
0%
#353645000000
1!
1%
#353650000000
0!
0%
#353655000000
1!
1%
#353660000000
0!
0%
#353665000000
1!
1%
#353670000000
0!
0%
#353675000000
1!
1%
#353680000000
0!
0%
#353685000000
1!
1%
#353690000000
0!
0%
#353695000000
1!
1%
#353700000000
0!
0%
#353705000000
1!
1%
#353710000000
0!
0%
#353715000000
1!
1%
#353720000000
0!
0%
#353725000000
1!
1%
#353730000000
0!
0%
#353735000000
1!
1%
#353740000000
0!
0%
#353745000000
1!
1%
#353750000000
0!
0%
#353755000000
1!
1%
#353760000000
0!
0%
#353765000000
1!
1%
#353770000000
0!
0%
#353775000000
1!
1%
#353780000000
0!
0%
#353785000000
1!
1%
#353790000000
0!
0%
#353795000000
1!
1%
#353800000000
0!
0%
#353805000000
1!
1%
#353810000000
0!
0%
#353815000000
1!
1%
#353820000000
0!
0%
#353825000000
1!
1%
#353830000000
0!
0%
#353835000000
1!
1%
#353840000000
0!
0%
#353845000000
1!
1%
#353850000000
0!
0%
#353855000000
1!
1%
#353860000000
0!
0%
#353865000000
1!
1%
#353870000000
0!
0%
#353875000000
1!
1%
#353880000000
0!
0%
#353885000000
1!
1%
#353890000000
0!
0%
#353895000000
1!
1%
#353900000000
0!
0%
#353905000000
1!
1%
#353910000000
0!
0%
#353915000000
1!
1%
#353920000000
0!
0%
#353925000000
1!
1%
#353930000000
0!
0%
#353935000000
1!
1%
#353940000000
0!
0%
#353945000000
1!
1%
#353950000000
0!
0%
#353955000000
1!
1%
#353960000000
0!
0%
#353965000000
1!
1%
#353970000000
0!
0%
#353975000000
1!
1%
#353980000000
0!
0%
#353985000000
1!
1%
#353990000000
0!
0%
#353995000000
1!
1%
#354000000000
0!
0%
#354005000000
1!
1%
#354010000000
0!
0%
#354015000000
1!
1%
#354020000000
0!
0%
#354025000000
1!
1%
#354030000000
0!
0%
#354035000000
1!
1%
#354040000000
0!
0%
#354045000000
1!
1%
#354050000000
0!
0%
#354055000000
1!
1%
#354060000000
0!
0%
#354065000000
1!
1%
#354070000000
0!
0%
#354075000000
1!
1%
#354080000000
0!
0%
#354085000000
1!
1%
#354090000000
0!
0%
#354095000000
1!
1%
#354100000000
0!
0%
#354105000000
1!
1%
#354110000000
0!
0%
#354115000000
1!
1%
#354120000000
0!
0%
#354125000000
1!
1%
#354130000000
0!
0%
#354135000000
1!
1%
#354140000000
0!
0%
#354145000000
1!
1%
#354150000000
0!
0%
#354155000000
1!
1%
#354160000000
0!
0%
#354165000000
1!
1%
#354170000000
0!
0%
#354175000000
1!
1%
#354180000000
0!
0%
#354185000000
1!
1%
#354190000000
0!
0%
#354195000000
1!
1%
#354200000000
0!
0%
#354205000000
1!
1%
#354210000000
0!
0%
#354215000000
1!
1%
#354220000000
0!
0%
#354225000000
1!
1%
#354230000000
0!
0%
#354235000000
1!
1%
#354240000000
0!
0%
#354245000000
1!
1%
#354250000000
0!
0%
#354255000000
1!
1%
#354260000000
0!
0%
#354265000000
1!
1%
#354270000000
0!
0%
#354275000000
1!
1%
#354280000000
0!
0%
#354285000000
1!
1%
#354290000000
0!
0%
#354295000000
1!
1%
#354300000000
0!
0%
#354305000000
1!
1%
#354310000000
0!
0%
#354315000000
1!
1%
#354320000000
0!
0%
#354325000000
1!
1%
#354330000000
0!
0%
#354335000000
1!
1%
#354340000000
0!
0%
#354345000000
1!
1%
#354350000000
0!
0%
#354355000000
1!
1%
#354360000000
0!
0%
#354365000000
1!
1%
#354370000000
0!
0%
#354375000000
1!
1%
#354380000000
0!
0%
#354385000000
1!
1%
#354390000000
0!
0%
#354395000000
1!
1%
#354400000000
0!
0%
#354405000000
1!
1%
#354410000000
0!
0%
#354415000000
1!
1%
#354420000000
0!
0%
#354425000000
1!
1%
#354430000000
0!
0%
#354435000000
1!
1%
#354440000000
0!
0%
#354445000000
1!
1%
#354450000000
0!
0%
#354455000000
1!
1%
#354460000000
0!
0%
#354465000000
1!
1%
#354470000000
0!
0%
#354475000000
1!
1%
#354480000000
0!
0%
#354485000000
1!
1%
#354490000000
0!
0%
#354495000000
1!
1%
#354500000000
0!
0%
#354505000000
1!
1%
#354510000000
0!
0%
#354515000000
1!
1%
#354520000000
0!
0%
#354525000000
1!
1%
#354530000000
0!
0%
#354535000000
1!
1%
#354540000000
0!
0%
#354545000000
1!
1%
#354550000000
0!
0%
#354555000000
1!
1%
#354560000000
0!
0%
#354565000000
1!
1%
#354570000000
0!
0%
#354575000000
1!
1%
#354580000000
0!
0%
#354585000000
1!
1%
#354590000000
0!
0%
#354595000000
1!
1%
#354600000000
0!
0%
#354605000000
1!
1%
#354610000000
0!
0%
#354615000000
1!
1%
#354620000000
0!
0%
#354625000000
1!
1%
#354630000000
0!
0%
#354635000000
1!
1%
#354640000000
0!
0%
#354645000000
1!
1%
#354650000000
0!
0%
#354655000000
1!
1%
#354660000000
0!
0%
#354665000000
1!
1%
#354670000000
0!
0%
#354675000000
1!
1%
#354680000000
0!
0%
#354685000000
1!
1%
#354690000000
0!
0%
#354695000000
1!
1%
#354700000000
0!
0%
#354705000000
1!
1%
#354710000000
0!
0%
#354715000000
1!
1%
#354720000000
0!
0%
#354725000000
1!
1%
#354730000000
0!
0%
#354735000000
1!
1%
#354740000000
0!
0%
#354745000000
1!
1%
#354750000000
0!
0%
#354755000000
1!
1%
#354760000000
0!
0%
#354765000000
1!
1%
#354770000000
0!
0%
#354775000000
1!
1%
#354780000000
0!
0%
#354785000000
1!
1%
#354790000000
0!
0%
#354795000000
1!
1%
#354800000000
0!
0%
#354805000000
1!
1%
#354810000000
0!
0%
#354815000000
1!
1%
#354820000000
0!
0%
#354825000000
1!
1%
#354830000000
0!
0%
#354835000000
1!
1%
#354840000000
0!
0%
#354845000000
1!
1%
#354850000000
0!
0%
#354855000000
1!
1%
#354860000000
0!
0%
#354865000000
1!
1%
#354870000000
0!
0%
#354875000000
1!
1%
#354880000000
0!
0%
#354885000000
1!
1%
#354890000000
0!
0%
#354895000000
1!
1%
#354900000000
0!
0%
#354905000000
1!
1%
#354910000000
0!
0%
#354915000000
1!
1%
#354920000000
0!
0%
#354925000000
1!
1%
#354930000000
0!
0%
#354935000000
1!
1%
#354940000000
0!
0%
#354945000000
1!
1%
#354950000000
0!
0%
#354955000000
1!
1%
#354960000000
0!
0%
#354965000000
1!
1%
#354970000000
0!
0%
#354975000000
1!
1%
#354980000000
0!
0%
#354985000000
1!
1%
#354990000000
0!
0%
#354995000000
1!
1%
#355000000000
0!
0%
#355005000000
1!
1%
#355010000000
0!
0%
#355015000000
1!
1%
#355020000000
0!
0%
#355025000000
1!
1%
#355030000000
0!
0%
#355035000000
1!
1%
#355040000000
0!
0%
#355045000000
1!
1%
#355050000000
0!
0%
#355055000000
1!
1%
#355060000000
0!
0%
#355065000000
1!
1%
#355070000000
0!
0%
#355075000000
1!
1%
#355080000000
0!
0%
#355085000000
1!
1%
#355090000000
0!
0%
#355095000000
1!
1%
#355100000000
0!
0%
#355105000000
1!
1%
#355110000000
0!
0%
#355115000000
1!
1%
#355120000000
0!
0%
#355125000000
1!
1%
#355130000000
0!
0%
#355135000000
1!
1%
#355140000000
0!
0%
#355145000000
1!
1%
#355150000000
0!
0%
#355155000000
1!
1%
#355160000000
0!
0%
#355165000000
1!
1%
#355170000000
0!
0%
#355175000000
1!
1%
#355180000000
0!
0%
#355185000000
1!
1%
#355190000000
0!
0%
#355195000000
1!
1%
#355200000000
0!
0%
#355205000000
1!
1%
#355210000000
0!
0%
#355215000000
1!
1%
#355220000000
0!
0%
#355225000000
1!
1%
#355230000000
0!
0%
#355235000000
1!
1%
#355240000000
0!
0%
#355245000000
1!
1%
#355250000000
0!
0%
#355255000000
1!
1%
#355260000000
0!
0%
#355265000000
1!
1%
#355270000000
0!
0%
#355275000000
1!
1%
#355280000000
0!
0%
#355285000000
1!
1%
#355290000000
0!
0%
#355295000000
1!
1%
#355300000000
0!
0%
#355305000000
1!
1%
#355310000000
0!
0%
#355315000000
1!
1%
#355320000000
0!
0%
#355325000000
1!
1%
#355330000000
0!
0%
#355335000000
1!
1%
#355340000000
0!
0%
#355345000000
1!
1%
#355350000000
0!
0%
#355355000000
1!
1%
#355360000000
0!
0%
#355365000000
1!
1%
#355370000000
0!
0%
#355375000000
1!
1%
#355380000000
0!
0%
#355385000000
1!
1%
#355390000000
0!
0%
#355395000000
1!
1%
#355400000000
0!
0%
#355405000000
1!
1%
#355410000000
0!
0%
#355415000000
1!
1%
#355420000000
0!
0%
#355425000000
1!
1%
#355430000000
0!
0%
#355435000000
1!
1%
#355440000000
0!
0%
#355445000000
1!
1%
#355450000000
0!
0%
#355455000000
1!
1%
#355460000000
0!
0%
#355465000000
1!
1%
#355470000000
0!
0%
#355475000000
1!
1%
#355480000000
0!
0%
#355485000000
1!
1%
#355490000000
0!
0%
#355495000000
1!
1%
#355500000000
0!
0%
#355505000000
1!
1%
#355510000000
0!
0%
#355515000000
1!
1%
#355520000000
0!
0%
#355525000000
1!
1%
#355530000000
0!
0%
#355535000000
1!
1%
#355540000000
0!
0%
#355545000000
1!
1%
#355550000000
0!
0%
#355555000000
1!
1%
#355560000000
0!
0%
#355565000000
1!
1%
#355570000000
0!
0%
#355575000000
1!
1%
#355580000000
0!
0%
#355585000000
1!
1%
#355590000000
0!
0%
#355595000000
1!
1%
#355600000000
0!
0%
#355605000000
1!
1%
#355610000000
0!
0%
#355615000000
1!
1%
#355620000000
0!
0%
#355625000000
1!
1%
#355630000000
0!
0%
#355635000000
1!
1%
#355640000000
0!
0%
#355645000000
1!
1%
#355650000000
0!
0%
#355655000000
1!
1%
#355660000000
0!
0%
#355665000000
1!
1%
#355670000000
0!
0%
#355675000000
1!
1%
#355680000000
0!
0%
#355685000000
1!
1%
#355690000000
0!
0%
#355695000000
1!
1%
#355700000000
0!
0%
#355705000000
1!
1%
#355710000000
0!
0%
#355715000000
1!
1%
#355720000000
0!
0%
#355725000000
1!
1%
#355730000000
0!
0%
#355735000000
1!
1%
#355740000000
0!
0%
#355745000000
1!
1%
#355750000000
0!
0%
#355755000000
1!
1%
#355760000000
0!
0%
#355765000000
1!
1%
#355770000000
0!
0%
#355775000000
1!
1%
#355780000000
0!
0%
#355785000000
1!
1%
#355790000000
0!
0%
#355795000000
1!
1%
#355800000000
0!
0%
#355805000000
1!
1%
#355810000000
0!
0%
#355815000000
1!
1%
#355820000000
0!
0%
#355825000000
1!
1%
#355830000000
0!
0%
#355835000000
1!
1%
#355840000000
0!
0%
#355845000000
1!
1%
#355850000000
0!
0%
#355855000000
1!
1%
#355860000000
0!
0%
#355865000000
1!
1%
#355870000000
0!
0%
#355875000000
1!
1%
#355880000000
0!
0%
#355885000000
1!
1%
#355890000000
0!
0%
#355895000000
1!
1%
#355900000000
0!
0%
#355905000000
1!
1%
#355910000000
0!
0%
#355915000000
1!
1%
#355920000000
0!
0%
#355925000000
1!
1%
#355930000000
0!
0%
#355935000000
1!
1%
#355940000000
0!
0%
#355945000000
1!
1%
#355950000000
0!
0%
#355955000000
1!
1%
#355960000000
0!
0%
#355965000000
1!
1%
#355970000000
0!
0%
#355975000000
1!
1%
#355980000000
0!
0%
#355985000000
1!
1%
#355990000000
0!
0%
#355995000000
1!
1%
#356000000000
0!
0%
#356005000000
1!
1%
#356010000000
0!
0%
#356015000000
1!
1%
#356020000000
0!
0%
#356025000000
1!
1%
#356030000000
0!
0%
#356035000000
1!
1%
#356040000000
0!
0%
#356045000000
1!
1%
#356050000000
0!
0%
#356055000000
1!
1%
#356060000000
0!
0%
#356065000000
1!
1%
#356070000000
0!
0%
#356075000000
1!
1%
#356080000000
0!
0%
#356085000000
1!
1%
#356090000000
0!
0%
#356095000000
1!
1%
#356100000000
0!
0%
#356105000000
1!
1%
#356110000000
0!
0%
#356115000000
1!
1%
#356120000000
0!
0%
#356125000000
1!
1%
#356130000000
0!
0%
#356135000000
1!
1%
#356140000000
0!
0%
#356145000000
1!
1%
#356150000000
0!
0%
#356155000000
1!
1%
#356160000000
0!
0%
#356165000000
1!
1%
#356170000000
0!
0%
#356175000000
1!
1%
#356180000000
0!
0%
#356185000000
1!
1%
#356190000000
0!
0%
#356195000000
1!
1%
#356200000000
0!
0%
#356205000000
1!
1%
#356210000000
0!
0%
#356215000000
1!
1%
#356220000000
0!
0%
#356225000000
1!
1%
#356230000000
0!
0%
#356235000000
1!
1%
#356240000000
0!
0%
#356245000000
1!
1%
#356250000000
0!
0%
#356255000000
1!
1%
#356260000000
0!
0%
#356265000000
1!
1%
#356270000000
0!
0%
#356275000000
1!
1%
#356280000000
0!
0%
#356285000000
1!
1%
#356290000000
0!
0%
#356295000000
1!
1%
#356300000000
0!
0%
#356305000000
1!
1%
#356310000000
0!
0%
#356315000000
1!
1%
#356320000000
0!
0%
#356325000000
1!
1%
#356330000000
0!
0%
#356335000000
1!
1%
#356340000000
0!
0%
#356345000000
1!
1%
#356350000000
0!
0%
#356355000000
1!
1%
#356360000000
0!
0%
#356365000000
1!
1%
#356370000000
0!
0%
#356375000000
1!
1%
#356380000000
0!
0%
#356385000000
1!
1%
#356390000000
0!
0%
#356395000000
1!
1%
#356400000000
0!
0%
#356405000000
1!
1%
#356410000000
0!
0%
#356415000000
1!
1%
#356420000000
0!
0%
#356425000000
1!
1%
#356430000000
0!
0%
#356435000000
1!
1%
#356440000000
0!
0%
#356445000000
1!
1%
#356450000000
0!
0%
#356455000000
1!
1%
#356460000000
0!
0%
#356465000000
1!
1%
#356470000000
0!
0%
#356475000000
1!
1%
#356480000000
0!
0%
#356485000000
1!
1%
#356490000000
0!
0%
#356495000000
1!
1%
#356500000000
0!
0%
#356505000000
1!
1%
#356510000000
0!
0%
#356515000000
1!
1%
#356520000000
0!
0%
#356525000000
1!
1%
#356530000000
0!
0%
#356535000000
1!
1%
#356540000000
0!
0%
#356545000000
1!
1%
#356550000000
0!
0%
#356555000000
1!
1%
#356560000000
0!
0%
#356565000000
1!
1%
#356570000000
0!
0%
#356575000000
1!
1%
#356580000000
0!
0%
#356585000000
1!
1%
#356590000000
0!
0%
#356595000000
1!
1%
#356600000000
0!
0%
#356605000000
1!
1%
#356610000000
0!
0%
#356615000000
1!
1%
#356620000000
0!
0%
#356625000000
1!
1%
#356630000000
0!
0%
#356635000000
1!
1%
#356640000000
0!
0%
#356645000000
1!
1%
#356650000000
0!
0%
#356655000000
1!
1%
#356660000000
0!
0%
#356665000000
1!
1%
#356670000000
0!
0%
#356675000000
1!
1%
#356680000000
0!
0%
#356685000000
1!
1%
#356690000000
0!
0%
#356695000000
1!
1%
#356700000000
0!
0%
#356705000000
1!
1%
#356710000000
0!
0%
#356715000000
1!
1%
#356720000000
0!
0%
#356725000000
1!
1%
#356730000000
0!
0%
#356735000000
1!
1%
#356740000000
0!
0%
#356745000000
1!
1%
#356750000000
0!
0%
#356755000000
1!
1%
#356760000000
0!
0%
#356765000000
1!
1%
#356770000000
0!
0%
#356775000000
1!
1%
#356780000000
0!
0%
#356785000000
1!
1%
#356790000000
0!
0%
#356795000000
1!
1%
#356800000000
0!
0%
#356805000000
1!
1%
#356810000000
0!
0%
#356815000000
1!
1%
#356820000000
0!
0%
#356825000000
1!
1%
#356830000000
0!
0%
#356835000000
1!
1%
#356840000000
0!
0%
#356845000000
1!
1%
#356850000000
0!
0%
#356855000000
1!
1%
#356860000000
0!
0%
#356865000000
1!
1%
#356870000000
0!
0%
#356875000000
1!
1%
#356880000000
0!
0%
#356885000000
1!
1%
#356890000000
0!
0%
#356895000000
1!
1%
#356900000000
0!
0%
#356905000000
1!
1%
#356910000000
0!
0%
#356915000000
1!
1%
#356920000000
0!
0%
#356925000000
1!
1%
#356930000000
0!
0%
#356935000000
1!
1%
#356940000000
0!
0%
#356945000000
1!
1%
#356950000000
0!
0%
#356955000000
1!
1%
#356960000000
0!
0%
#356965000000
1!
1%
#356970000000
0!
0%
#356975000000
1!
1%
#356980000000
0!
0%
#356985000000
1!
1%
#356990000000
0!
0%
#356995000000
1!
1%
#357000000000
0!
0%
#357005000000
1!
1%
#357010000000
0!
0%
#357015000000
1!
1%
#357020000000
0!
0%
#357025000000
1!
1%
#357030000000
0!
0%
#357035000000
1!
1%
#357040000000
0!
0%
#357045000000
1!
1%
#357050000000
0!
0%
#357055000000
1!
1%
#357060000000
0!
0%
#357065000000
1!
1%
#357070000000
0!
0%
#357075000000
1!
1%
#357080000000
0!
0%
#357085000000
1!
1%
#357090000000
0!
0%
#357095000000
1!
1%
#357100000000
0!
0%
#357105000000
1!
1%
#357110000000
0!
0%
#357115000000
1!
1%
#357120000000
0!
0%
#357125000000
1!
1%
#357130000000
0!
0%
#357135000000
1!
1%
#357140000000
0!
0%
#357145000000
1!
1%
#357150000000
0!
0%
#357155000000
1!
1%
#357160000000
0!
0%
#357165000000
1!
1%
#357170000000
0!
0%
#357175000000
1!
1%
#357180000000
0!
0%
#357185000000
1!
1%
#357190000000
0!
0%
#357195000000
1!
1%
#357200000000
0!
0%
#357205000000
1!
1%
#357210000000
0!
0%
#357215000000
1!
1%
#357220000000
0!
0%
#357225000000
1!
1%
#357230000000
0!
0%
#357235000000
1!
1%
#357240000000
0!
0%
#357245000000
1!
1%
#357250000000
0!
0%
#357255000000
1!
1%
#357260000000
0!
0%
#357265000000
1!
1%
#357270000000
0!
0%
#357275000000
1!
1%
#357280000000
0!
0%
#357285000000
1!
1%
#357290000000
0!
0%
#357295000000
1!
1%
#357300000000
0!
0%
#357305000000
1!
1%
#357310000000
0!
0%
#357315000000
1!
1%
#357320000000
0!
0%
#357325000000
1!
1%
#357330000000
0!
0%
#357335000000
1!
1%
#357340000000
0!
0%
#357345000000
1!
1%
#357350000000
0!
0%
#357355000000
1!
1%
#357360000000
0!
0%
#357365000000
1!
1%
#357370000000
0!
0%
#357375000000
1!
1%
#357380000000
0!
0%
#357385000000
1!
1%
#357390000000
0!
0%
#357395000000
1!
1%
#357400000000
0!
0%
#357405000000
1!
1%
#357410000000
0!
0%
#357415000000
1!
1%
#357420000000
0!
0%
#357425000000
1!
1%
#357430000000
0!
0%
#357435000000
1!
1%
#357440000000
0!
0%
#357445000000
1!
1%
#357450000000
0!
0%
#357455000000
1!
1%
#357460000000
0!
0%
#357465000000
1!
1%
#357470000000
0!
0%
#357475000000
1!
1%
#357480000000
0!
0%
#357485000000
1!
1%
#357490000000
0!
0%
#357495000000
1!
1%
#357500000000
0!
0%
#357505000000
1!
1%
#357510000000
0!
0%
#357515000000
1!
1%
#357520000000
0!
0%
#357525000000
1!
1%
#357530000000
0!
0%
#357535000000
1!
1%
#357540000000
0!
0%
#357545000000
1!
1%
#357550000000
0!
0%
#357555000000
1!
1%
#357560000000
0!
0%
#357565000000
1!
1%
#357570000000
0!
0%
#357575000000
1!
1%
#357580000000
0!
0%
#357585000000
1!
1%
#357590000000
0!
0%
#357595000000
1!
1%
#357600000000
0!
0%
#357605000000
1!
1%
#357610000000
0!
0%
#357615000000
1!
1%
#357620000000
0!
0%
#357625000000
1!
1%
#357630000000
0!
0%
#357635000000
1!
1%
#357640000000
0!
0%
#357645000000
1!
1%
#357650000000
0!
0%
#357655000000
1!
1%
#357660000000
0!
0%
#357665000000
1!
1%
#357670000000
0!
0%
#357675000000
1!
1%
#357680000000
0!
0%
#357685000000
1!
1%
#357690000000
0!
0%
#357695000000
1!
1%
#357700000000
0!
0%
#357705000000
1!
1%
#357710000000
0!
0%
#357715000000
1!
1%
#357720000000
0!
0%
#357725000000
1!
1%
#357730000000
0!
0%
#357735000000
1!
1%
#357740000000
0!
0%
#357745000000
1!
1%
#357750000000
0!
0%
#357755000000
1!
1%
#357760000000
0!
0%
#357765000000
1!
1%
#357770000000
0!
0%
#357775000000
1!
1%
#357780000000
0!
0%
#357785000000
1!
1%
#357790000000
0!
0%
#357795000000
1!
1%
#357800000000
0!
0%
#357805000000
1!
1%
#357810000000
0!
0%
#357815000000
1!
1%
#357820000000
0!
0%
#357825000000
1!
1%
#357830000000
0!
0%
#357835000000
1!
1%
#357840000000
0!
0%
#357845000000
1!
1%
#357850000000
0!
0%
#357855000000
1!
1%
#357860000000
0!
0%
#357865000000
1!
1%
#357870000000
0!
0%
#357875000000
1!
1%
#357880000000
0!
0%
#357885000000
1!
1%
#357890000000
0!
0%
#357895000000
1!
1%
#357900000000
0!
0%
#357905000000
1!
1%
#357910000000
0!
0%
#357915000000
1!
1%
#357920000000
0!
0%
#357925000000
1!
1%
#357930000000
0!
0%
#357935000000
1!
1%
#357940000000
0!
0%
#357945000000
1!
1%
#357950000000
0!
0%
#357955000000
1!
1%
#357960000000
0!
0%
#357965000000
1!
1%
#357970000000
0!
0%
#357975000000
1!
1%
#357980000000
0!
0%
#357985000000
1!
1%
#357990000000
0!
0%
#357995000000
1!
1%
#358000000000
0!
0%
#358005000000
1!
1%
#358010000000
0!
0%
#358015000000
1!
1%
#358020000000
0!
0%
#358025000000
1!
1%
#358030000000
0!
0%
#358035000000
1!
1%
#358040000000
0!
0%
#358045000000
1!
1%
#358050000000
0!
0%
#358055000000
1!
1%
#358060000000
0!
0%
#358065000000
1!
1%
#358070000000
0!
0%
#358075000000
1!
1%
#358080000000
0!
0%
#358085000000
1!
1%
#358090000000
0!
0%
#358095000000
1!
1%
#358100000000
0!
0%
#358105000000
1!
1%
#358110000000
0!
0%
#358115000000
1!
1%
#358120000000
0!
0%
#358125000000
1!
1%
#358130000000
0!
0%
#358135000000
1!
1%
#358140000000
0!
0%
#358145000000
1!
1%
#358150000000
0!
0%
#358155000000
1!
1%
#358160000000
0!
0%
#358165000000
1!
1%
#358170000000
0!
0%
#358175000000
1!
1%
#358180000000
0!
0%
#358185000000
1!
1%
#358190000000
0!
0%
#358195000000
1!
1%
#358200000000
0!
0%
#358205000000
1!
1%
#358210000000
0!
0%
#358215000000
1!
1%
#358220000000
0!
0%
#358225000000
1!
1%
#358230000000
0!
0%
#358235000000
1!
1%
#358240000000
0!
0%
#358245000000
1!
1%
#358250000000
0!
0%
#358255000000
1!
1%
#358260000000
0!
0%
#358265000000
1!
1%
#358270000000
0!
0%
#358275000000
1!
1%
#358280000000
0!
0%
#358285000000
1!
1%
#358290000000
0!
0%
#358295000000
1!
1%
#358300000000
0!
0%
#358305000000
1!
1%
#358310000000
0!
0%
#358315000000
1!
1%
#358320000000
0!
0%
#358325000000
1!
1%
#358330000000
0!
0%
#358335000000
1!
1%
#358340000000
0!
0%
#358345000000
1!
1%
#358350000000
0!
0%
#358355000000
1!
1%
#358360000000
0!
0%
#358365000000
1!
1%
#358370000000
0!
0%
#358375000000
1!
1%
#358380000000
0!
0%
#358385000000
1!
1%
#358390000000
0!
0%
#358395000000
1!
1%
#358400000000
0!
0%
#358405000000
1!
1%
#358410000000
0!
0%
#358415000000
1!
1%
#358420000000
0!
0%
#358425000000
1!
1%
#358430000000
0!
0%
#358435000000
1!
1%
#358440000000
0!
0%
#358445000000
1!
1%
#358450000000
0!
0%
#358455000000
1!
1%
#358460000000
0!
0%
#358465000000
1!
1%
#358470000000
0!
0%
#358475000000
1!
1%
#358480000000
0!
0%
#358485000000
1!
1%
#358490000000
0!
0%
#358495000000
1!
1%
#358500000000
0!
0%
#358505000000
1!
1%
#358510000000
0!
0%
#358515000000
1!
1%
#358520000000
0!
0%
#358525000000
1!
1%
#358530000000
0!
0%
#358535000000
1!
1%
#358540000000
0!
0%
#358545000000
1!
1%
#358550000000
0!
0%
#358555000000
1!
1%
#358560000000
0!
0%
#358565000000
1!
1%
#358570000000
0!
0%
#358575000000
1!
1%
#358580000000
0!
0%
#358585000000
1!
1%
#358590000000
0!
0%
#358595000000
1!
1%
#358600000000
0!
0%
#358605000000
1!
1%
#358610000000
0!
0%
#358615000000
1!
1%
#358620000000
0!
0%
#358625000000
1!
1%
#358630000000
0!
0%
#358635000000
1!
1%
#358640000000
0!
0%
#358645000000
1!
1%
#358650000000
0!
0%
#358655000000
1!
1%
#358660000000
0!
0%
#358665000000
1!
1%
#358670000000
0!
0%
#358675000000
1!
1%
#358680000000
0!
0%
#358685000000
1!
1%
#358690000000
0!
0%
#358695000000
1!
1%
#358700000000
0!
0%
#358705000000
1!
1%
#358710000000
0!
0%
#358715000000
1!
1%
#358720000000
0!
0%
#358725000000
1!
1%
#358730000000
0!
0%
#358735000000
1!
1%
#358740000000
0!
0%
#358745000000
1!
1%
#358750000000
0!
0%
#358755000000
1!
1%
#358760000000
0!
0%
#358765000000
1!
1%
#358770000000
0!
0%
#358775000000
1!
1%
#358780000000
0!
0%
#358785000000
1!
1%
#358790000000
0!
0%
#358795000000
1!
1%
#358800000000
0!
0%
#358805000000
1!
1%
#358810000000
0!
0%
#358815000000
1!
1%
#358820000000
0!
0%
#358825000000
1!
1%
#358830000000
0!
0%
#358835000000
1!
1%
#358840000000
0!
0%
#358845000000
1!
1%
#358850000000
0!
0%
#358855000000
1!
1%
#358860000000
0!
0%
#358865000000
1!
1%
#358870000000
0!
0%
#358875000000
1!
1%
#358880000000
0!
0%
#358885000000
1!
1%
#358890000000
0!
0%
#358895000000
1!
1%
#358900000000
0!
0%
#358905000000
1!
1%
#358910000000
0!
0%
#358915000000
1!
1%
#358920000000
0!
0%
#358925000000
1!
1%
#358930000000
0!
0%
#358935000000
1!
1%
#358940000000
0!
0%
#358945000000
1!
1%
#358950000000
0!
0%
#358955000000
1!
1%
#358960000000
0!
0%
#358965000000
1!
1%
#358970000000
0!
0%
#358975000000
1!
1%
#358980000000
0!
0%
#358985000000
1!
1%
#358990000000
0!
0%
#358995000000
1!
1%
#359000000000
0!
0%
#359005000000
1!
1%
#359010000000
0!
0%
#359015000000
1!
1%
#359020000000
0!
0%
#359025000000
1!
1%
#359030000000
0!
0%
#359035000000
1!
1%
#359040000000
0!
0%
#359045000000
1!
1%
#359050000000
0!
0%
#359055000000
1!
1%
#359060000000
0!
0%
#359065000000
1!
1%
#359070000000
0!
0%
#359075000000
1!
1%
#359080000000
0!
0%
#359085000000
1!
1%
#359090000000
0!
0%
#359095000000
1!
1%
#359100000000
0!
0%
#359105000000
1!
1%
#359110000000
0!
0%
#359115000000
1!
1%
#359120000000
0!
0%
#359125000000
1!
1%
#359130000000
0!
0%
#359135000000
1!
1%
#359140000000
0!
0%
#359145000000
1!
1%
#359150000000
0!
0%
#359155000000
1!
1%
#359160000000
0!
0%
#359165000000
1!
1%
#359170000000
0!
0%
#359175000000
1!
1%
#359180000000
0!
0%
#359185000000
1!
1%
#359190000000
0!
0%
#359195000000
1!
1%
#359200000000
0!
0%
#359205000000
1!
1%
#359210000000
0!
0%
#359215000000
1!
1%
#359220000000
0!
0%
#359225000000
1!
1%
#359230000000
0!
0%
#359235000000
1!
1%
#359240000000
0!
0%
#359245000000
1!
1%
#359250000000
0!
0%
#359255000000
1!
1%
#359260000000
0!
0%
#359265000000
1!
1%
#359270000000
0!
0%
#359275000000
1!
1%
#359280000000
0!
0%
#359285000000
1!
1%
#359290000000
0!
0%
#359295000000
1!
1%
#359300000000
0!
0%
#359305000000
1!
1%
#359310000000
0!
0%
#359315000000
1!
1%
#359320000000
0!
0%
#359325000000
1!
1%
#359330000000
0!
0%
#359335000000
1!
1%
#359340000000
0!
0%
#359345000000
1!
1%
#359350000000
0!
0%
#359355000000
1!
1%
#359360000000
0!
0%
#359365000000
1!
1%
#359370000000
0!
0%
#359375000000
1!
1%
#359380000000
0!
0%
#359385000000
1!
1%
#359390000000
0!
0%
#359395000000
1!
1%
#359400000000
0!
0%
#359405000000
1!
1%
#359410000000
0!
0%
#359415000000
1!
1%
#359420000000
0!
0%
#359425000000
1!
1%
#359430000000
0!
0%
#359435000000
1!
1%
#359440000000
0!
0%
#359445000000
1!
1%
#359450000000
0!
0%
#359455000000
1!
1%
#359460000000
0!
0%
#359465000000
1!
1%
#359470000000
0!
0%
#359475000000
1!
1%
#359480000000
0!
0%
#359485000000
1!
1%
#359490000000
0!
0%
#359495000000
1!
1%
#359500000000
0!
0%
#359505000000
1!
1%
#359510000000
0!
0%
#359515000000
1!
1%
#359520000000
0!
0%
#359525000000
1!
1%
#359530000000
0!
0%
#359535000000
1!
1%
#359540000000
0!
0%
#359545000000
1!
1%
#359550000000
0!
0%
#359555000000
1!
1%
#359560000000
0!
0%
#359565000000
1!
1%
#359570000000
0!
0%
#359575000000
1!
1%
#359580000000
0!
0%
#359585000000
1!
1%
#359590000000
0!
0%
#359595000000
1!
1%
#359600000000
0!
0%
#359605000000
1!
1%
#359610000000
0!
0%
#359615000000
1!
1%
#359620000000
0!
0%
#359625000000
1!
1%
#359630000000
0!
0%
#359635000000
1!
1%
#359640000000
0!
0%
#359645000000
1!
1%
#359650000000
0!
0%
#359655000000
1!
1%
#359660000000
0!
0%
#359665000000
1!
1%
#359670000000
0!
0%
#359675000000
1!
1%
#359680000000
0!
0%
#359685000000
1!
1%
#359690000000
0!
0%
#359695000000
1!
1%
#359700000000
0!
0%
#359705000000
1!
1%
#359710000000
0!
0%
#359715000000
1!
1%
#359720000000
0!
0%
#359725000000
1!
1%
#359730000000
0!
0%
#359735000000
1!
1%
#359740000000
0!
0%
#359745000000
1!
1%
#359750000000
0!
0%
#359755000000
1!
1%
#359760000000
0!
0%
#359765000000
1!
1%
#359770000000
0!
0%
#359775000000
1!
1%
#359780000000
0!
0%
#359785000000
1!
1%
#359790000000
0!
0%
#359795000000
1!
1%
#359800000000
0!
0%
#359805000000
1!
1%
#359810000000
0!
0%
#359815000000
1!
1%
#359820000000
0!
0%
#359825000000
1!
1%
#359830000000
0!
0%
#359835000000
1!
1%
#359840000000
0!
0%
#359845000000
1!
1%
#359850000000
0!
0%
#359855000000
1!
1%
#359860000000
0!
0%
#359865000000
1!
1%
#359870000000
0!
0%
#359875000000
1!
1%
#359880000000
0!
0%
#359885000000
1!
1%
#359890000000
0!
0%
#359895000000
1!
1%
#359900000000
0!
0%
#359905000000
1!
1%
#359910000000
0!
0%
#359915000000
1!
1%
#359920000000
0!
0%
#359925000000
1!
1%
#359930000000
0!
0%
#359935000000
1!
1%
#359940000000
0!
0%
#359945000000
1!
1%
#359950000000
0!
0%
#359955000000
1!
1%
#359960000000
0!
0%
#359965000000
1!
1%
#359970000000
0!
0%
#359975000000
1!
1%
#359980000000
0!
0%
#359985000000
1!
1%
#359990000000
0!
0%
#359995000000
1!
1%
#360000000000
0!
0%
#360005000000
1!
1%
#360010000000
0!
0%
#360015000000
1!
1%
#360020000000
0!
0%
#360025000000
1!
1%
#360030000000
0!
0%
#360035000000
1!
1%
#360040000000
0!
0%
#360045000000
1!
1%
#360050000000
0!
0%
#360055000000
1!
1%
#360060000000
0!
0%
#360065000000
1!
1%
#360070000000
0!
0%
#360075000000
1!
1%
#360080000000
0!
0%
#360085000000
1!
1%
#360090000000
0!
0%
#360095000000
1!
1%
#360100000000
0!
0%
#360105000000
1!
1%
#360110000000
0!
0%
#360115000000
1!
1%
#360120000000
0!
0%
#360125000000
1!
1%
#360130000000
0!
0%
#360135000000
1!
1%
#360140000000
0!
0%
#360145000000
1!
1%
#360150000000
0!
0%
#360155000000
1!
1%
#360160000000
0!
0%
#360165000000
1!
1%
#360170000000
0!
0%
#360175000000
1!
1%
#360180000000
0!
0%
#360185000000
1!
1%
#360190000000
0!
0%
#360195000000
1!
1%
#360200000000
0!
0%
#360205000000
1!
1%
#360210000000
0!
0%
#360215000000
1!
1%
#360220000000
0!
0%
#360225000000
1!
1%
#360230000000
0!
0%
#360235000000
1!
1%
#360240000000
0!
0%
#360245000000
1!
1%
#360250000000
0!
0%
#360255000000
1!
1%
#360260000000
0!
0%
#360265000000
1!
1%
#360270000000
0!
0%
#360275000000
1!
1%
#360280000000
0!
0%
#360285000000
1!
1%
#360290000000
0!
0%
#360295000000
1!
1%
#360300000000
0!
0%
#360305000000
1!
1%
#360310000000
0!
0%
#360315000000
1!
1%
#360320000000
0!
0%
#360325000000
1!
1%
#360330000000
0!
0%
#360335000000
1!
1%
#360340000000
0!
0%
#360345000000
1!
1%
#360350000000
0!
0%
#360355000000
1!
1%
#360360000000
0!
0%
#360365000000
1!
1%
#360370000000
0!
0%
#360375000000
1!
1%
#360380000000
0!
0%
#360385000000
1!
1%
#360390000000
0!
0%
#360395000000
1!
1%
#360400000000
0!
0%
#360405000000
1!
1%
#360410000000
0!
0%
#360415000000
1!
1%
#360420000000
0!
0%
#360425000000
1!
1%
#360430000000
0!
0%
#360435000000
1!
1%
#360440000000
0!
0%
#360445000000
1!
1%
#360450000000
0!
0%
#360455000000
1!
1%
#360460000000
0!
0%
#360465000000
1!
1%
#360470000000
0!
0%
#360475000000
1!
1%
#360480000000
0!
0%
#360485000000
1!
1%
#360490000000
0!
0%
#360495000000
1!
1%
#360500000000
0!
0%
#360505000000
1!
1%
#360510000000
0!
0%
#360515000000
1!
1%
#360520000000
0!
0%
#360525000000
1!
1%
#360530000000
0!
0%
#360535000000
1!
1%
#360540000000
0!
0%
#360545000000
1!
1%
#360550000000
0!
0%
#360555000000
1!
1%
#360560000000
0!
0%
#360565000000
1!
1%
#360570000000
0!
0%
#360575000000
1!
1%
#360580000000
0!
0%
#360585000000
1!
1%
#360590000000
0!
0%
#360595000000
1!
1%
#360600000000
0!
0%
#360605000000
1!
1%
#360610000000
0!
0%
#360615000000
1!
1%
#360620000000
0!
0%
#360625000000
1!
1%
#360630000000
0!
0%
#360635000000
1!
1%
#360640000000
0!
0%
#360645000000
1!
1%
#360650000000
0!
0%
#360655000000
1!
1%
#360660000000
0!
0%
#360665000000
1!
1%
#360670000000
0!
0%
#360675000000
1!
1%
#360680000000
0!
0%
#360685000000
1!
1%
#360690000000
0!
0%
#360695000000
1!
1%
#360700000000
0!
0%
#360705000000
1!
1%
#360710000000
0!
0%
#360715000000
1!
1%
#360720000000
0!
0%
#360725000000
1!
1%
#360730000000
0!
0%
#360735000000
1!
1%
#360740000000
0!
0%
#360745000000
1!
1%
#360750000000
0!
0%
#360755000000
1!
1%
#360760000000
0!
0%
#360765000000
1!
1%
#360770000000
0!
0%
#360775000000
1!
1%
#360780000000
0!
0%
#360785000000
1!
1%
#360790000000
0!
0%
#360795000000
1!
1%
#360800000000
0!
0%
#360805000000
1!
1%
#360810000000
0!
0%
#360815000000
1!
1%
#360820000000
0!
0%
#360825000000
1!
1%
#360830000000
0!
0%
#360835000000
1!
1%
#360840000000
0!
0%
#360845000000
1!
1%
#360850000000
0!
0%
#360855000000
1!
1%
#360860000000
0!
0%
#360865000000
1!
1%
#360870000000
0!
0%
#360875000000
1!
1%
#360880000000
0!
0%
#360885000000
1!
1%
#360890000000
0!
0%
#360895000000
1!
1%
#360900000000
0!
0%
#360905000000
1!
1%
#360910000000
0!
0%
#360915000000
1!
1%
#360920000000
0!
0%
#360925000000
1!
1%
#360930000000
0!
0%
#360935000000
1!
1%
#360940000000
0!
0%
#360945000000
1!
1%
#360950000000
0!
0%
#360955000000
1!
1%
#360960000000
0!
0%
#360965000000
1!
1%
#360970000000
0!
0%
#360975000000
1!
1%
#360980000000
0!
0%
#360985000000
1!
1%
#360990000000
0!
0%
#360995000000
1!
1%
#361000000000
0!
0%
#361005000000
1!
1%
#361010000000
0!
0%
#361015000000
1!
1%
#361020000000
0!
0%
#361025000000
1!
1%
#361030000000
0!
0%
#361035000000
1!
1%
#361040000000
0!
0%
#361045000000
1!
1%
#361050000000
0!
0%
#361055000000
1!
1%
#361060000000
0!
0%
#361065000000
1!
1%
#361070000000
0!
0%
#361075000000
1!
1%
#361080000000
0!
0%
#361085000000
1!
1%
#361090000000
0!
0%
#361095000000
1!
1%
#361100000000
0!
0%
#361105000000
1!
1%
#361110000000
0!
0%
#361115000000
1!
1%
#361120000000
0!
0%
#361125000000
1!
1%
#361130000000
0!
0%
#361135000000
1!
1%
#361140000000
0!
0%
#361145000000
1!
1%
#361150000000
0!
0%
#361155000000
1!
1%
#361160000000
0!
0%
#361165000000
1!
1%
#361170000000
0!
0%
#361175000000
1!
1%
#361180000000
0!
0%
#361185000000
1!
1%
#361190000000
0!
0%
#361195000000
1!
1%
#361200000000
0!
0%
#361205000000
1!
1%
#361210000000
0!
0%
#361215000000
1!
1%
#361220000000
0!
0%
#361225000000
1!
1%
#361230000000
0!
0%
#361235000000
1!
1%
#361240000000
0!
0%
#361245000000
1!
1%
#361250000000
0!
0%
#361255000000
1!
1%
#361260000000
0!
0%
#361265000000
1!
1%
#361270000000
0!
0%
#361275000000
1!
1%
#361280000000
0!
0%
#361285000000
1!
1%
#361290000000
0!
0%
#361295000000
1!
1%
#361300000000
0!
0%
#361305000000
1!
1%
#361310000000
0!
0%
#361315000000
1!
1%
#361320000000
0!
0%
#361325000000
1!
1%
#361330000000
0!
0%
#361335000000
1!
1%
#361340000000
0!
0%
#361345000000
1!
1%
#361350000000
0!
0%
#361355000000
1!
1%
#361360000000
0!
0%
#361365000000
1!
1%
#361370000000
0!
0%
#361375000000
1!
1%
#361380000000
0!
0%
#361385000000
1!
1%
#361390000000
0!
0%
#361395000000
1!
1%
#361400000000
0!
0%
#361405000000
1!
1%
#361410000000
0!
0%
#361415000000
1!
1%
#361420000000
0!
0%
#361425000000
1!
1%
#361430000000
0!
0%
#361435000000
1!
1%
#361440000000
0!
0%
#361445000000
1!
1%
#361450000000
0!
0%
#361455000000
1!
1%
#361460000000
0!
0%
#361465000000
1!
1%
#361470000000
0!
0%
#361475000000
1!
1%
#361480000000
0!
0%
#361485000000
1!
1%
#361490000000
0!
0%
#361495000000
1!
1%
#361500000000
0!
0%
#361505000000
1!
1%
#361510000000
0!
0%
#361515000000
1!
1%
#361520000000
0!
0%
#361525000000
1!
1%
#361530000000
0!
0%
#361535000000
1!
1%
#361540000000
0!
0%
#361545000000
1!
1%
#361550000000
0!
0%
#361555000000
1!
1%
#361560000000
0!
0%
#361565000000
1!
1%
#361570000000
0!
0%
#361575000000
1!
1%
#361580000000
0!
0%
#361585000000
1!
1%
#361590000000
0!
0%
#361595000000
1!
1%
#361600000000
0!
0%
#361605000000
1!
1%
#361610000000
0!
0%
#361615000000
1!
1%
#361620000000
0!
0%
#361625000000
1!
1%
#361630000000
0!
0%
#361635000000
1!
1%
#361640000000
0!
0%
#361645000000
1!
1%
#361650000000
0!
0%
#361655000000
1!
1%
#361660000000
0!
0%
#361665000000
1!
1%
#361670000000
0!
0%
#361675000000
1!
1%
#361680000000
0!
0%
#361685000000
1!
1%
#361690000000
0!
0%
#361695000000
1!
1%
#361700000000
0!
0%
#361705000000
1!
1%
#361710000000
0!
0%
#361715000000
1!
1%
#361720000000
0!
0%
#361725000000
1!
1%
#361730000000
0!
0%
#361735000000
1!
1%
#361740000000
0!
0%
#361745000000
1!
1%
#361750000000
0!
0%
#361755000000
1!
1%
#361760000000
0!
0%
#361765000000
1!
1%
#361770000000
0!
0%
#361775000000
1!
1%
#361780000000
0!
0%
#361785000000
1!
1%
#361790000000
0!
0%
#361795000000
1!
1%
#361800000000
0!
0%
#361805000000
1!
1%
#361810000000
0!
0%
#361815000000
1!
1%
#361820000000
0!
0%
#361825000000
1!
1%
#361830000000
0!
0%
#361835000000
1!
1%
#361840000000
0!
0%
#361845000000
1!
1%
#361850000000
0!
0%
#361855000000
1!
1%
#361860000000
0!
0%
#361865000000
1!
1%
#361870000000
0!
0%
#361875000000
1!
1%
#361880000000
0!
0%
#361885000000
1!
1%
#361890000000
0!
0%
#361895000000
1!
1%
#361900000000
0!
0%
#361905000000
1!
1%
#361910000000
0!
0%
#361915000000
1!
1%
#361920000000
0!
0%
#361925000000
1!
1%
#361930000000
0!
0%
#361935000000
1!
1%
#361940000000
0!
0%
#361945000000
1!
1%
#361950000000
0!
0%
#361955000000
1!
1%
#361960000000
0!
0%
#361965000000
1!
1%
#361970000000
0!
0%
#361975000000
1!
1%
#361980000000
0!
0%
#361985000000
1!
1%
#361990000000
0!
0%
#361995000000
1!
1%
#362000000000
0!
0%
#362005000000
1!
1%
#362010000000
0!
0%
#362015000000
1!
1%
#362020000000
0!
0%
#362025000000
1!
1%
#362030000000
0!
0%
#362035000000
1!
1%
#362040000000
0!
0%
#362045000000
1!
1%
#362050000000
0!
0%
#362055000000
1!
1%
#362060000000
0!
0%
#362065000000
1!
1%
#362070000000
0!
0%
#362075000000
1!
1%
#362080000000
0!
0%
#362085000000
1!
1%
#362090000000
0!
0%
#362095000000
1!
1%
#362100000000
0!
0%
#362105000000
1!
1%
#362110000000
0!
0%
#362115000000
1!
1%
#362120000000
0!
0%
#362125000000
1!
1%
#362130000000
0!
0%
#362135000000
1!
1%
#362140000000
0!
0%
#362145000000
1!
1%
#362150000000
0!
0%
#362155000000
1!
1%
#362160000000
0!
0%
#362165000000
1!
1%
#362170000000
0!
0%
#362175000000
1!
1%
#362180000000
0!
0%
#362185000000
1!
1%
#362190000000
0!
0%
#362195000000
1!
1%
#362200000000
0!
0%
#362205000000
1!
1%
#362210000000
0!
0%
#362215000000
1!
1%
#362220000000
0!
0%
#362225000000
1!
1%
#362230000000
0!
0%
#362235000000
1!
1%
#362240000000
0!
0%
#362245000000
1!
1%
#362250000000
0!
0%
#362255000000
1!
1%
#362260000000
0!
0%
#362265000000
1!
1%
#362270000000
0!
0%
#362275000000
1!
1%
#362280000000
0!
0%
#362285000000
1!
1%
#362290000000
0!
0%
#362295000000
1!
1%
#362300000000
0!
0%
#362305000000
1!
1%
#362310000000
0!
0%
#362315000000
1!
1%
#362320000000
0!
0%
#362325000000
1!
1%
#362330000000
0!
0%
#362335000000
1!
1%
#362340000000
0!
0%
#362345000000
1!
1%
#362350000000
0!
0%
#362355000000
1!
1%
#362360000000
0!
0%
#362365000000
1!
1%
#362370000000
0!
0%
#362375000000
1!
1%
#362380000000
0!
0%
#362385000000
1!
1%
#362390000000
0!
0%
#362395000000
1!
1%
#362400000000
0!
0%
#362405000000
1!
1%
#362410000000
0!
0%
#362415000000
1!
1%
#362420000000
0!
0%
#362425000000
1!
1%
#362430000000
0!
0%
#362435000000
1!
1%
#362440000000
0!
0%
#362445000000
1!
1%
#362450000000
0!
0%
#362455000000
1!
1%
#362460000000
0!
0%
#362465000000
1!
1%
#362470000000
0!
0%
#362475000000
1!
1%
#362480000000
0!
0%
#362485000000
1!
1%
#362490000000
0!
0%
#362495000000
1!
1%
#362500000000
0!
0%
#362505000000
1!
1%
#362510000000
0!
0%
#362515000000
1!
1%
#362520000000
0!
0%
#362525000000
1!
1%
#362530000000
0!
0%
#362535000000
1!
1%
#362540000000
0!
0%
#362545000000
1!
1%
#362550000000
0!
0%
#362555000000
1!
1%
#362560000000
0!
0%
#362565000000
1!
1%
#362570000000
0!
0%
#362575000000
1!
1%
#362580000000
0!
0%
#362585000000
1!
1%
#362590000000
0!
0%
#362595000000
1!
1%
#362600000000
0!
0%
#362605000000
1!
1%
#362610000000
0!
0%
#362615000000
1!
1%
#362620000000
0!
0%
#362625000000
1!
1%
#362630000000
0!
0%
#362635000000
1!
1%
#362640000000
0!
0%
#362645000000
1!
1%
#362650000000
0!
0%
#362655000000
1!
1%
#362660000000
0!
0%
#362665000000
1!
1%
#362670000000
0!
0%
#362675000000
1!
1%
#362680000000
0!
0%
#362685000000
1!
1%
#362690000000
0!
0%
#362695000000
1!
1%
#362700000000
0!
0%
#362705000000
1!
1%
#362710000000
0!
0%
#362715000000
1!
1%
#362720000000
0!
0%
#362725000000
1!
1%
#362730000000
0!
0%
#362735000000
1!
1%
#362740000000
0!
0%
#362745000000
1!
1%
#362750000000
0!
0%
#362755000000
1!
1%
#362760000000
0!
0%
#362765000000
1!
1%
#362770000000
0!
0%
#362775000000
1!
1%
#362780000000
0!
0%
#362785000000
1!
1%
#362790000000
0!
0%
#362795000000
1!
1%
#362800000000
0!
0%
#362805000000
1!
1%
#362810000000
0!
0%
#362815000000
1!
1%
#362820000000
0!
0%
#362825000000
1!
1%
#362830000000
0!
0%
#362835000000
1!
1%
#362840000000
0!
0%
#362845000000
1!
1%
#362850000000
0!
0%
#362855000000
1!
1%
#362860000000
0!
0%
#362865000000
1!
1%
#362870000000
0!
0%
#362875000000
1!
1%
#362880000000
0!
0%
#362885000000
1!
1%
#362890000000
0!
0%
#362895000000
1!
1%
#362900000000
0!
0%
#362905000000
1!
1%
#362910000000
0!
0%
#362915000000
1!
1%
#362920000000
0!
0%
#362925000000
1!
1%
#362930000000
0!
0%
#362935000000
1!
1%
#362940000000
0!
0%
#362945000000
1!
1%
#362950000000
0!
0%
#362955000000
1!
1%
#362960000000
0!
0%
#362965000000
1!
1%
#362970000000
0!
0%
#362975000000
1!
1%
#362980000000
0!
0%
#362985000000
1!
1%
#362990000000
0!
0%
#362995000000
1!
1%
#363000000000
0!
0%
#363005000000
1!
1%
#363010000000
0!
0%
#363015000000
1!
1%
#363020000000
0!
0%
#363025000000
1!
1%
#363030000000
0!
0%
#363035000000
1!
1%
#363040000000
0!
0%
#363045000000
1!
1%
#363050000000
0!
0%
#363055000000
1!
1%
#363060000000
0!
0%
#363065000000
1!
1%
#363070000000
0!
0%
#363075000000
1!
1%
#363080000000
0!
0%
#363085000000
1!
1%
#363090000000
0!
0%
#363095000000
1!
1%
#363100000000
0!
0%
#363105000000
1!
1%
#363110000000
0!
0%
#363115000000
1!
1%
#363120000000
0!
0%
#363125000000
1!
1%
#363130000000
0!
0%
#363135000000
1!
1%
#363140000000
0!
0%
#363145000000
1!
1%
#363150000000
0!
0%
#363155000000
1!
1%
#363160000000
0!
0%
#363165000000
1!
1%
#363170000000
0!
0%
#363175000000
1!
1%
#363180000000
0!
0%
#363185000000
1!
1%
#363190000000
0!
0%
#363195000000
1!
1%
#363200000000
0!
0%
#363205000000
1!
1%
#363210000000
0!
0%
#363215000000
1!
1%
#363220000000
0!
0%
#363225000000
1!
1%
#363230000000
0!
0%
#363235000000
1!
1%
#363240000000
0!
0%
#363245000000
1!
1%
#363250000000
0!
0%
#363255000000
1!
1%
#363260000000
0!
0%
#363265000000
1!
1%
#363270000000
0!
0%
#363275000000
1!
1%
#363280000000
0!
0%
#363285000000
1!
1%
#363290000000
0!
0%
#363295000000
1!
1%
#363300000000
0!
0%
#363305000000
1!
1%
#363310000000
0!
0%
#363315000000
1!
1%
#363320000000
0!
0%
#363325000000
1!
1%
#363330000000
0!
0%
#363335000000
1!
1%
#363340000000
0!
0%
#363345000000
1!
1%
#363350000000
0!
0%
#363355000000
1!
1%
#363360000000
0!
0%
#363365000000
1!
1%
#363370000000
0!
0%
#363375000000
1!
1%
#363380000000
0!
0%
#363385000000
1!
1%
#363390000000
0!
0%
#363395000000
1!
1%
#363400000000
0!
0%
#363405000000
1!
1%
#363410000000
0!
0%
#363415000000
1!
1%
#363420000000
0!
0%
#363425000000
1!
1%
#363430000000
0!
0%
#363435000000
1!
1%
#363440000000
0!
0%
#363445000000
1!
1%
#363450000000
0!
0%
#363455000000
1!
1%
#363460000000
0!
0%
#363465000000
1!
1%
#363470000000
0!
0%
#363475000000
1!
1%
#363480000000
0!
0%
#363485000000
1!
1%
#363490000000
0!
0%
#363495000000
1!
1%
#363500000000
0!
0%
#363505000000
1!
1%
#363510000000
0!
0%
#363515000000
1!
1%
#363520000000
0!
0%
#363525000000
1!
1%
#363530000000
0!
0%
#363535000000
1!
1%
#363540000000
0!
0%
#363545000000
1!
1%
#363550000000
0!
0%
#363555000000
1!
1%
#363560000000
0!
0%
#363565000000
1!
1%
#363570000000
0!
0%
#363575000000
1!
1%
#363580000000
0!
0%
#363585000000
1!
1%
#363590000000
0!
0%
#363595000000
1!
1%
#363600000000
0!
0%
#363605000000
1!
1%
#363610000000
0!
0%
#363615000000
1!
1%
#363620000000
0!
0%
#363625000000
1!
1%
#363630000000
0!
0%
#363635000000
1!
1%
#363640000000
0!
0%
#363645000000
1!
1%
#363650000000
0!
0%
#363655000000
1!
1%
#363660000000
0!
0%
#363665000000
1!
1%
#363670000000
0!
0%
#363675000000
1!
1%
#363680000000
0!
0%
#363685000000
1!
1%
#363690000000
0!
0%
#363695000000
1!
1%
#363700000000
0!
0%
#363705000000
1!
1%
#363710000000
0!
0%
#363715000000
1!
1%
#363720000000
0!
0%
#363725000000
1!
1%
#363730000000
0!
0%
#363735000000
1!
1%
#363740000000
0!
0%
#363745000000
1!
1%
#363750000000
0!
0%
#363755000000
1!
1%
#363760000000
0!
0%
#363765000000
1!
1%
#363770000000
0!
0%
#363775000000
1!
1%
#363780000000
0!
0%
#363785000000
1!
1%
#363790000000
0!
0%
#363795000000
1!
1%
#363800000000
0!
0%
#363805000000
1!
1%
#363810000000
0!
0%
#363815000000
1!
1%
#363820000000
0!
0%
#363825000000
1!
1%
#363830000000
0!
0%
#363835000000
1!
1%
#363840000000
0!
0%
#363845000000
1!
1%
#363850000000
0!
0%
#363855000000
1!
1%
#363860000000
0!
0%
#363865000000
1!
1%
#363870000000
0!
0%
#363875000000
1!
1%
#363880000000
0!
0%
#363885000000
1!
1%
#363890000000
0!
0%
#363895000000
1!
1%
#363900000000
0!
0%
#363905000000
1!
1%
#363910000000
0!
0%
#363915000000
1!
1%
#363920000000
0!
0%
#363925000000
1!
1%
#363930000000
0!
0%
#363935000000
1!
1%
#363940000000
0!
0%
#363945000000
1!
1%
#363950000000
0!
0%
#363955000000
1!
1%
#363960000000
0!
0%
#363965000000
1!
1%
#363970000000
0!
0%
#363975000000
1!
1%
#363980000000
0!
0%
#363985000000
1!
1%
#363990000000
0!
0%
#363995000000
1!
1%
#364000000000
0!
0%
#364005000000
1!
1%
#364010000000
0!
0%
#364015000000
1!
1%
#364020000000
0!
0%
#364025000000
1!
1%
#364030000000
0!
0%
#364035000000
1!
1%
#364040000000
0!
0%
#364045000000
1!
1%
#364050000000
0!
0%
#364055000000
1!
1%
#364060000000
0!
0%
#364065000000
1!
1%
#364070000000
0!
0%
#364075000000
1!
1%
#364080000000
0!
0%
#364085000000
1!
1%
#364090000000
0!
0%
#364095000000
1!
1%
#364100000000
0!
0%
#364105000000
1!
1%
#364110000000
0!
0%
#364115000000
1!
1%
#364120000000
0!
0%
#364125000000
1!
1%
#364130000000
0!
0%
#364135000000
1!
1%
#364140000000
0!
0%
#364145000000
1!
1%
#364150000000
0!
0%
#364155000000
1!
1%
#364160000000
0!
0%
#364165000000
1!
1%
#364170000000
0!
0%
#364175000000
1!
1%
#364180000000
0!
0%
#364185000000
1!
1%
#364190000000
0!
0%
#364195000000
1!
1%
#364200000000
0!
0%
#364205000000
1!
1%
#364210000000
0!
0%
#364215000000
1!
1%
#364220000000
0!
0%
#364225000000
1!
1%
#364230000000
0!
0%
#364235000000
1!
1%
#364240000000
0!
0%
#364245000000
1!
1%
#364250000000
0!
0%
#364255000000
1!
1%
#364260000000
0!
0%
#364265000000
1!
1%
#364270000000
0!
0%
#364275000000
1!
1%
#364280000000
0!
0%
#364285000000
1!
1%
#364290000000
0!
0%
#364295000000
1!
1%
#364300000000
0!
0%
#364305000000
1!
1%
#364310000000
0!
0%
#364315000000
1!
1%
#364320000000
0!
0%
#364325000000
1!
1%
#364330000000
0!
0%
#364335000000
1!
1%
#364340000000
0!
0%
#364345000000
1!
1%
#364350000000
0!
0%
#364355000000
1!
1%
#364360000000
0!
0%
#364365000000
1!
1%
#364370000000
0!
0%
#364375000000
1!
1%
#364380000000
0!
0%
#364385000000
1!
1%
#364390000000
0!
0%
#364395000000
1!
1%
#364400000000
0!
0%
#364405000000
1!
1%
#364410000000
0!
0%
#364415000000
1!
1%
#364420000000
0!
0%
#364425000000
1!
1%
#364430000000
0!
0%
#364435000000
1!
1%
#364440000000
0!
0%
#364445000000
1!
1%
#364450000000
0!
0%
#364455000000
1!
1%
#364460000000
0!
0%
#364465000000
1!
1%
#364470000000
0!
0%
#364475000000
1!
1%
#364480000000
0!
0%
#364485000000
1!
1%
#364490000000
0!
0%
#364495000000
1!
1%
#364500000000
0!
0%
#364505000000
1!
1%
#364510000000
0!
0%
#364515000000
1!
1%
#364520000000
0!
0%
#364525000000
1!
1%
#364530000000
0!
0%
#364535000000
1!
1%
#364540000000
0!
0%
#364545000000
1!
1%
#364550000000
0!
0%
#364555000000
1!
1%
#364560000000
0!
0%
#364565000000
1!
1%
#364570000000
0!
0%
#364575000000
1!
1%
#364580000000
0!
0%
#364585000000
1!
1%
#364590000000
0!
0%
#364595000000
1!
1%
#364600000000
0!
0%
#364605000000
1!
1%
#364610000000
0!
0%
#364615000000
1!
1%
#364620000000
0!
0%
#364625000000
1!
1%
#364630000000
0!
0%
#364635000000
1!
1%
#364640000000
0!
0%
#364645000000
1!
1%
#364650000000
0!
0%
#364655000000
1!
1%
#364660000000
0!
0%
#364665000000
1!
1%
#364670000000
0!
0%
#364675000000
1!
1%
#364680000000
0!
0%
#364685000000
1!
1%
#364690000000
0!
0%
#364695000000
1!
1%
#364700000000
0!
0%
#364705000000
1!
1%
#364710000000
0!
0%
#364715000000
1!
1%
#364720000000
0!
0%
#364725000000
1!
1%
#364730000000
0!
0%
#364735000000
1!
1%
#364740000000
0!
0%
#364745000000
1!
1%
#364750000000
0!
0%
#364755000000
1!
1%
#364760000000
0!
0%
#364765000000
1!
1%
#364770000000
0!
0%
#364775000000
1!
1%
#364780000000
0!
0%
#364785000000
1!
1%
#364790000000
0!
0%
#364795000000
1!
1%
#364800000000
0!
0%
#364805000000
1!
1%
#364810000000
0!
0%
#364815000000
1!
1%
#364820000000
0!
0%
#364825000000
1!
1%
#364830000000
0!
0%
#364835000000
1!
1%
#364840000000
0!
0%
#364845000000
1!
1%
#364850000000
0!
0%
#364855000000
1!
1%
#364860000000
0!
0%
#364865000000
1!
1%
#364870000000
0!
0%
#364875000000
1!
1%
#364880000000
0!
0%
#364885000000
1!
1%
#364890000000
0!
0%
#364895000000
1!
1%
#364900000000
0!
0%
#364905000000
1!
1%
#364910000000
0!
0%
#364915000000
1!
1%
#364920000000
0!
0%
#364925000000
1!
1%
#364930000000
0!
0%
#364935000000
1!
1%
#364940000000
0!
0%
#364945000000
1!
1%
#364950000000
0!
0%
#364955000000
1!
1%
#364960000000
0!
0%
#364965000000
1!
1%
#364970000000
0!
0%
#364975000000
1!
1%
#364980000000
0!
0%
#364985000000
1!
1%
#364990000000
0!
0%
#364995000000
1!
1%
#365000000000
0!
0%
#365005000000
1!
1%
#365010000000
0!
0%
#365015000000
1!
1%
#365020000000
0!
0%
#365025000000
1!
1%
#365030000000
0!
0%
#365035000000
1!
1%
#365040000000
0!
0%
#365045000000
1!
1%
#365050000000
0!
0%
#365055000000
1!
1%
#365060000000
0!
0%
#365065000000
1!
1%
#365070000000
0!
0%
#365075000000
1!
1%
#365080000000
0!
0%
#365085000000
1!
1%
#365090000000
0!
0%
#365095000000
1!
1%
#365100000000
0!
0%
#365105000000
1!
1%
#365110000000
0!
0%
#365115000000
1!
1%
#365120000000
0!
0%
#365125000000
1!
1%
#365130000000
0!
0%
#365135000000
1!
1%
#365140000000
0!
0%
#365145000000
1!
1%
#365150000000
0!
0%
#365155000000
1!
1%
#365160000000
0!
0%
#365165000000
1!
1%
#365170000000
0!
0%
#365175000000
1!
1%
#365180000000
0!
0%
#365185000000
1!
1%
#365190000000
0!
0%
#365195000000
1!
1%
#365200000000
0!
0%
#365205000000
1!
1%
#365210000000
0!
0%
#365215000000
1!
1%
#365220000000
0!
0%
#365225000000
1!
1%
#365230000000
0!
0%
#365235000000
1!
1%
#365240000000
0!
0%
#365245000000
1!
1%
#365250000000
0!
0%
#365255000000
1!
1%
#365260000000
0!
0%
#365265000000
1!
1%
#365270000000
0!
0%
#365275000000
1!
1%
#365280000000
0!
0%
#365285000000
1!
1%
#365290000000
0!
0%
#365295000000
1!
1%
#365300000000
0!
0%
#365305000000
1!
1%
#365310000000
0!
0%
#365315000000
1!
1%
#365320000000
0!
0%
#365325000000
1!
1%
#365330000000
0!
0%
#365335000000
1!
1%
#365340000000
0!
0%
#365345000000
1!
1%
#365350000000
0!
0%
#365355000000
1!
1%
#365360000000
0!
0%
#365365000000
1!
1%
#365370000000
0!
0%
#365375000000
1!
1%
#365380000000
0!
0%
#365385000000
1!
1%
#365390000000
0!
0%
#365395000000
1!
1%
#365400000000
0!
0%
#365405000000
1!
1%
#365410000000
0!
0%
#365415000000
1!
1%
#365420000000
0!
0%
#365425000000
1!
1%
#365430000000
0!
0%
#365435000000
1!
1%
#365440000000
0!
0%
#365445000000
1!
1%
#365450000000
0!
0%
#365455000000
1!
1%
#365460000000
0!
0%
#365465000000
1!
1%
#365470000000
0!
0%
#365475000000
1!
1%
#365480000000
0!
0%
#365485000000
1!
1%
#365490000000
0!
0%
#365495000000
1!
1%
#365500000000
0!
0%
#365505000000
1!
1%
#365510000000
0!
0%
#365515000000
1!
1%
#365520000000
0!
0%
#365525000000
1!
1%
#365530000000
0!
0%
#365535000000
1!
1%
#365540000000
0!
0%
#365545000000
1!
1%
#365550000000
0!
0%
#365555000000
1!
1%
#365560000000
0!
0%
#365565000000
1!
1%
#365570000000
0!
0%
#365575000000
1!
1%
#365580000000
0!
0%
#365585000000
1!
1%
#365590000000
0!
0%
#365595000000
1!
1%
#365600000000
0!
0%
#365605000000
1!
1%
#365610000000
0!
0%
#365615000000
1!
1%
#365620000000
0!
0%
#365625000000
1!
1%
#365630000000
0!
0%
#365635000000
1!
1%
#365640000000
0!
0%
#365645000000
1!
1%
#365650000000
0!
0%
#365655000000
1!
1%
#365660000000
0!
0%
#365665000000
1!
1%
#365670000000
0!
0%
#365675000000
1!
1%
#365680000000
0!
0%
#365685000000
1!
1%
#365690000000
0!
0%
#365695000000
1!
1%
#365700000000
0!
0%
#365705000000
1!
1%
#365710000000
0!
0%
#365715000000
1!
1%
#365720000000
0!
0%
#365725000000
1!
1%
#365730000000
0!
0%
#365735000000
1!
1%
#365740000000
0!
0%
#365745000000
1!
1%
#365750000000
0!
0%
#365755000000
1!
1%
#365760000000
0!
0%
#365765000000
1!
1%
#365770000000
0!
0%
#365775000000
1!
1%
#365780000000
0!
0%
#365785000000
1!
1%
#365790000000
0!
0%
#365795000000
1!
1%
#365800000000
0!
0%
#365805000000
1!
1%
#365810000000
0!
0%
#365815000000
1!
1%
#365820000000
0!
0%
#365825000000
1!
1%
#365830000000
0!
0%
#365835000000
1!
1%
#365840000000
0!
0%
#365845000000
1!
1%
#365850000000
0!
0%
#365855000000
1!
1%
#365860000000
0!
0%
#365865000000
1!
1%
#365870000000
0!
0%
#365875000000
1!
1%
#365880000000
0!
0%
#365885000000
1!
1%
#365890000000
0!
0%
#365895000000
1!
1%
#365900000000
0!
0%
#365905000000
1!
1%
#365910000000
0!
0%
#365915000000
1!
1%
#365920000000
0!
0%
#365925000000
1!
1%
#365930000000
0!
0%
#365935000000
1!
1%
#365940000000
0!
0%
#365945000000
1!
1%
#365950000000
0!
0%
#365955000000
1!
1%
#365960000000
0!
0%
#365965000000
1!
1%
#365970000000
0!
0%
#365975000000
1!
1%
#365980000000
0!
0%
#365985000000
1!
1%
#365990000000
0!
0%
#365995000000
1!
1%
#366000000000
0!
0%
#366005000000
1!
1%
#366010000000
0!
0%
#366015000000
1!
1%
#366020000000
0!
0%
#366025000000
1!
1%
#366030000000
0!
0%
#366035000000
1!
1%
#366040000000
0!
0%
#366045000000
1!
1%
#366050000000
0!
0%
#366055000000
1!
1%
#366060000000
0!
0%
#366065000000
1!
1%
#366070000000
0!
0%
#366075000000
1!
1%
#366080000000
0!
0%
#366085000000
1!
1%
#366090000000
0!
0%
#366095000000
1!
1%
#366100000000
0!
0%
#366105000000
1!
1%
#366110000000
0!
0%
#366115000000
1!
1%
#366120000000
0!
0%
#366125000000
1!
1%
#366130000000
0!
0%
#366135000000
1!
1%
#366140000000
0!
0%
#366145000000
1!
1%
#366150000000
0!
0%
#366155000000
1!
1%
#366160000000
0!
0%
#366165000000
1!
1%
#366170000000
0!
0%
#366175000000
1!
1%
#366180000000
0!
0%
#366185000000
1!
1%
#366190000000
0!
0%
#366195000000
1!
1%
#366200000000
0!
0%
#366205000000
1!
1%
#366210000000
0!
0%
#366215000000
1!
1%
#366220000000
0!
0%
#366225000000
1!
1%
#366230000000
0!
0%
#366235000000
1!
1%
#366240000000
0!
0%
#366245000000
1!
1%
#366250000000
0!
0%
#366255000000
1!
1%
#366260000000
0!
0%
#366265000000
1!
1%
#366270000000
0!
0%
#366275000000
1!
1%
#366280000000
0!
0%
#366285000000
1!
1%
#366290000000
0!
0%
#366295000000
1!
1%
#366300000000
0!
0%
#366305000000
1!
1%
#366310000000
0!
0%
#366315000000
1!
1%
#366320000000
0!
0%
#366325000000
1!
1%
#366330000000
0!
0%
#366335000000
1!
1%
#366340000000
0!
0%
#366345000000
1!
1%
#366350000000
0!
0%
#366355000000
1!
1%
#366360000000
0!
0%
#366365000000
1!
1%
#366370000000
0!
0%
#366375000000
1!
1%
#366380000000
0!
0%
#366385000000
1!
1%
#366390000000
0!
0%
#366395000000
1!
1%
#366400000000
0!
0%
#366405000000
1!
1%
#366410000000
0!
0%
#366415000000
1!
1%
#366420000000
0!
0%
#366425000000
1!
1%
#366430000000
0!
0%
#366435000000
1!
1%
#366440000000
0!
0%
#366445000000
1!
1%
#366450000000
0!
0%
#366455000000
1!
1%
#366460000000
0!
0%
#366465000000
1!
1%
#366470000000
0!
0%
#366475000000
1!
1%
#366480000000
0!
0%
#366485000000
1!
1%
#366490000000
0!
0%
#366495000000
1!
1%
#366500000000
0!
0%
#366505000000
1!
1%
#366510000000
0!
0%
#366515000000
1!
1%
#366520000000
0!
0%
#366525000000
1!
1%
#366530000000
0!
0%
#366535000000
1!
1%
#366540000000
0!
0%
#366545000000
1!
1%
#366550000000
0!
0%
#366555000000
1!
1%
#366560000000
0!
0%
#366565000000
1!
1%
#366570000000
0!
0%
#366575000000
1!
1%
#366580000000
0!
0%
#366585000000
1!
1%
#366590000000
0!
0%
#366595000000
1!
1%
#366600000000
0!
0%
#366605000000
1!
1%
#366610000000
0!
0%
#366615000000
1!
1%
#366620000000
0!
0%
#366625000000
1!
1%
#366630000000
0!
0%
#366635000000
1!
1%
#366640000000
0!
0%
#366645000000
1!
1%
#366650000000
0!
0%
#366655000000
1!
1%
#366660000000
0!
0%
#366665000000
1!
1%
#366670000000
0!
0%
#366675000000
1!
1%
#366680000000
0!
0%
#366685000000
1!
1%
#366690000000
0!
0%
#366695000000
1!
1%
#366700000000
0!
0%
#366705000000
1!
1%
#366710000000
0!
0%
#366715000000
1!
1%
#366720000000
0!
0%
#366725000000
1!
1%
#366730000000
0!
0%
#366735000000
1!
1%
#366740000000
0!
0%
#366745000000
1!
1%
#366750000000
0!
0%
#366755000000
1!
1%
#366760000000
0!
0%
#366765000000
1!
1%
#366770000000
0!
0%
#366775000000
1!
1%
#366780000000
0!
0%
#366785000000
1!
1%
#366790000000
0!
0%
#366795000000
1!
1%
#366800000000
0!
0%
#366805000000
1!
1%
#366810000000
0!
0%
#366815000000
1!
1%
#366820000000
0!
0%
#366825000000
1!
1%
#366830000000
0!
0%
#366835000000
1!
1%
#366840000000
0!
0%
#366845000000
1!
1%
#366850000000
0!
0%
#366855000000
1!
1%
#366860000000
0!
0%
#366865000000
1!
1%
#366870000000
0!
0%
#366875000000
1!
1%
#366880000000
0!
0%
#366885000000
1!
1%
#366890000000
0!
0%
#366895000000
1!
1%
#366900000000
0!
0%
#366905000000
1!
1%
#366910000000
0!
0%
#366915000000
1!
1%
#366920000000
0!
0%
#366925000000
1!
1%
#366930000000
0!
0%
#366935000000
1!
1%
#366940000000
0!
0%
#366945000000
1!
1%
#366950000000
0!
0%
#366955000000
1!
1%
#366960000000
0!
0%
#366965000000
1!
1%
#366970000000
0!
0%
#366975000000
1!
1%
#366980000000
0!
0%
#366985000000
1!
1%
#366990000000
0!
0%
#366995000000
1!
1%
#367000000000
0!
0%
#367005000000
1!
1%
#367010000000
0!
0%
#367015000000
1!
1%
#367020000000
0!
0%
#367025000000
1!
1%
#367030000000
0!
0%
#367035000000
1!
1%
#367040000000
0!
0%
#367045000000
1!
1%
#367050000000
0!
0%
#367055000000
1!
1%
#367060000000
0!
0%
#367065000000
1!
1%
#367070000000
0!
0%
#367075000000
1!
1%
#367080000000
0!
0%
#367085000000
1!
1%
#367090000000
0!
0%
#367095000000
1!
1%
#367100000000
0!
0%
#367105000000
1!
1%
#367110000000
0!
0%
#367115000000
1!
1%
#367120000000
0!
0%
#367125000000
1!
1%
#367130000000
0!
0%
#367135000000
1!
1%
#367140000000
0!
0%
#367145000000
1!
1%
#367150000000
0!
0%
#367155000000
1!
1%
#367160000000
0!
0%
#367165000000
1!
1%
#367170000000
0!
0%
#367175000000
1!
1%
#367180000000
0!
0%
#367185000000
1!
1%
#367190000000
0!
0%
#367195000000
1!
1%
#367200000000
0!
0%
#367205000000
1!
1%
#367210000000
0!
0%
#367215000000
1!
1%
#367220000000
0!
0%
#367225000000
1!
1%
#367230000000
0!
0%
#367235000000
1!
1%
#367240000000
0!
0%
#367245000000
1!
1%
#367250000000
0!
0%
#367255000000
1!
1%
#367260000000
0!
0%
#367265000000
1!
1%
#367270000000
0!
0%
#367275000000
1!
1%
#367280000000
0!
0%
#367285000000
1!
1%
#367290000000
0!
0%
#367295000000
1!
1%
#367300000000
0!
0%
#367305000000
1!
1%
#367310000000
0!
0%
#367315000000
1!
1%
#367320000000
0!
0%
#367325000000
1!
1%
#367330000000
0!
0%
#367335000000
1!
1%
#367340000000
0!
0%
#367345000000
1!
1%
#367350000000
0!
0%
#367355000000
1!
1%
#367360000000
0!
0%
#367365000000
1!
1%
#367370000000
0!
0%
#367375000000
1!
1%
#367380000000
0!
0%
#367385000000
1!
1%
#367390000000
0!
0%
#367395000000
1!
1%
#367400000000
0!
0%
#367405000000
1!
1%
#367410000000
0!
0%
#367415000000
1!
1%
#367420000000
0!
0%
#367425000000
1!
1%
#367430000000
0!
0%
#367435000000
1!
1%
#367440000000
0!
0%
#367445000000
1!
1%
#367450000000
0!
0%
#367455000000
1!
1%
#367460000000
0!
0%
#367465000000
1!
1%
#367470000000
0!
0%
#367475000000
1!
1%
#367480000000
0!
0%
#367485000000
1!
1%
#367490000000
0!
0%
#367495000000
1!
1%
#367500000000
0!
0%
#367505000000
1!
1%
#367510000000
0!
0%
#367515000000
1!
1%
#367520000000
0!
0%
#367525000000
1!
1%
#367530000000
0!
0%
#367535000000
1!
1%
#367540000000
0!
0%
#367545000000
1!
1%
#367550000000
0!
0%
#367555000000
1!
1%
#367560000000
0!
0%
#367565000000
1!
1%
#367570000000
0!
0%
#367575000000
1!
1%
#367580000000
0!
0%
#367585000000
1!
1%
#367590000000
0!
0%
#367595000000
1!
1%
#367600000000
0!
0%
#367605000000
1!
1%
#367610000000
0!
0%
#367615000000
1!
1%
#367620000000
0!
0%
#367625000000
1!
1%
#367630000000
0!
0%
#367635000000
1!
1%
#367640000000
0!
0%
#367645000000
1!
1%
#367650000000
0!
0%
#367655000000
1!
1%
#367660000000
0!
0%
#367665000000
1!
1%
#367670000000
0!
0%
#367675000000
1!
1%
#367680000000
0!
0%
#367685000000
1!
1%
#367690000000
0!
0%
#367695000000
1!
1%
#367700000000
0!
0%
#367705000000
1!
1%
#367710000000
0!
0%
#367715000000
1!
1%
#367720000000
0!
0%
#367725000000
1!
1%
#367730000000
0!
0%
#367735000000
1!
1%
#367740000000
0!
0%
#367745000000
1!
1%
#367750000000
0!
0%
#367755000000
1!
1%
#367760000000
0!
0%
#367765000000
1!
1%
#367770000000
0!
0%
#367775000000
1!
1%
#367780000000
0!
0%
#367785000000
1!
1%
#367790000000
0!
0%
#367795000000
1!
1%
#367800000000
0!
0%
#367805000000
1!
1%
#367810000000
0!
0%
#367815000000
1!
1%
#367820000000
0!
0%
#367825000000
1!
1%
#367830000000
0!
0%
#367835000000
1!
1%
#367840000000
0!
0%
#367845000000
1!
1%
#367850000000
0!
0%
#367855000000
1!
1%
#367860000000
0!
0%
#367865000000
1!
1%
#367870000000
0!
0%
#367875000000
1!
1%
#367880000000
0!
0%
#367885000000
1!
1%
#367890000000
0!
0%
#367895000000
1!
1%
#367900000000
0!
0%
#367905000000
1!
1%
#367910000000
0!
0%
#367915000000
1!
1%
#367920000000
0!
0%
#367925000000
1!
1%
#367930000000
0!
0%
#367935000000
1!
1%
#367940000000
0!
0%
#367945000000
1!
1%
#367950000000
0!
0%
#367955000000
1!
1%
#367960000000
0!
0%
#367965000000
1!
1%
#367970000000
0!
0%
#367975000000
1!
1%
#367980000000
0!
0%
#367985000000
1!
1%
#367990000000
0!
0%
#367995000000
1!
1%
#368000000000
0!
0%
#368005000000
1!
1%
#368010000000
0!
0%
#368015000000
1!
1%
#368020000000
0!
0%
#368025000000
1!
1%
#368030000000
0!
0%
#368035000000
1!
1%
#368040000000
0!
0%
#368045000000
1!
1%
#368050000000
0!
0%
#368055000000
1!
1%
#368060000000
0!
0%
#368065000000
1!
1%
#368070000000
0!
0%
#368075000000
1!
1%
#368080000000
0!
0%
#368085000000
1!
1%
#368090000000
0!
0%
#368095000000
1!
1%
#368100000000
0!
0%
#368105000000
1!
1%
#368110000000
0!
0%
#368115000000
1!
1%
#368120000000
0!
0%
#368125000000
1!
1%
#368130000000
0!
0%
#368135000000
1!
1%
#368140000000
0!
0%
#368145000000
1!
1%
#368150000000
0!
0%
#368155000000
1!
1%
#368160000000
0!
0%
#368165000000
1!
1%
#368170000000
0!
0%
#368175000000
1!
1%
#368180000000
0!
0%
#368185000000
1!
1%
#368190000000
0!
0%
#368195000000
1!
1%
#368200000000
0!
0%
#368205000000
1!
1%
#368210000000
0!
0%
#368215000000
1!
1%
#368220000000
0!
0%
#368225000000
1!
1%
#368230000000
0!
0%
#368235000000
1!
1%
#368240000000
0!
0%
#368245000000
1!
1%
#368250000000
0!
0%
#368255000000
1!
1%
#368260000000
0!
0%
#368265000000
1!
1%
#368270000000
0!
0%
#368275000000
1!
1%
#368280000000
0!
0%
#368285000000
1!
1%
#368290000000
0!
0%
#368295000000
1!
1%
#368300000000
0!
0%
#368305000000
1!
1%
#368310000000
0!
0%
#368315000000
1!
1%
#368320000000
0!
0%
#368325000000
1!
1%
#368330000000
0!
0%
#368335000000
1!
1%
#368340000000
0!
0%
#368345000000
1!
1%
#368350000000
0!
0%
#368355000000
1!
1%
#368360000000
0!
0%
#368365000000
1!
1%
#368370000000
0!
0%
#368375000000
1!
1%
#368380000000
0!
0%
#368385000000
1!
1%
#368390000000
0!
0%
#368395000000
1!
1%
#368400000000
0!
0%
#368405000000
1!
1%
#368410000000
0!
0%
#368415000000
1!
1%
#368420000000
0!
0%
#368425000000
1!
1%
#368430000000
0!
0%
#368435000000
1!
1%
#368440000000
0!
0%
#368445000000
1!
1%
#368450000000
0!
0%
#368455000000
1!
1%
#368460000000
0!
0%
#368465000000
1!
1%
#368470000000
0!
0%
#368475000000
1!
1%
#368480000000
0!
0%
#368485000000
1!
1%
#368490000000
0!
0%
#368495000000
1!
1%
#368500000000
0!
0%
#368505000000
1!
1%
#368510000000
0!
0%
#368515000000
1!
1%
#368520000000
0!
0%
#368525000000
1!
1%
#368530000000
0!
0%
#368535000000
1!
1%
#368540000000
0!
0%
#368545000000
1!
1%
#368550000000
0!
0%
#368555000000
1!
1%
#368560000000
0!
0%
#368565000000
1!
1%
#368570000000
0!
0%
#368575000000
1!
1%
#368580000000
0!
0%
#368585000000
1!
1%
#368590000000
0!
0%
#368595000000
1!
1%
#368600000000
0!
0%
#368605000000
1!
1%
#368610000000
0!
0%
#368615000000
1!
1%
#368620000000
0!
0%
#368625000000
1!
1%
#368630000000
0!
0%
#368635000000
1!
1%
#368640000000
0!
0%
#368645000000
1!
1%
#368650000000
0!
0%
#368655000000
1!
1%
#368660000000
0!
0%
#368665000000
1!
1%
#368670000000
0!
0%
#368675000000
1!
1%
#368680000000
0!
0%
#368685000000
1!
1%
#368690000000
0!
0%
#368695000000
1!
1%
#368700000000
0!
0%
#368705000000
1!
1%
#368710000000
0!
0%
#368715000000
1!
1%
#368720000000
0!
0%
#368725000000
1!
1%
#368730000000
0!
0%
#368735000000
1!
1%
#368740000000
0!
0%
#368745000000
1!
1%
#368750000000
0!
0%
#368755000000
1!
1%
#368760000000
0!
0%
#368765000000
1!
1%
#368770000000
0!
0%
#368775000000
1!
1%
#368780000000
0!
0%
#368785000000
1!
1%
#368790000000
0!
0%
#368795000000
1!
1%
#368800000000
0!
0%
#368805000000
1!
1%
#368810000000
0!
0%
#368815000000
1!
1%
#368820000000
0!
0%
#368825000000
1!
1%
#368830000000
0!
0%
#368835000000
1!
1%
#368840000000
0!
0%
#368845000000
1!
1%
#368850000000
0!
0%
#368855000000
1!
1%
#368860000000
0!
0%
#368865000000
1!
1%
#368870000000
0!
0%
#368875000000
1!
1%
#368880000000
0!
0%
#368885000000
1!
1%
#368890000000
0!
0%
#368895000000
1!
1%
#368900000000
0!
0%
#368905000000
1!
1%
#368910000000
0!
0%
#368915000000
1!
1%
#368920000000
0!
0%
#368925000000
1!
1%
#368930000000
0!
0%
#368935000000
1!
1%
#368940000000
0!
0%
#368945000000
1!
1%
#368950000000
0!
0%
#368955000000
1!
1%
#368960000000
0!
0%
#368965000000
1!
1%
#368970000000
0!
0%
#368975000000
1!
1%
#368980000000
0!
0%
#368985000000
1!
1%
#368990000000
0!
0%
#368995000000
1!
1%
#369000000000
0!
0%
#369005000000
1!
1%
#369010000000
0!
0%
#369015000000
1!
1%
#369020000000
0!
0%
#369025000000
1!
1%
#369030000000
0!
0%
#369035000000
1!
1%
#369040000000
0!
0%
#369045000000
1!
1%
#369050000000
0!
0%
#369055000000
1!
1%
#369060000000
0!
0%
#369065000000
1!
1%
#369070000000
0!
0%
#369075000000
1!
1%
#369080000000
0!
0%
#369085000000
1!
1%
#369090000000
0!
0%
#369095000000
1!
1%
#369100000000
0!
0%
#369105000000
1!
1%
#369110000000
0!
0%
#369115000000
1!
1%
#369120000000
0!
0%
#369125000000
1!
1%
#369130000000
0!
0%
#369135000000
1!
1%
#369140000000
0!
0%
#369145000000
1!
1%
#369150000000
0!
0%
#369155000000
1!
1%
#369160000000
0!
0%
#369165000000
1!
1%
#369170000000
0!
0%
#369175000000
1!
1%
#369180000000
0!
0%
#369185000000
1!
1%
#369190000000
0!
0%
#369195000000
1!
1%
#369200000000
0!
0%
#369205000000
1!
1%
#369210000000
0!
0%
#369215000000
1!
1%
#369220000000
0!
0%
#369225000000
1!
1%
#369230000000
0!
0%
#369235000000
1!
1%
#369240000000
0!
0%
#369245000000
1!
1%
#369250000000
0!
0%
#369255000000
1!
1%
#369260000000
0!
0%
#369265000000
1!
1%
#369270000000
0!
0%
#369275000000
1!
1%
#369280000000
0!
0%
#369285000000
1!
1%
#369290000000
0!
0%
#369295000000
1!
1%
#369300000000
0!
0%
#369305000000
1!
1%
#369310000000
0!
0%
#369315000000
1!
1%
#369320000000
0!
0%
#369325000000
1!
1%
#369330000000
0!
0%
#369335000000
1!
1%
#369340000000
0!
0%
#369345000000
1!
1%
#369350000000
0!
0%
#369355000000
1!
1%
#369360000000
0!
0%
#369365000000
1!
1%
#369370000000
0!
0%
#369375000000
1!
1%
#369380000000
0!
0%
#369385000000
1!
1%
#369390000000
0!
0%
#369395000000
1!
1%
#369400000000
0!
0%
#369405000000
1!
1%
#369410000000
0!
0%
#369415000000
1!
1%
#369420000000
0!
0%
#369425000000
1!
1%
#369430000000
0!
0%
#369435000000
1!
1%
#369440000000
0!
0%
#369445000000
1!
1%
#369450000000
0!
0%
#369455000000
1!
1%
#369460000000
0!
0%
#369465000000
1!
1%
#369470000000
0!
0%
#369475000000
1!
1%
#369480000000
0!
0%
#369485000000
1!
1%
#369490000000
0!
0%
#369495000000
1!
1%
#369500000000
0!
0%
#369505000000
1!
1%
#369510000000
0!
0%
#369515000000
1!
1%
#369520000000
0!
0%
#369525000000
1!
1%
#369530000000
0!
0%
#369535000000
1!
1%
#369540000000
0!
0%
#369545000000
1!
1%
#369550000000
0!
0%
#369555000000
1!
1%
#369560000000
0!
0%
#369565000000
1!
1%
#369570000000
0!
0%
#369575000000
1!
1%
#369580000000
0!
0%
#369585000000
1!
1%
#369590000000
0!
0%
#369595000000
1!
1%
#369600000000
0!
0%
#369605000000
1!
1%
#369610000000
0!
0%
#369615000000
1!
1%
#369620000000
0!
0%
#369625000000
1!
1%
#369630000000
0!
0%
#369635000000
1!
1%
#369640000000
0!
0%
#369645000000
1!
1%
#369650000000
0!
0%
#369655000000
1!
1%
#369660000000
0!
0%
#369665000000
1!
1%
#369670000000
0!
0%
#369675000000
1!
1%
#369680000000
0!
0%
#369685000000
1!
1%
#369690000000
0!
0%
#369695000000
1!
1%
#369700000000
0!
0%
#369705000000
1!
1%
#369710000000
0!
0%
#369715000000
1!
1%
#369720000000
0!
0%
#369725000000
1!
1%
#369730000000
0!
0%
#369735000000
1!
1%
#369740000000
0!
0%
#369745000000
1!
1%
#369750000000
0!
0%
#369755000000
1!
1%
#369760000000
0!
0%
#369765000000
1!
1%
#369770000000
0!
0%
#369775000000
1!
1%
#369780000000
0!
0%
#369785000000
1!
1%
#369790000000
0!
0%
#369795000000
1!
1%
#369800000000
0!
0%
#369805000000
1!
1%
#369810000000
0!
0%
#369815000000
1!
1%
#369820000000
0!
0%
#369825000000
1!
1%
#369830000000
0!
0%
#369835000000
1!
1%
#369840000000
0!
0%
#369845000000
1!
1%
#369850000000
0!
0%
#369855000000
1!
1%
#369860000000
0!
0%
#369865000000
1!
1%
#369870000000
0!
0%
#369875000000
1!
1%
#369880000000
0!
0%
#369885000000
1!
1%
#369890000000
0!
0%
#369895000000
1!
1%
#369900000000
0!
0%
#369905000000
1!
1%
#369910000000
0!
0%
#369915000000
1!
1%
#369920000000
0!
0%
#369925000000
1!
1%
#369930000000
0!
0%
#369935000000
1!
1%
#369940000000
0!
0%
#369945000000
1!
1%
#369950000000
0!
0%
#369955000000
1!
1%
#369960000000
0!
0%
#369965000000
1!
1%
#369970000000
0!
0%
#369975000000
1!
1%
#369980000000
0!
0%
#369985000000
1!
1%
#369990000000
0!
0%
#369995000000
1!
1%
#370000000000
0!
0%
#370005000000
1!
1%
#370010000000
0!
0%
#370015000000
1!
1%
#370020000000
0!
0%
#370025000000
1!
1%
#370030000000
0!
0%
#370035000000
1!
1%
#370040000000
0!
0%
#370045000000
1!
1%
#370050000000
0!
0%
#370055000000
1!
1%
#370060000000
0!
0%
#370065000000
1!
1%
#370070000000
0!
0%
#370075000000
1!
1%
#370080000000
0!
0%
#370085000000
1!
1%
#370090000000
0!
0%
#370095000000
1!
1%
#370100000000
0!
0%
#370105000000
1!
1%
#370110000000
0!
0%
#370115000000
1!
1%
#370120000000
0!
0%
#370125000000
1!
1%
#370130000000
0!
0%
#370135000000
1!
1%
#370140000000
0!
0%
#370145000000
1!
1%
#370150000000
0!
0%
#370155000000
1!
1%
#370160000000
0!
0%
#370165000000
1!
1%
#370170000000
0!
0%
#370175000000
1!
1%
#370180000000
0!
0%
#370185000000
1!
1%
#370190000000
0!
0%
#370195000000
1!
1%
#370200000000
0!
0%
#370205000000
1!
1%
#370210000000
0!
0%
#370215000000
1!
1%
#370220000000
0!
0%
#370225000000
1!
1%
#370230000000
0!
0%
#370235000000
1!
1%
#370240000000
0!
0%
#370245000000
1!
1%
#370250000000
0!
0%
#370255000000
1!
1%
#370260000000
0!
0%
#370265000000
1!
1%
#370270000000
0!
0%
#370275000000
1!
1%
#370280000000
0!
0%
#370285000000
1!
1%
#370290000000
0!
0%
#370295000000
1!
1%
#370300000000
0!
0%
#370305000000
1!
1%
#370310000000
0!
0%
#370315000000
1!
1%
#370320000000
0!
0%
#370325000000
1!
1%
#370330000000
0!
0%
#370335000000
1!
1%
#370340000000
0!
0%
#370345000000
1!
1%
#370350000000
0!
0%
#370355000000
1!
1%
#370360000000
0!
0%
#370365000000
1!
1%
#370370000000
0!
0%
#370375000000
1!
1%
#370380000000
0!
0%
#370385000000
1!
1%
#370390000000
0!
0%
#370395000000
1!
1%
#370400000000
0!
0%
#370405000000
1!
1%
#370410000000
0!
0%
#370415000000
1!
1%
#370420000000
0!
0%
#370425000000
1!
1%
#370430000000
0!
0%
#370435000000
1!
1%
#370440000000
0!
0%
#370445000000
1!
1%
#370450000000
0!
0%
#370455000000
1!
1%
#370460000000
0!
0%
#370465000000
1!
1%
#370470000000
0!
0%
#370475000000
1!
1%
#370480000000
0!
0%
#370485000000
1!
1%
#370490000000
0!
0%
#370495000000
1!
1%
#370500000000
0!
0%
#370505000000
1!
1%
#370510000000
0!
0%
#370515000000
1!
1%
#370520000000
0!
0%
#370525000000
1!
1%
#370530000000
0!
0%
#370535000000
1!
1%
#370540000000
0!
0%
#370545000000
1!
1%
#370550000000
0!
0%
#370555000000
1!
1%
#370560000000
0!
0%
#370565000000
1!
1%
#370570000000
0!
0%
#370575000000
1!
1%
#370580000000
0!
0%
#370585000000
1!
1%
#370590000000
0!
0%
#370595000000
1!
1%
#370600000000
0!
0%
#370605000000
1!
1%
#370610000000
0!
0%
#370615000000
1!
1%
#370620000000
0!
0%
#370625000000
1!
1%
#370630000000
0!
0%
#370635000000
1!
1%
#370640000000
0!
0%
#370645000000
1!
1%
#370650000000
0!
0%
#370655000000
1!
1%
#370660000000
0!
0%
#370665000000
1!
1%
#370670000000
0!
0%
#370675000000
1!
1%
#370680000000
0!
0%
#370685000000
1!
1%
#370690000000
0!
0%
#370695000000
1!
1%
#370700000000
0!
0%
#370705000000
1!
1%
#370710000000
0!
0%
#370715000000
1!
1%
#370720000000
0!
0%
#370725000000
1!
1%
#370730000000
0!
0%
#370735000000
1!
1%
#370740000000
0!
0%
#370745000000
1!
1%
#370750000000
0!
0%
#370755000000
1!
1%
#370760000000
0!
0%
#370765000000
1!
1%
#370770000000
0!
0%
#370775000000
1!
1%
#370780000000
0!
0%
#370785000000
1!
1%
#370790000000
0!
0%
#370795000000
1!
1%
#370800000000
0!
0%
#370805000000
1!
1%
#370810000000
0!
0%
#370815000000
1!
1%
#370820000000
0!
0%
#370825000000
1!
1%
#370830000000
0!
0%
#370835000000
1!
1%
#370840000000
0!
0%
#370845000000
1!
1%
#370850000000
0!
0%
#370855000000
1!
1%
#370860000000
0!
0%
#370865000000
1!
1%
#370870000000
0!
0%
#370875000000
1!
1%
#370880000000
0!
0%
#370885000000
1!
1%
#370890000000
0!
0%
#370895000000
1!
1%
#370900000000
0!
0%
#370905000000
1!
1%
#370910000000
0!
0%
#370915000000
1!
1%
#370920000000
0!
0%
#370925000000
1!
1%
#370930000000
0!
0%
#370935000000
1!
1%
#370940000000
0!
0%
#370945000000
1!
1%
#370950000000
0!
0%
#370955000000
1!
1%
#370960000000
0!
0%
#370965000000
1!
1%
#370970000000
0!
0%
#370975000000
1!
1%
#370980000000
0!
0%
#370985000000
1!
1%
#370990000000
0!
0%
#370995000000
1!
1%
#371000000000
0!
0%
#371005000000
1!
1%
#371010000000
0!
0%
#371015000000
1!
1%
#371020000000
0!
0%
#371025000000
1!
1%
#371030000000
0!
0%
#371035000000
1!
1%
#371040000000
0!
0%
#371045000000
1!
1%
#371050000000
0!
0%
#371055000000
1!
1%
#371060000000
0!
0%
#371065000000
1!
1%
#371070000000
0!
0%
#371075000000
1!
1%
#371080000000
0!
0%
#371085000000
1!
1%
#371090000000
0!
0%
#371095000000
1!
1%
#371100000000
0!
0%
#371105000000
1!
1%
#371110000000
0!
0%
#371115000000
1!
1%
#371120000000
0!
0%
#371125000000
1!
1%
#371130000000
0!
0%
#371135000000
1!
1%
#371140000000
0!
0%
#371145000000
1!
1%
#371150000000
0!
0%
#371155000000
1!
1%
#371160000000
0!
0%
#371165000000
1!
1%
#371170000000
0!
0%
#371175000000
1!
1%
#371180000000
0!
0%
#371185000000
1!
1%
#371190000000
0!
0%
#371195000000
1!
1%
#371200000000
0!
0%
#371205000000
1!
1%
#371210000000
0!
0%
#371215000000
1!
1%
#371220000000
0!
0%
#371225000000
1!
1%
#371230000000
0!
0%
#371235000000
1!
1%
#371240000000
0!
0%
#371245000000
1!
1%
#371250000000
0!
0%
#371255000000
1!
1%
#371260000000
0!
0%
#371265000000
1!
1%
#371270000000
0!
0%
#371275000000
1!
1%
#371280000000
0!
0%
#371285000000
1!
1%
#371290000000
0!
0%
#371295000000
1!
1%
#371300000000
0!
0%
#371305000000
1!
1%
#371310000000
0!
0%
#371315000000
1!
1%
#371320000000
0!
0%
#371325000000
1!
1%
#371330000000
0!
0%
#371335000000
1!
1%
#371340000000
0!
0%
#371345000000
1!
1%
#371350000000
0!
0%
#371355000000
1!
1%
#371360000000
0!
0%
#371365000000
1!
1%
#371370000000
0!
0%
#371375000000
1!
1%
#371380000000
0!
0%
#371385000000
1!
1%
#371390000000
0!
0%
#371395000000
1!
1%
#371400000000
0!
0%
#371405000000
1!
1%
#371410000000
0!
0%
#371415000000
1!
1%
#371420000000
0!
0%
#371425000000
1!
1%
#371430000000
0!
0%
#371435000000
1!
1%
#371440000000
0!
0%
#371445000000
1!
1%
#371450000000
0!
0%
#371455000000
1!
1%
#371460000000
0!
0%
#371465000000
1!
1%
#371470000000
0!
0%
#371475000000
1!
1%
#371480000000
0!
0%
#371485000000
1!
1%
#371490000000
0!
0%
#371495000000
1!
1%
#371500000000
0!
0%
#371505000000
1!
1%
#371510000000
0!
0%
#371515000000
1!
1%
#371520000000
0!
0%
#371525000000
1!
1%
#371530000000
0!
0%
#371535000000
1!
1%
#371540000000
0!
0%
#371545000000
1!
1%
#371550000000
0!
0%
#371555000000
1!
1%
#371560000000
0!
0%
#371565000000
1!
1%
#371570000000
0!
0%
#371575000000
1!
1%
#371580000000
0!
0%
#371585000000
1!
1%
#371590000000
0!
0%
#371595000000
1!
1%
#371600000000
0!
0%
#371605000000
1!
1%
#371610000000
0!
0%
#371615000000
1!
1%
#371620000000
0!
0%
#371625000000
1!
1%
#371630000000
0!
0%
#371635000000
1!
1%
#371640000000
0!
0%
#371645000000
1!
1%
#371650000000
0!
0%
#371655000000
1!
1%
#371660000000
0!
0%
#371665000000
1!
1%
#371670000000
0!
0%
#371675000000
1!
1%
#371680000000
0!
0%
#371685000000
1!
1%
#371690000000
0!
0%
#371695000000
1!
1%
#371700000000
0!
0%
#371705000000
1!
1%
#371710000000
0!
0%
#371715000000
1!
1%
#371720000000
0!
0%
#371725000000
1!
1%
#371730000000
0!
0%
#371735000000
1!
1%
#371740000000
0!
0%
#371745000000
1!
1%
#371750000000
0!
0%
#371755000000
1!
1%
#371760000000
0!
0%
#371765000000
1!
1%
#371770000000
0!
0%
#371775000000
1!
1%
#371780000000
0!
0%
#371785000000
1!
1%
#371790000000
0!
0%
#371795000000
1!
1%
#371800000000
0!
0%
#371805000000
1!
1%
#371810000000
0!
0%
#371815000000
1!
1%
#371820000000
0!
0%
#371825000000
1!
1%
#371830000000
0!
0%
#371835000000
1!
1%
#371840000000
0!
0%
#371845000000
1!
1%
#371850000000
0!
0%
#371855000000
1!
1%
#371860000000
0!
0%
#371865000000
1!
1%
#371870000000
0!
0%
#371875000000
1!
1%
#371880000000
0!
0%
#371885000000
1!
1%
#371890000000
0!
0%
#371895000000
1!
1%
#371900000000
0!
0%
#371905000000
1!
1%
#371910000000
0!
0%
#371915000000
1!
1%
#371920000000
0!
0%
#371925000000
1!
1%
#371930000000
0!
0%
#371935000000
1!
1%
#371940000000
0!
0%
#371945000000
1!
1%
#371950000000
0!
0%
#371955000000
1!
1%
#371960000000
0!
0%
#371965000000
1!
1%
#371970000000
0!
0%
#371975000000
1!
1%
#371980000000
0!
0%
#371985000000
1!
1%
#371990000000
0!
0%
#371995000000
1!
1%
#372000000000
0!
0%
#372005000000
1!
1%
#372010000000
0!
0%
#372015000000
1!
1%
#372020000000
0!
0%
#372025000000
1!
1%
#372030000000
0!
0%
#372035000000
1!
1%
#372040000000
0!
0%
#372045000000
1!
1%
#372050000000
0!
0%
#372055000000
1!
1%
#372060000000
0!
0%
#372065000000
1!
1%
#372070000000
0!
0%
#372075000000
1!
1%
#372080000000
0!
0%
#372085000000
1!
1%
#372090000000
0!
0%
#372095000000
1!
1%
#372100000000
0!
0%
#372105000000
1!
1%
#372110000000
0!
0%
#372115000000
1!
1%
#372120000000
0!
0%
#372125000000
1!
1%
#372130000000
0!
0%
#372135000000
1!
1%
#372140000000
0!
0%
#372145000000
1!
1%
#372150000000
0!
0%
#372155000000
1!
1%
#372160000000
0!
0%
#372165000000
1!
1%
#372170000000
0!
0%
#372175000000
1!
1%
#372180000000
0!
0%
#372185000000
1!
1%
#372190000000
0!
0%
#372195000000
1!
1%
#372200000000
0!
0%
#372205000000
1!
1%
#372210000000
0!
0%
#372215000000
1!
1%
#372220000000
0!
0%
#372225000000
1!
1%
#372230000000
0!
0%
#372235000000
1!
1%
#372240000000
0!
0%
#372245000000
1!
1%
#372250000000
0!
0%
#372255000000
1!
1%
#372260000000
0!
0%
#372265000000
1!
1%
#372270000000
0!
0%
#372275000000
1!
1%
#372280000000
0!
0%
#372285000000
1!
1%
#372290000000
0!
0%
#372295000000
1!
1%
#372300000000
0!
0%
#372305000000
1!
1%
#372310000000
0!
0%
#372315000000
1!
1%
#372320000000
0!
0%
#372325000000
1!
1%
#372330000000
0!
0%
#372335000000
1!
1%
#372340000000
0!
0%
#372345000000
1!
1%
#372350000000
0!
0%
#372355000000
1!
1%
#372360000000
0!
0%
#372365000000
1!
1%
#372370000000
0!
0%
#372375000000
1!
1%
#372380000000
0!
0%
#372385000000
1!
1%
#372390000000
0!
0%
#372395000000
1!
1%
#372400000000
0!
0%
#372405000000
1!
1%
#372410000000
0!
0%
#372415000000
1!
1%
#372420000000
0!
0%
#372425000000
1!
1%
#372430000000
0!
0%
#372435000000
1!
1%
#372440000000
0!
0%
#372445000000
1!
1%
#372450000000
0!
0%
#372455000000
1!
1%
#372460000000
0!
0%
#372465000000
1!
1%
#372470000000
0!
0%
#372475000000
1!
1%
#372480000000
0!
0%
#372485000000
1!
1%
#372490000000
0!
0%
#372495000000
1!
1%
#372500000000
0!
0%
#372505000000
1!
1%
#372510000000
0!
0%
#372515000000
1!
1%
#372520000000
0!
0%
#372525000000
1!
1%
#372530000000
0!
0%
#372535000000
1!
1%
#372540000000
0!
0%
#372545000000
1!
1%
#372550000000
0!
0%
#372555000000
1!
1%
#372560000000
0!
0%
#372565000000
1!
1%
#372570000000
0!
0%
#372575000000
1!
1%
#372580000000
0!
0%
#372585000000
1!
1%
#372590000000
0!
0%
#372595000000
1!
1%
#372600000000
0!
0%
#372605000000
1!
1%
#372610000000
0!
0%
#372615000000
1!
1%
#372620000000
0!
0%
#372625000000
1!
1%
#372630000000
0!
0%
#372635000000
1!
1%
#372640000000
0!
0%
#372645000000
1!
1%
#372650000000
0!
0%
#372655000000
1!
1%
#372660000000
0!
0%
#372665000000
1!
1%
#372670000000
0!
0%
#372675000000
1!
1%
#372680000000
0!
0%
#372685000000
1!
1%
#372690000000
0!
0%
#372695000000
1!
1%
#372700000000
0!
0%
#372705000000
1!
1%
#372710000000
0!
0%
#372715000000
1!
1%
#372720000000
0!
0%
#372725000000
1!
1%
#372730000000
0!
0%
#372735000000
1!
1%
#372740000000
0!
0%
#372745000000
1!
1%
#372750000000
0!
0%
#372755000000
1!
1%
#372760000000
0!
0%
#372765000000
1!
1%
#372770000000
0!
0%
#372775000000
1!
1%
#372780000000
0!
0%
#372785000000
1!
1%
#372790000000
0!
0%
#372795000000
1!
1%
#372800000000
0!
0%
#372805000000
1!
1%
#372810000000
0!
0%
#372815000000
1!
1%
#372820000000
0!
0%
#372825000000
1!
1%
#372830000000
0!
0%
#372835000000
1!
1%
#372840000000
0!
0%
#372845000000
1!
1%
#372850000000
0!
0%
#372855000000
1!
1%
#372860000000
0!
0%
#372865000000
1!
1%
#372870000000
0!
0%
#372875000000
1!
1%
#372880000000
0!
0%
#372885000000
1!
1%
#372890000000
0!
0%
#372895000000
1!
1%
#372900000000
0!
0%
#372905000000
1!
1%
#372910000000
0!
0%
#372915000000
1!
1%
#372920000000
0!
0%
#372925000000
1!
1%
#372930000000
0!
0%
#372935000000
1!
1%
#372940000000
0!
0%
#372945000000
1!
1%
#372950000000
0!
0%
#372955000000
1!
1%
#372960000000
0!
0%
#372965000000
1!
1%
#372970000000
0!
0%
#372975000000
1!
1%
#372980000000
0!
0%
#372985000000
1!
1%
#372990000000
0!
0%
#372995000000
1!
1%
#373000000000
0!
0%
#373005000000
1!
1%
#373010000000
0!
0%
#373015000000
1!
1%
#373020000000
0!
0%
#373025000000
1!
1%
#373030000000
0!
0%
#373035000000
1!
1%
#373040000000
0!
0%
#373045000000
1!
1%
#373050000000
0!
0%
#373055000000
1!
1%
#373060000000
0!
0%
#373065000000
1!
1%
#373070000000
0!
0%
#373075000000
1!
1%
#373080000000
0!
0%
#373085000000
1!
1%
#373090000000
0!
0%
#373095000000
1!
1%
#373100000000
0!
0%
#373105000000
1!
1%
#373110000000
0!
0%
#373115000000
1!
1%
#373120000000
0!
0%
#373125000000
1!
1%
#373130000000
0!
0%
#373135000000
1!
1%
#373140000000
0!
0%
#373145000000
1!
1%
#373150000000
0!
0%
#373155000000
1!
1%
#373160000000
0!
0%
#373165000000
1!
1%
#373170000000
0!
0%
#373175000000
1!
1%
#373180000000
0!
0%
#373185000000
1!
1%
#373190000000
0!
0%
#373195000000
1!
1%
#373200000000
0!
0%
#373205000000
1!
1%
#373210000000
0!
0%
#373215000000
1!
1%
#373220000000
0!
0%
#373225000000
1!
1%
#373230000000
0!
0%
#373235000000
1!
1%
#373240000000
0!
0%
#373245000000
1!
1%
#373250000000
0!
0%
#373255000000
1!
1%
#373260000000
0!
0%
#373265000000
1!
1%
#373270000000
0!
0%
#373275000000
1!
1%
#373280000000
0!
0%
#373285000000
1!
1%
#373290000000
0!
0%
#373295000000
1!
1%
#373300000000
0!
0%
#373305000000
1!
1%
#373310000000
0!
0%
#373315000000
1!
1%
#373320000000
0!
0%
#373325000000
1!
1%
#373330000000
0!
0%
#373335000000
1!
1%
#373340000000
0!
0%
#373345000000
1!
1%
#373350000000
0!
0%
#373355000000
1!
1%
#373360000000
0!
0%
#373365000000
1!
1%
#373370000000
0!
0%
#373375000000
1!
1%
#373380000000
0!
0%
#373385000000
1!
1%
#373390000000
0!
0%
#373395000000
1!
1%
#373400000000
0!
0%
#373405000000
1!
1%
#373410000000
0!
0%
#373415000000
1!
1%
#373420000000
0!
0%
#373425000000
1!
1%
#373430000000
0!
0%
#373435000000
1!
1%
#373440000000
0!
0%
#373445000000
1!
1%
#373450000000
0!
0%
#373455000000
1!
1%
#373460000000
0!
0%
#373465000000
1!
1%
#373470000000
0!
0%
#373475000000
1!
1%
#373480000000
0!
0%
#373485000000
1!
1%
#373490000000
0!
0%
#373495000000
1!
1%
#373500000000
0!
0%
#373505000000
1!
1%
#373510000000
0!
0%
#373515000000
1!
1%
#373520000000
0!
0%
#373525000000
1!
1%
#373530000000
0!
0%
#373535000000
1!
1%
#373540000000
0!
0%
#373545000000
1!
1%
#373550000000
0!
0%
#373555000000
1!
1%
#373560000000
0!
0%
#373565000000
1!
1%
#373570000000
0!
0%
#373575000000
1!
1%
#373580000000
0!
0%
#373585000000
1!
1%
#373590000000
0!
0%
#373595000000
1!
1%
#373600000000
0!
0%
#373605000000
1!
1%
#373610000000
0!
0%
#373615000000
1!
1%
#373620000000
0!
0%
#373625000000
1!
1%
#373630000000
0!
0%
#373635000000
1!
1%
#373640000000
0!
0%
#373645000000
1!
1%
#373650000000
0!
0%
#373655000000
1!
1%
#373660000000
0!
0%
#373665000000
1!
1%
#373670000000
0!
0%
#373675000000
1!
1%
#373680000000
0!
0%
#373685000000
1!
1%
#373690000000
0!
0%
#373695000000
1!
1%
#373700000000
0!
0%
#373705000000
1!
1%
#373710000000
0!
0%
#373715000000
1!
1%
#373720000000
0!
0%
#373725000000
1!
1%
#373730000000
0!
0%
#373735000000
1!
1%
#373740000000
0!
0%
#373745000000
1!
1%
#373750000000
0!
0%
#373755000000
1!
1%
#373760000000
0!
0%
#373765000000
1!
1%
#373770000000
0!
0%
#373775000000
1!
1%
#373780000000
0!
0%
#373785000000
1!
1%
#373790000000
0!
0%
#373795000000
1!
1%
#373800000000
0!
0%
#373805000000
1!
1%
#373810000000
0!
0%
#373815000000
1!
1%
#373820000000
0!
0%
#373825000000
1!
1%
#373830000000
0!
0%
#373835000000
1!
1%
#373840000000
0!
0%
#373845000000
1!
1%
#373850000000
0!
0%
#373855000000
1!
1%
#373860000000
0!
0%
#373865000000
1!
1%
#373870000000
0!
0%
#373875000000
1!
1%
#373880000000
0!
0%
#373885000000
1!
1%
#373890000000
0!
0%
#373895000000
1!
1%
#373900000000
0!
0%
#373905000000
1!
1%
#373910000000
0!
0%
#373915000000
1!
1%
#373920000000
0!
0%
#373925000000
1!
1%
#373930000000
0!
0%
#373935000000
1!
1%
#373940000000
0!
0%
#373945000000
1!
1%
#373950000000
0!
0%
#373955000000
1!
1%
#373960000000
0!
0%
#373965000000
1!
1%
#373970000000
0!
0%
#373975000000
1!
1%
#373980000000
0!
0%
#373985000000
1!
1%
#373990000000
0!
0%
#373995000000
1!
1%
#374000000000
0!
0%
#374005000000
1!
1%
#374010000000
0!
0%
#374015000000
1!
1%
#374020000000
0!
0%
#374025000000
1!
1%
#374030000000
0!
0%
#374035000000
1!
1%
#374040000000
0!
0%
#374045000000
1!
1%
#374050000000
0!
0%
#374055000000
1!
1%
#374060000000
0!
0%
#374065000000
1!
1%
#374070000000
0!
0%
#374075000000
1!
1%
#374080000000
0!
0%
#374085000000
1!
1%
#374090000000
0!
0%
#374095000000
1!
1%
#374100000000
0!
0%
#374105000000
1!
1%
#374110000000
0!
0%
#374115000000
1!
1%
#374120000000
0!
0%
#374125000000
1!
1%
#374130000000
0!
0%
#374135000000
1!
1%
#374140000000
0!
0%
#374145000000
1!
1%
#374150000000
0!
0%
#374155000000
1!
1%
#374160000000
0!
0%
#374165000000
1!
1%
#374170000000
0!
0%
#374175000000
1!
1%
#374180000000
0!
0%
#374185000000
1!
1%
#374190000000
0!
0%
#374195000000
1!
1%
#374200000000
0!
0%
#374205000000
1!
1%
#374210000000
0!
0%
#374215000000
1!
1%
#374220000000
0!
0%
#374225000000
1!
1%
#374230000000
0!
0%
#374235000000
1!
1%
#374240000000
0!
0%
#374245000000
1!
1%
#374250000000
0!
0%
#374255000000
1!
1%
#374260000000
0!
0%
#374265000000
1!
1%
#374270000000
0!
0%
#374275000000
1!
1%
#374280000000
0!
0%
#374285000000
1!
1%
#374290000000
0!
0%
#374295000000
1!
1%
#374300000000
0!
0%
#374305000000
1!
1%
#374310000000
0!
0%
#374315000000
1!
1%
#374320000000
0!
0%
#374325000000
1!
1%
#374330000000
0!
0%
#374335000000
1!
1%
#374340000000
0!
0%
#374345000000
1!
1%
#374350000000
0!
0%
#374355000000
1!
1%
#374360000000
0!
0%
#374365000000
1!
1%
#374370000000
0!
0%
#374375000000
1!
1%
#374380000000
0!
0%
#374385000000
1!
1%
#374390000000
0!
0%
#374395000000
1!
1%
#374400000000
0!
0%
#374405000000
1!
1%
#374410000000
0!
0%
#374415000000
1!
1%
#374420000000
0!
0%
#374425000000
1!
1%
#374430000000
0!
0%
#374435000000
1!
1%
#374440000000
0!
0%
#374445000000
1!
1%
#374450000000
0!
0%
#374455000000
1!
1%
#374460000000
0!
0%
#374465000000
1!
1%
#374470000000
0!
0%
#374475000000
1!
1%
#374480000000
0!
0%
#374485000000
1!
1%
#374490000000
0!
0%
#374495000000
1!
1%
#374500000000
0!
0%
#374505000000
1!
1%
#374510000000
0!
0%
#374515000000
1!
1%
#374520000000
0!
0%
#374525000000
1!
1%
#374530000000
0!
0%
#374535000000
1!
1%
#374540000000
0!
0%
#374545000000
1!
1%
#374550000000
0!
0%
#374555000000
1!
1%
#374560000000
0!
0%
#374565000000
1!
1%
#374570000000
0!
0%
#374575000000
1!
1%
#374580000000
0!
0%
#374585000000
1!
1%
#374590000000
0!
0%
#374595000000
1!
1%
#374600000000
0!
0%
#374605000000
1!
1%
#374610000000
0!
0%
#374615000000
1!
1%
#374620000000
0!
0%
#374625000000
1!
1%
#374630000000
0!
0%
#374635000000
1!
1%
#374640000000
0!
0%
#374645000000
1!
1%
#374650000000
0!
0%
#374655000000
1!
1%
#374660000000
0!
0%
#374665000000
1!
1%
#374670000000
0!
0%
#374675000000
1!
1%
#374680000000
0!
0%
#374685000000
1!
1%
#374690000000
0!
0%
#374695000000
1!
1%
#374700000000
0!
0%
#374705000000
1!
1%
#374710000000
0!
0%
#374715000000
1!
1%
#374720000000
0!
0%
#374725000000
1!
1%
#374730000000
0!
0%
#374735000000
1!
1%
#374740000000
0!
0%
#374745000000
1!
1%
#374750000000
0!
0%
#374755000000
1!
1%
#374760000000
0!
0%
#374765000000
1!
1%
#374770000000
0!
0%
#374775000000
1!
1%
#374780000000
0!
0%
#374785000000
1!
1%
#374790000000
0!
0%
#374795000000
1!
1%
#374800000000
0!
0%
#374805000000
1!
1%
#374810000000
0!
0%
#374815000000
1!
1%
#374820000000
0!
0%
#374825000000
1!
1%
#374830000000
0!
0%
#374835000000
1!
1%
#374840000000
0!
0%
#374845000000
1!
1%
#374850000000
0!
0%
#374855000000
1!
1%
#374860000000
0!
0%
#374865000000
1!
1%
#374870000000
0!
0%
#374875000000
1!
1%
#374880000000
0!
0%
#374885000000
1!
1%
#374890000000
0!
0%
#374895000000
1!
1%
#374900000000
0!
0%
#374905000000
1!
1%
#374910000000
0!
0%
#374915000000
1!
1%
#374920000000
0!
0%
#374925000000
1!
1%
#374930000000
0!
0%
#374935000000
1!
1%
#374940000000
0!
0%
#374945000000
1!
1%
#374950000000
0!
0%
#374955000000
1!
1%
#374960000000
0!
0%
#374965000000
1!
1%
#374970000000
0!
0%
#374975000000
1!
1%
#374980000000
0!
0%
#374985000000
1!
1%
#374990000000
0!
0%
#374995000000
1!
1%
#375000000000
0!
0%
#375005000000
1!
1%
#375010000000
0!
0%
#375015000000
1!
1%
#375020000000
0!
0%
#375025000000
1!
1%
#375030000000
0!
0%
#375035000000
1!
1%
#375040000000
0!
0%
#375045000000
1!
1%
#375050000000
0!
0%
#375055000000
1!
1%
#375060000000
0!
0%
#375065000000
1!
1%
#375070000000
0!
0%
#375075000000
1!
1%
#375080000000
0!
0%
#375085000000
1!
1%
#375090000000
0!
0%
#375095000000
1!
1%
#375100000000
0!
0%
#375105000000
1!
1%
#375110000000
0!
0%
#375115000000
1!
1%
#375120000000
0!
0%
#375125000000
1!
1%
#375130000000
0!
0%
#375135000000
1!
1%
#375140000000
0!
0%
#375145000000
1!
1%
#375150000000
0!
0%
#375155000000
1!
1%
#375160000000
0!
0%
#375165000000
1!
1%
#375170000000
0!
0%
#375175000000
1!
1%
#375180000000
0!
0%
#375185000000
1!
1%
#375190000000
0!
0%
#375195000000
1!
1%
#375200000000
0!
0%
#375205000000
1!
1%
#375210000000
0!
0%
#375215000000
1!
1%
#375220000000
0!
0%
#375225000000
1!
1%
#375230000000
0!
0%
#375235000000
1!
1%
#375240000000
0!
0%
#375245000000
1!
1%
#375250000000
0!
0%
#375255000000
1!
1%
#375260000000
0!
0%
#375265000000
1!
1%
#375270000000
0!
0%
#375275000000
1!
1%
#375280000000
0!
0%
#375285000000
1!
1%
#375290000000
0!
0%
#375295000000
1!
1%
#375300000000
0!
0%
#375305000000
1!
1%
#375310000000
0!
0%
#375315000000
1!
1%
#375320000000
0!
0%
#375325000000
1!
1%
#375330000000
0!
0%
#375335000000
1!
1%
#375340000000
0!
0%
#375345000000
1!
1%
#375350000000
0!
0%
#375355000000
1!
1%
#375360000000
0!
0%
#375365000000
1!
1%
#375370000000
0!
0%
#375375000000
1!
1%
#375380000000
0!
0%
#375385000000
1!
1%
#375390000000
0!
0%
#375395000000
1!
1%
#375400000000
0!
0%
#375405000000
1!
1%
#375410000000
0!
0%
#375415000000
1!
1%
#375420000000
0!
0%
#375425000000
1!
1%
#375430000000
0!
0%
#375435000000
1!
1%
#375440000000
0!
0%
#375445000000
1!
1%
#375450000000
0!
0%
#375455000000
1!
1%
#375460000000
0!
0%
#375465000000
1!
1%
#375470000000
0!
0%
#375475000000
1!
1%
#375480000000
0!
0%
#375485000000
1!
1%
#375490000000
0!
0%
#375495000000
1!
1%
#375500000000
0!
0%
#375505000000
1!
1%
#375510000000
0!
0%
#375515000000
1!
1%
#375520000000
0!
0%
#375525000000
1!
1%
#375530000000
0!
0%
#375535000000
1!
1%
#375540000000
0!
0%
#375545000000
1!
1%
#375550000000
0!
0%
#375555000000
1!
1%
#375560000000
0!
0%
#375565000000
1!
1%
#375570000000
0!
0%
#375575000000
1!
1%
#375580000000
0!
0%
#375585000000
1!
1%
#375590000000
0!
0%
#375595000000
1!
1%
#375600000000
0!
0%
#375605000000
1!
1%
#375610000000
0!
0%
#375615000000
1!
1%
#375620000000
0!
0%
#375625000000
1!
1%
#375630000000
0!
0%
#375635000000
1!
1%
#375640000000
0!
0%
#375645000000
1!
1%
#375650000000
0!
0%
#375655000000
1!
1%
#375660000000
0!
0%
#375665000000
1!
1%
#375670000000
0!
0%
#375675000000
1!
1%
#375680000000
0!
0%
#375685000000
1!
1%
#375690000000
0!
0%
#375695000000
1!
1%
#375700000000
0!
0%
#375705000000
1!
1%
#375710000000
0!
0%
#375715000000
1!
1%
#375720000000
0!
0%
#375725000000
1!
1%
#375730000000
0!
0%
#375735000000
1!
1%
#375740000000
0!
0%
#375745000000
1!
1%
#375750000000
0!
0%
#375755000000
1!
1%
#375760000000
0!
0%
#375765000000
1!
1%
#375770000000
0!
0%
#375775000000
1!
1%
#375780000000
0!
0%
#375785000000
1!
1%
#375790000000
0!
0%
#375795000000
1!
1%
#375800000000
0!
0%
#375805000000
1!
1%
#375810000000
0!
0%
#375815000000
1!
1%
#375820000000
0!
0%
#375825000000
1!
1%
#375830000000
0!
0%
#375835000000
1!
1%
#375840000000
0!
0%
#375845000000
1!
1%
#375850000000
0!
0%
#375855000000
1!
1%
#375860000000
0!
0%
#375865000000
1!
1%
#375870000000
0!
0%
#375875000000
1!
1%
#375880000000
0!
0%
#375885000000
1!
1%
#375890000000
0!
0%
#375895000000
1!
1%
#375900000000
0!
0%
#375905000000
1!
1%
#375910000000
0!
0%
#375915000000
1!
1%
#375920000000
0!
0%
#375925000000
1!
1%
#375930000000
0!
0%
#375935000000
1!
1%
#375940000000
0!
0%
#375945000000
1!
1%
#375950000000
0!
0%
#375955000000
1!
1%
#375960000000
0!
0%
#375965000000
1!
1%
#375970000000
0!
0%
#375975000000
1!
1%
#375980000000
0!
0%
#375985000000
1!
1%
#375990000000
0!
0%
#375995000000
1!
1%
#376000000000
0!
0%
#376005000000
1!
1%
#376010000000
0!
0%
#376015000000
1!
1%
#376020000000
0!
0%
#376025000000
1!
1%
#376030000000
0!
0%
#376035000000
1!
1%
#376040000000
0!
0%
#376045000000
1!
1%
#376050000000
0!
0%
#376055000000
1!
1%
#376060000000
0!
0%
#376065000000
1!
1%
#376070000000
0!
0%
#376075000000
1!
1%
#376080000000
0!
0%
#376085000000
1!
1%
#376090000000
0!
0%
#376095000000
1!
1%
#376100000000
0!
0%
#376105000000
1!
1%
#376110000000
0!
0%
#376115000000
1!
1%
#376120000000
0!
0%
#376125000000
1!
1%
#376130000000
0!
0%
#376135000000
1!
1%
#376140000000
0!
0%
#376145000000
1!
1%
#376150000000
0!
0%
#376155000000
1!
1%
#376160000000
0!
0%
#376165000000
1!
1%
#376170000000
0!
0%
#376175000000
1!
1%
#376180000000
0!
0%
#376185000000
1!
1%
#376190000000
0!
0%
#376195000000
1!
1%
#376200000000
0!
0%
#376205000000
1!
1%
#376210000000
0!
0%
#376215000000
1!
1%
#376220000000
0!
0%
#376225000000
1!
1%
#376230000000
0!
0%
#376235000000
1!
1%
#376240000000
0!
0%
#376245000000
1!
1%
#376250000000
0!
0%
#376255000000
1!
1%
#376260000000
0!
0%
#376265000000
1!
1%
#376270000000
0!
0%
#376275000000
1!
1%
#376280000000
0!
0%
#376285000000
1!
1%
#376290000000
0!
0%
#376295000000
1!
1%
#376300000000
0!
0%
#376305000000
1!
1%
#376310000000
0!
0%
#376315000000
1!
1%
#376320000000
0!
0%
#376325000000
1!
1%
#376330000000
0!
0%
#376335000000
1!
1%
#376340000000
0!
0%
#376345000000
1!
1%
#376350000000
0!
0%
#376355000000
1!
1%
#376360000000
0!
0%
#376365000000
1!
1%
#376370000000
0!
0%
#376375000000
1!
1%
#376380000000
0!
0%
#376385000000
1!
1%
#376390000000
0!
0%
#376395000000
1!
1%
#376400000000
0!
0%
#376405000000
1!
1%
#376410000000
0!
0%
#376415000000
1!
1%
#376420000000
0!
0%
#376425000000
1!
1%
#376430000000
0!
0%
#376435000000
1!
1%
#376440000000
0!
0%
#376445000000
1!
1%
#376450000000
0!
0%
#376455000000
1!
1%
#376460000000
0!
0%
#376465000000
1!
1%
#376470000000
0!
0%
#376475000000
1!
1%
#376480000000
0!
0%
#376485000000
1!
1%
#376490000000
0!
0%
#376495000000
1!
1%
#376500000000
0!
0%
#376505000000
1!
1%
#376510000000
0!
0%
#376515000000
1!
1%
#376520000000
0!
0%
#376525000000
1!
1%
#376530000000
0!
0%
#376535000000
1!
1%
#376540000000
0!
0%
#376545000000
1!
1%
#376550000000
0!
0%
#376555000000
1!
1%
#376560000000
0!
0%
#376565000000
1!
1%
#376570000000
0!
0%
#376575000000
1!
1%
#376580000000
0!
0%
#376585000000
1!
1%
#376590000000
0!
0%
#376595000000
1!
1%
#376600000000
0!
0%
#376605000000
1!
1%
#376610000000
0!
0%
#376615000000
1!
1%
#376620000000
0!
0%
#376625000000
1!
1%
#376630000000
0!
0%
#376635000000
1!
1%
#376640000000
0!
0%
#376645000000
1!
1%
#376650000000
0!
0%
#376655000000
1!
1%
#376660000000
0!
0%
#376665000000
1!
1%
#376670000000
0!
0%
#376675000000
1!
1%
#376680000000
0!
0%
#376685000000
1!
1%
#376690000000
0!
0%
#376695000000
1!
1%
#376700000000
0!
0%
#376705000000
1!
1%
#376710000000
0!
0%
#376715000000
1!
1%
#376720000000
0!
0%
#376725000000
1!
1%
#376730000000
0!
0%
#376735000000
1!
1%
#376740000000
0!
0%
#376745000000
1!
1%
#376750000000
0!
0%
#376755000000
1!
1%
#376760000000
0!
0%
#376765000000
1!
1%
#376770000000
0!
0%
#376775000000
1!
1%
#376780000000
0!
0%
#376785000000
1!
1%
#376790000000
0!
0%
#376795000000
1!
1%
#376800000000
0!
0%
#376805000000
1!
1%
#376810000000
0!
0%
#376815000000
1!
1%
#376820000000
0!
0%
#376825000000
1!
1%
#376830000000
0!
0%
#376835000000
1!
1%
#376840000000
0!
0%
#376845000000
1!
1%
#376850000000
0!
0%
#376855000000
1!
1%
#376860000000
0!
0%
#376865000000
1!
1%
#376870000000
0!
0%
#376875000000
1!
1%
#376880000000
0!
0%
#376885000000
1!
1%
#376890000000
0!
0%
#376895000000
1!
1%
#376900000000
0!
0%
#376905000000
1!
1%
#376910000000
0!
0%
#376915000000
1!
1%
#376920000000
0!
0%
#376925000000
1!
1%
#376930000000
0!
0%
#376935000000
1!
1%
#376940000000
0!
0%
#376945000000
1!
1%
#376950000000
0!
0%
#376955000000
1!
1%
#376960000000
0!
0%
#376965000000
1!
1%
#376970000000
0!
0%
#376975000000
1!
1%
#376980000000
0!
0%
#376985000000
1!
1%
#376990000000
0!
0%
#376995000000
1!
1%
#377000000000
0!
0%
#377005000000
1!
1%
#377010000000
0!
0%
#377015000000
1!
1%
#377020000000
0!
0%
#377025000000
1!
1%
#377030000000
0!
0%
#377035000000
1!
1%
#377040000000
0!
0%
#377045000000
1!
1%
#377050000000
0!
0%
#377055000000
1!
1%
#377060000000
0!
0%
#377065000000
1!
1%
#377070000000
0!
0%
#377075000000
1!
1%
#377080000000
0!
0%
#377085000000
1!
1%
#377090000000
0!
0%
#377095000000
1!
1%
#377100000000
0!
0%
#377105000000
1!
1%
#377110000000
0!
0%
#377115000000
1!
1%
#377120000000
0!
0%
#377125000000
1!
1%
#377130000000
0!
0%
#377135000000
1!
1%
#377140000000
0!
0%
#377145000000
1!
1%
#377150000000
0!
0%
#377155000000
1!
1%
#377160000000
0!
0%
#377165000000
1!
1%
#377170000000
0!
0%
#377175000000
1!
1%
#377180000000
0!
0%
#377185000000
1!
1%
#377190000000
0!
0%
#377195000000
1!
1%
#377200000000
0!
0%
#377205000000
1!
1%
#377210000000
0!
0%
#377215000000
1!
1%
#377220000000
0!
0%
#377225000000
1!
1%
#377230000000
0!
0%
#377235000000
1!
1%
#377240000000
0!
0%
#377245000000
1!
1%
#377250000000
0!
0%
#377255000000
1!
1%
#377260000000
0!
0%
#377265000000
1!
1%
#377270000000
0!
0%
#377275000000
1!
1%
#377280000000
0!
0%
#377285000000
1!
1%
#377290000000
0!
0%
#377295000000
1!
1%
#377300000000
0!
0%
#377305000000
1!
1%
#377310000000
0!
0%
#377315000000
1!
1%
#377320000000
0!
0%
#377325000000
1!
1%
#377330000000
0!
0%
#377335000000
1!
1%
#377340000000
0!
0%
#377345000000
1!
1%
#377350000000
0!
0%
#377355000000
1!
1%
#377360000000
0!
0%
#377365000000
1!
1%
#377370000000
0!
0%
#377375000000
1!
1%
#377380000000
0!
0%
#377385000000
1!
1%
#377390000000
0!
0%
#377395000000
1!
1%
#377400000000
0!
0%
#377405000000
1!
1%
#377410000000
0!
0%
#377415000000
1!
1%
#377420000000
0!
0%
#377425000000
1!
1%
#377430000000
0!
0%
#377435000000
1!
1%
#377440000000
0!
0%
#377445000000
1!
1%
#377450000000
0!
0%
#377455000000
1!
1%
#377460000000
0!
0%
#377465000000
1!
1%
#377470000000
0!
0%
#377475000000
1!
1%
#377480000000
0!
0%
#377485000000
1!
1%
#377490000000
0!
0%
#377495000000
1!
1%
#377500000000
0!
0%
#377505000000
1!
1%
#377510000000
0!
0%
#377515000000
1!
1%
#377520000000
0!
0%
#377525000000
1!
1%
#377530000000
0!
0%
#377535000000
1!
1%
#377540000000
0!
0%
#377545000000
1!
1%
#377550000000
0!
0%
#377555000000
1!
1%
#377560000000
0!
0%
#377565000000
1!
1%
#377570000000
0!
0%
#377575000000
1!
1%
#377580000000
0!
0%
#377585000000
1!
1%
#377590000000
0!
0%
#377595000000
1!
1%
#377600000000
0!
0%
#377605000000
1!
1%
#377610000000
0!
0%
#377615000000
1!
1%
#377620000000
0!
0%
#377625000000
1!
1%
#377630000000
0!
0%
#377635000000
1!
1%
#377640000000
0!
0%
#377645000000
1!
1%
#377650000000
0!
0%
#377655000000
1!
1%
#377660000000
0!
0%
#377665000000
1!
1%
#377670000000
0!
0%
#377675000000
1!
1%
#377680000000
0!
0%
#377685000000
1!
1%
#377690000000
0!
0%
#377695000000
1!
1%
#377700000000
0!
0%
#377705000000
1!
1%
#377710000000
0!
0%
#377715000000
1!
1%
#377720000000
0!
0%
#377725000000
1!
1%
#377730000000
0!
0%
#377735000000
1!
1%
#377740000000
0!
0%
#377745000000
1!
1%
#377750000000
0!
0%
#377755000000
1!
1%
#377760000000
0!
0%
#377765000000
1!
1%
#377770000000
0!
0%
#377775000000
1!
1%
#377780000000
0!
0%
#377785000000
1!
1%
#377790000000
0!
0%
#377795000000
1!
1%
#377800000000
0!
0%
#377805000000
1!
1%
#377810000000
0!
0%
#377815000000
1!
1%
#377820000000
0!
0%
#377825000000
1!
1%
#377830000000
0!
0%
#377835000000
1!
1%
#377840000000
0!
0%
#377845000000
1!
1%
#377850000000
0!
0%
#377855000000
1!
1%
#377860000000
0!
0%
#377865000000
1!
1%
#377870000000
0!
0%
#377875000000
1!
1%
#377880000000
0!
0%
#377885000000
1!
1%
#377890000000
0!
0%
#377895000000
1!
1%
#377900000000
0!
0%
#377905000000
1!
1%
#377910000000
0!
0%
#377915000000
1!
1%
#377920000000
0!
0%
#377925000000
1!
1%
#377930000000
0!
0%
#377935000000
1!
1%
#377940000000
0!
0%
#377945000000
1!
1%
#377950000000
0!
0%
#377955000000
1!
1%
#377960000000
0!
0%
#377965000000
1!
1%
#377970000000
0!
0%
#377975000000
1!
1%
#377980000000
0!
0%
#377985000000
1!
1%
#377990000000
0!
0%
#377995000000
1!
1%
#378000000000
0!
0%
#378005000000
1!
1%
#378010000000
0!
0%
#378015000000
1!
1%
#378020000000
0!
0%
#378025000000
1!
1%
#378030000000
0!
0%
#378035000000
1!
1%
#378040000000
0!
0%
#378045000000
1!
1%
#378050000000
0!
0%
#378055000000
1!
1%
#378060000000
0!
0%
#378065000000
1!
1%
#378070000000
0!
0%
#378075000000
1!
1%
#378080000000
0!
0%
#378085000000
1!
1%
#378090000000
0!
0%
#378095000000
1!
1%
#378100000000
0!
0%
#378105000000
1!
1%
#378110000000
0!
0%
#378115000000
1!
1%
#378120000000
0!
0%
#378125000000
1!
1%
#378130000000
0!
0%
#378135000000
1!
1%
#378140000000
0!
0%
#378145000000
1!
1%
#378150000000
0!
0%
#378155000000
1!
1%
#378160000000
0!
0%
#378165000000
1!
1%
#378170000000
0!
0%
#378175000000
1!
1%
#378180000000
0!
0%
#378185000000
1!
1%
#378190000000
0!
0%
#378195000000
1!
1%
#378200000000
0!
0%
#378205000000
1!
1%
#378210000000
0!
0%
#378215000000
1!
1%
#378220000000
0!
0%
#378225000000
1!
1%
#378230000000
0!
0%
#378235000000
1!
1%
#378240000000
0!
0%
#378245000000
1!
1%
#378250000000
0!
0%
#378255000000
1!
1%
#378260000000
0!
0%
#378265000000
1!
1%
#378270000000
0!
0%
#378275000000
1!
1%
#378280000000
0!
0%
#378285000000
1!
1%
#378290000000
0!
0%
#378295000000
1!
1%
#378300000000
0!
0%
#378305000000
1!
1%
#378310000000
0!
0%
#378315000000
1!
1%
#378320000000
0!
0%
#378325000000
1!
1%
#378330000000
0!
0%
#378335000000
1!
1%
#378340000000
0!
0%
#378345000000
1!
1%
#378350000000
0!
0%
#378355000000
1!
1%
#378360000000
0!
0%
#378365000000
1!
1%
#378370000000
0!
0%
#378375000000
1!
1%
#378380000000
0!
0%
#378385000000
1!
1%
#378390000000
0!
0%
#378395000000
1!
1%
#378400000000
0!
0%
#378405000000
1!
1%
#378410000000
0!
0%
#378415000000
1!
1%
#378420000000
0!
0%
#378425000000
1!
1%
#378430000000
0!
0%
#378435000000
1!
1%
#378440000000
0!
0%
#378445000000
1!
1%
#378450000000
0!
0%
#378455000000
1!
1%
#378460000000
0!
0%
#378465000000
1!
1%
#378470000000
0!
0%
#378475000000
1!
1%
#378480000000
0!
0%
#378485000000
1!
1%
#378490000000
0!
0%
#378495000000
1!
1%
#378500000000
0!
0%
#378505000000
1!
1%
#378510000000
0!
0%
#378515000000
1!
1%
#378520000000
0!
0%
#378525000000
1!
1%
#378530000000
0!
0%
#378535000000
1!
1%
#378540000000
0!
0%
#378545000000
1!
1%
#378550000000
0!
0%
#378555000000
1!
1%
#378560000000
0!
0%
#378565000000
1!
1%
#378570000000
0!
0%
#378575000000
1!
1%
#378580000000
0!
0%
#378585000000
1!
1%
#378590000000
0!
0%
#378595000000
1!
1%
#378600000000
0!
0%
#378605000000
1!
1%
#378610000000
0!
0%
#378615000000
1!
1%
#378620000000
0!
0%
#378625000000
1!
1%
#378630000000
0!
0%
#378635000000
1!
1%
#378640000000
0!
0%
#378645000000
1!
1%
#378650000000
0!
0%
#378655000000
1!
1%
#378660000000
0!
0%
#378665000000
1!
1%
#378670000000
0!
0%
#378675000000
1!
1%
#378680000000
0!
0%
#378685000000
1!
1%
#378690000000
0!
0%
#378695000000
1!
1%
#378700000000
0!
0%
#378705000000
1!
1%
#378710000000
0!
0%
#378715000000
1!
1%
#378720000000
0!
0%
#378725000000
1!
1%
#378730000000
0!
0%
#378735000000
1!
1%
#378740000000
0!
0%
#378745000000
1!
1%
#378750000000
0!
0%
#378755000000
1!
1%
#378760000000
0!
0%
#378765000000
1!
1%
#378770000000
0!
0%
#378775000000
1!
1%
#378780000000
0!
0%
#378785000000
1!
1%
#378790000000
0!
0%
#378795000000
1!
1%
#378800000000
0!
0%
#378805000000
1!
1%
#378810000000
0!
0%
#378815000000
1!
1%
#378820000000
0!
0%
#378825000000
1!
1%
#378830000000
0!
0%
#378835000000
1!
1%
#378840000000
0!
0%
#378845000000
1!
1%
#378850000000
0!
0%
#378855000000
1!
1%
#378860000000
0!
0%
#378865000000
1!
1%
#378870000000
0!
0%
#378875000000
1!
1%
#378880000000
0!
0%
#378885000000
1!
1%
#378890000000
0!
0%
#378895000000
1!
1%
#378900000000
0!
0%
#378905000000
1!
1%
#378910000000
0!
0%
#378915000000
1!
1%
#378920000000
0!
0%
#378925000000
1!
1%
#378930000000
0!
0%
#378935000000
1!
1%
#378940000000
0!
0%
#378945000000
1!
1%
#378950000000
0!
0%
#378955000000
1!
1%
#378960000000
0!
0%
#378965000000
1!
1%
#378970000000
0!
0%
#378975000000
1!
1%
#378980000000
0!
0%
#378985000000
1!
1%
#378990000000
0!
0%
#378995000000
1!
1%
#379000000000
0!
0%
#379005000000
1!
1%
#379010000000
0!
0%
#379015000000
1!
1%
#379020000000
0!
0%
#379025000000
1!
1%
#379030000000
0!
0%
#379035000000
1!
1%
#379040000000
0!
0%
#379045000000
1!
1%
#379050000000
0!
0%
#379055000000
1!
1%
#379060000000
0!
0%
#379065000000
1!
1%
#379070000000
0!
0%
#379075000000
1!
1%
#379080000000
0!
0%
#379085000000
1!
1%
#379090000000
0!
0%
#379095000000
1!
1%
#379100000000
0!
0%
#379105000000
1!
1%
#379110000000
0!
0%
#379115000000
1!
1%
#379120000000
0!
0%
#379125000000
1!
1%
#379130000000
0!
0%
#379135000000
1!
1%
#379140000000
0!
0%
#379145000000
1!
1%
#379150000000
0!
0%
#379155000000
1!
1%
#379160000000
0!
0%
#379165000000
1!
1%
#379170000000
0!
0%
#379175000000
1!
1%
#379180000000
0!
0%
#379185000000
1!
1%
#379190000000
0!
0%
#379195000000
1!
1%
#379200000000
0!
0%
#379205000000
1!
1%
#379210000000
0!
0%
#379215000000
1!
1%
#379220000000
0!
0%
#379225000000
1!
1%
#379230000000
0!
0%
#379235000000
1!
1%
#379240000000
0!
0%
#379245000000
1!
1%
#379250000000
0!
0%
#379255000000
1!
1%
#379260000000
0!
0%
#379265000000
1!
1%
#379270000000
0!
0%
#379275000000
1!
1%
#379280000000
0!
0%
#379285000000
1!
1%
#379290000000
0!
0%
#379295000000
1!
1%
#379300000000
0!
0%
#379305000000
1!
1%
#379310000000
0!
0%
#379315000000
1!
1%
#379320000000
0!
0%
#379325000000
1!
1%
#379330000000
0!
0%
#379335000000
1!
1%
#379340000000
0!
0%
#379345000000
1!
1%
#379350000000
0!
0%
#379355000000
1!
1%
#379360000000
0!
0%
#379365000000
1!
1%
#379370000000
0!
0%
#379375000000
1!
1%
#379380000000
0!
0%
#379385000000
1!
1%
#379390000000
0!
0%
#379395000000
1!
1%
#379400000000
0!
0%
#379405000000
1!
1%
#379410000000
0!
0%
#379415000000
1!
1%
#379420000000
0!
0%
#379425000000
1!
1%
#379430000000
0!
0%
#379435000000
1!
1%
#379440000000
0!
0%
#379445000000
1!
1%
#379450000000
0!
0%
#379455000000
1!
1%
#379460000000
0!
0%
#379465000000
1!
1%
#379470000000
0!
0%
#379475000000
1!
1%
#379480000000
0!
0%
#379485000000
1!
1%
#379490000000
0!
0%
#379495000000
1!
1%
#379500000000
0!
0%
#379505000000
1!
1%
#379510000000
0!
0%
#379515000000
1!
1%
#379520000000
0!
0%
#379525000000
1!
1%
#379530000000
0!
0%
#379535000000
1!
1%
#379540000000
0!
0%
#379545000000
1!
1%
#379550000000
0!
0%
#379555000000
1!
1%
#379560000000
0!
0%
#379565000000
1!
1%
#379570000000
0!
0%
#379575000000
1!
1%
#379580000000
0!
0%
#379585000000
1!
1%
#379590000000
0!
0%
#379595000000
1!
1%
#379600000000
0!
0%
#379605000000
1!
1%
#379610000000
0!
0%
#379615000000
1!
1%
#379620000000
0!
0%
#379625000000
1!
1%
#379630000000
0!
0%
#379635000000
1!
1%
#379640000000
0!
0%
#379645000000
1!
1%
#379650000000
0!
0%
#379655000000
1!
1%
#379660000000
0!
0%
#379665000000
1!
1%
#379670000000
0!
0%
#379675000000
1!
1%
#379680000000
0!
0%
#379685000000
1!
1%
#379690000000
0!
0%
#379695000000
1!
1%
#379700000000
0!
0%
#379705000000
1!
1%
#379710000000
0!
0%
#379715000000
1!
1%
#379720000000
0!
0%
#379725000000
1!
1%
#379730000000
0!
0%
#379735000000
1!
1%
#379740000000
0!
0%
#379745000000
1!
1%
#379750000000
0!
0%
#379755000000
1!
1%
#379760000000
0!
0%
#379765000000
1!
1%
#379770000000
0!
0%
#379775000000
1!
1%
#379780000000
0!
0%
#379785000000
1!
1%
#379790000000
0!
0%
#379795000000
1!
1%
#379800000000
0!
0%
#379805000000
1!
1%
#379810000000
0!
0%
#379815000000
1!
1%
#379820000000
0!
0%
#379825000000
1!
1%
#379830000000
0!
0%
#379835000000
1!
1%
#379840000000
0!
0%
#379845000000
1!
1%
#379850000000
0!
0%
#379855000000
1!
1%
#379860000000
0!
0%
#379865000000
1!
1%
#379870000000
0!
0%
#379875000000
1!
1%
#379880000000
0!
0%
#379885000000
1!
1%
#379890000000
0!
0%
#379895000000
1!
1%
#379900000000
0!
0%
#379905000000
1!
1%
#379910000000
0!
0%
#379915000000
1!
1%
#379920000000
0!
0%
#379925000000
1!
1%
#379930000000
0!
0%
#379935000000
1!
1%
#379940000000
0!
0%
#379945000000
1!
1%
#379950000000
0!
0%
#379955000000
1!
1%
#379960000000
0!
0%
#379965000000
1!
1%
#379970000000
0!
0%
#379975000000
1!
1%
#379980000000
0!
0%
#379985000000
1!
1%
#379990000000
0!
0%
#379995000000
1!
1%
#380000000000
0!
0%
#380005000000
1!
1%
#380010000000
0!
0%
#380015000000
1!
1%
#380020000000
0!
0%
#380025000000
1!
1%
#380030000000
0!
0%
#380035000000
1!
1%
#380040000000
0!
0%
#380045000000
1!
1%
#380050000000
0!
0%
#380055000000
1!
1%
#380060000000
0!
0%
#380065000000
1!
1%
#380070000000
0!
0%
#380075000000
1!
1%
#380080000000
0!
0%
#380085000000
1!
1%
#380090000000
0!
0%
#380095000000
1!
1%
#380100000000
0!
0%
#380105000000
1!
1%
#380110000000
0!
0%
#380115000000
1!
1%
#380120000000
0!
0%
#380125000000
1!
1%
#380130000000
0!
0%
#380135000000
1!
1%
#380140000000
0!
0%
#380145000000
1!
1%
#380150000000
0!
0%
#380155000000
1!
1%
#380160000000
0!
0%
#380165000000
1!
1%
#380170000000
0!
0%
#380175000000
1!
1%
#380180000000
0!
0%
#380185000000
1!
1%
#380190000000
0!
0%
#380195000000
1!
1%
#380200000000
0!
0%
#380205000000
1!
1%
#380210000000
0!
0%
#380215000000
1!
1%
#380220000000
0!
0%
#380225000000
1!
1%
#380230000000
0!
0%
#380235000000
1!
1%
#380240000000
0!
0%
#380245000000
1!
1%
#380250000000
0!
0%
#380255000000
1!
1%
#380260000000
0!
0%
#380265000000
1!
1%
#380270000000
0!
0%
#380275000000
1!
1%
#380280000000
0!
0%
#380285000000
1!
1%
#380290000000
0!
0%
#380295000000
1!
1%
#380300000000
0!
0%
#380305000000
1!
1%
#380310000000
0!
0%
#380315000000
1!
1%
#380320000000
0!
0%
#380325000000
1!
1%
#380330000000
0!
0%
#380335000000
1!
1%
#380340000000
0!
0%
#380345000000
1!
1%
#380350000000
0!
0%
#380355000000
1!
1%
#380360000000
0!
0%
#380365000000
1!
1%
#380370000000
0!
0%
#380375000000
1!
1%
#380380000000
0!
0%
#380385000000
1!
1%
#380390000000
0!
0%
#380395000000
1!
1%
#380400000000
0!
0%
#380405000000
1!
1%
#380410000000
0!
0%
#380415000000
1!
1%
#380420000000
0!
0%
#380425000000
1!
1%
#380430000000
0!
0%
#380435000000
1!
1%
#380440000000
0!
0%
#380445000000
1!
1%
#380450000000
0!
0%
#380455000000
1!
1%
#380460000000
0!
0%
#380465000000
1!
1%
#380470000000
0!
0%
#380475000000
1!
1%
#380480000000
0!
0%
#380485000000
1!
1%
#380490000000
0!
0%
#380495000000
1!
1%
#380500000000
0!
0%
#380505000000
1!
1%
#380510000000
0!
0%
#380515000000
1!
1%
#380520000000
0!
0%
#380525000000
1!
1%
#380530000000
0!
0%
#380535000000
1!
1%
#380540000000
0!
0%
#380545000000
1!
1%
#380550000000
0!
0%
#380555000000
1!
1%
#380560000000
0!
0%
#380565000000
1!
1%
#380570000000
0!
0%
#380575000000
1!
1%
#380580000000
0!
0%
#380585000000
1!
1%
#380590000000
0!
0%
#380595000000
1!
1%
#380600000000
0!
0%
#380605000000
1!
1%
#380610000000
0!
0%
#380615000000
1!
1%
#380620000000
0!
0%
#380625000000
1!
1%
#380630000000
0!
0%
#380635000000
1!
1%
#380640000000
0!
0%
#380645000000
1!
1%
#380650000000
0!
0%
#380655000000
1!
1%
#380660000000
0!
0%
#380665000000
1!
1%
#380670000000
0!
0%
#380675000000
1!
1%
#380680000000
0!
0%
#380685000000
1!
1%
#380690000000
0!
0%
#380695000000
1!
1%
#380700000000
0!
0%
#380705000000
1!
1%
#380710000000
0!
0%
#380715000000
1!
1%
#380720000000
0!
0%
#380725000000
1!
1%
#380730000000
0!
0%
#380735000000
1!
1%
#380740000000
0!
0%
#380745000000
1!
1%
#380750000000
0!
0%
#380755000000
1!
1%
#380760000000
0!
0%
#380765000000
1!
1%
#380770000000
0!
0%
#380775000000
1!
1%
#380780000000
0!
0%
#380785000000
1!
1%
#380790000000
0!
0%
#380795000000
1!
1%
#380800000000
0!
0%
#380805000000
1!
1%
#380810000000
0!
0%
#380815000000
1!
1%
#380820000000
0!
0%
#380825000000
1!
1%
#380830000000
0!
0%
#380835000000
1!
1%
#380840000000
0!
0%
#380845000000
1!
1%
#380850000000
0!
0%
#380855000000
1!
1%
#380860000000
0!
0%
#380865000000
1!
1%
#380870000000
0!
0%
#380875000000
1!
1%
#380880000000
0!
0%
#380885000000
1!
1%
#380890000000
0!
0%
#380895000000
1!
1%
#380900000000
0!
0%
#380905000000
1!
1%
#380910000000
0!
0%
#380915000000
1!
1%
#380920000000
0!
0%
#380925000000
1!
1%
#380930000000
0!
0%
#380935000000
1!
1%
#380940000000
0!
0%
#380945000000
1!
1%
#380950000000
0!
0%
#380955000000
1!
1%
#380960000000
0!
0%
#380965000000
1!
1%
#380970000000
0!
0%
#380975000000
1!
1%
#380980000000
0!
0%
#380985000000
1!
1%
#380990000000
0!
0%
#380995000000
1!
1%
#381000000000
0!
0%
#381005000000
1!
1%
#381010000000
0!
0%
#381015000000
1!
1%
#381020000000
0!
0%
#381025000000
1!
1%
#381030000000
0!
0%
#381035000000
1!
1%
#381040000000
0!
0%
#381045000000
1!
1%
#381050000000
0!
0%
#381055000000
1!
1%
#381060000000
0!
0%
#381065000000
1!
1%
#381070000000
0!
0%
#381075000000
1!
1%
#381080000000
0!
0%
#381085000000
1!
1%
#381090000000
0!
0%
#381095000000
1!
1%
#381100000000
0!
0%
#381105000000
1!
1%
#381110000000
0!
0%
#381115000000
1!
1%
#381120000000
0!
0%
#381125000000
1!
1%
#381130000000
0!
0%
#381135000000
1!
1%
#381140000000
0!
0%
#381145000000
1!
1%
#381150000000
0!
0%
#381155000000
1!
1%
#381160000000
0!
0%
#381165000000
1!
1%
#381170000000
0!
0%
#381175000000
1!
1%
#381180000000
0!
0%
#381185000000
1!
1%
#381190000000
0!
0%
#381195000000
1!
1%
#381200000000
0!
0%
#381205000000
1!
1%
#381210000000
0!
0%
#381215000000
1!
1%
#381220000000
0!
0%
#381225000000
1!
1%
#381230000000
0!
0%
#381235000000
1!
1%
#381240000000
0!
0%
#381245000000
1!
1%
#381250000000
0!
0%
#381255000000
1!
1%
#381260000000
0!
0%
#381265000000
1!
1%
#381270000000
0!
0%
#381275000000
1!
1%
#381280000000
0!
0%
#381285000000
1!
1%
#381290000000
0!
0%
#381295000000
1!
1%
#381300000000
0!
0%
#381305000000
1!
1%
#381310000000
0!
0%
#381315000000
1!
1%
#381320000000
0!
0%
#381325000000
1!
1%
#381330000000
0!
0%
#381335000000
1!
1%
#381340000000
0!
0%
#381345000000
1!
1%
#381350000000
0!
0%
#381355000000
1!
1%
#381360000000
0!
0%
#381365000000
1!
1%
#381370000000
0!
0%
#381375000000
1!
1%
#381380000000
0!
0%
#381385000000
1!
1%
#381390000000
0!
0%
#381395000000
1!
1%
#381400000000
0!
0%
#381405000000
1!
1%
#381410000000
0!
0%
#381415000000
1!
1%
#381420000000
0!
0%
#381425000000
1!
1%
#381430000000
0!
0%
#381435000000
1!
1%
#381440000000
0!
0%
#381445000000
1!
1%
#381450000000
0!
0%
#381455000000
1!
1%
#381460000000
0!
0%
#381465000000
1!
1%
#381470000000
0!
0%
#381475000000
1!
1%
#381480000000
0!
0%
#381485000000
1!
1%
#381490000000
0!
0%
#381495000000
1!
1%
#381500000000
0!
0%
#381505000000
1!
1%
#381510000000
0!
0%
#381515000000
1!
1%
#381520000000
0!
0%
#381525000000
1!
1%
#381530000000
0!
0%
#381535000000
1!
1%
#381540000000
0!
0%
#381545000000
1!
1%
#381550000000
0!
0%
#381555000000
1!
1%
#381560000000
0!
0%
#381565000000
1!
1%
#381570000000
0!
0%
#381575000000
1!
1%
#381580000000
0!
0%
#381585000000
1!
1%
#381590000000
0!
0%
#381595000000
1!
1%
#381600000000
0!
0%
#381605000000
1!
1%
#381610000000
0!
0%
#381615000000
1!
1%
#381620000000
0!
0%
#381625000000
1!
1%
#381630000000
0!
0%
#381635000000
1!
1%
#381640000000
0!
0%
#381645000000
1!
1%
#381650000000
0!
0%
#381655000000
1!
1%
#381660000000
0!
0%
#381665000000
1!
1%
#381670000000
0!
0%
#381675000000
1!
1%
#381680000000
0!
0%
#381685000000
1!
1%
#381690000000
0!
0%
#381695000000
1!
1%
#381700000000
0!
0%
#381705000000
1!
1%
#381710000000
0!
0%
#381715000000
1!
1%
#381720000000
0!
0%
#381725000000
1!
1%
#381730000000
0!
0%
#381735000000
1!
1%
#381740000000
0!
0%
#381745000000
1!
1%
#381750000000
0!
0%
#381755000000
1!
1%
#381760000000
0!
0%
#381765000000
1!
1%
#381770000000
0!
0%
#381775000000
1!
1%
#381780000000
0!
0%
#381785000000
1!
1%
#381790000000
0!
0%
#381795000000
1!
1%
#381800000000
0!
0%
#381805000000
1!
1%
#381810000000
0!
0%
#381815000000
1!
1%
#381820000000
0!
0%
#381825000000
1!
1%
#381830000000
0!
0%
#381835000000
1!
1%
#381840000000
0!
0%
#381845000000
1!
1%
#381850000000
0!
0%
#381855000000
1!
1%
#381860000000
0!
0%
#381865000000
1!
1%
#381870000000
0!
0%
#381875000000
1!
1%
#381880000000
0!
0%
#381885000000
1!
1%
#381890000000
0!
0%
#381895000000
1!
1%
#381900000000
0!
0%
#381905000000
1!
1%
#381910000000
0!
0%
#381915000000
1!
1%
#381920000000
0!
0%
#381925000000
1!
1%
#381930000000
0!
0%
#381935000000
1!
1%
#381940000000
0!
0%
#381945000000
1!
1%
#381950000000
0!
0%
#381955000000
1!
1%
#381960000000
0!
0%
#381965000000
1!
1%
#381970000000
0!
0%
#381975000000
1!
1%
#381980000000
0!
0%
#381985000000
1!
1%
#381990000000
0!
0%
#381995000000
1!
1%
#382000000000
0!
0%
#382005000000
1!
1%
#382010000000
0!
0%
#382015000000
1!
1%
#382020000000
0!
0%
#382025000000
1!
1%
#382030000000
0!
0%
#382035000000
1!
1%
#382040000000
0!
0%
#382045000000
1!
1%
#382050000000
0!
0%
#382055000000
1!
1%
#382060000000
0!
0%
#382065000000
1!
1%
#382070000000
0!
0%
#382075000000
1!
1%
#382080000000
0!
0%
#382085000000
1!
1%
#382090000000
0!
0%
#382095000000
1!
1%
#382100000000
0!
0%
#382105000000
1!
1%
#382110000000
0!
0%
#382115000000
1!
1%
#382120000000
0!
0%
#382125000000
1!
1%
#382130000000
0!
0%
#382135000000
1!
1%
#382140000000
0!
0%
#382145000000
1!
1%
#382150000000
0!
0%
#382155000000
1!
1%
#382160000000
0!
0%
#382165000000
1!
1%
#382170000000
0!
0%
#382175000000
1!
1%
#382180000000
0!
0%
#382185000000
1!
1%
#382190000000
0!
0%
#382195000000
1!
1%
#382200000000
0!
0%
#382205000000
1!
1%
#382210000000
0!
0%
#382215000000
1!
1%
#382220000000
0!
0%
#382225000000
1!
1%
#382230000000
0!
0%
#382235000000
1!
1%
#382240000000
0!
0%
#382245000000
1!
1%
#382250000000
0!
0%
#382255000000
1!
1%
#382260000000
0!
0%
#382265000000
1!
1%
#382270000000
0!
0%
#382275000000
1!
1%
#382280000000
0!
0%
#382285000000
1!
1%
#382290000000
0!
0%
#382295000000
1!
1%
#382300000000
0!
0%
#382305000000
1!
1%
#382310000000
0!
0%
#382315000000
1!
1%
#382320000000
0!
0%
#382325000000
1!
1%
#382330000000
0!
0%
#382335000000
1!
1%
#382340000000
0!
0%
#382345000000
1!
1%
#382350000000
0!
0%
#382355000000
1!
1%
#382360000000
0!
0%
#382365000000
1!
1%
#382370000000
0!
0%
#382375000000
1!
1%
#382380000000
0!
0%
#382385000000
1!
1%
#382390000000
0!
0%
#382395000000
1!
1%
#382400000000
0!
0%
#382405000000
1!
1%
#382410000000
0!
0%
#382415000000
1!
1%
#382420000000
0!
0%
#382425000000
1!
1%
#382430000000
0!
0%
#382435000000
1!
1%
#382440000000
0!
0%
#382445000000
1!
1%
#382450000000
0!
0%
#382455000000
1!
1%
#382460000000
0!
0%
#382465000000
1!
1%
#382470000000
0!
0%
#382475000000
1!
1%
#382480000000
0!
0%
#382485000000
1!
1%
#382490000000
0!
0%
#382495000000
1!
1%
#382500000000
0!
0%
#382505000000
1!
1%
#382510000000
0!
0%
#382515000000
1!
1%
#382520000000
0!
0%
#382525000000
1!
1%
#382530000000
0!
0%
#382535000000
1!
1%
#382540000000
0!
0%
#382545000000
1!
1%
#382550000000
0!
0%
#382555000000
1!
1%
#382560000000
0!
0%
#382565000000
1!
1%
#382570000000
0!
0%
#382575000000
1!
1%
#382580000000
0!
0%
#382585000000
1!
1%
#382590000000
0!
0%
#382595000000
1!
1%
#382600000000
0!
0%
#382605000000
1!
1%
#382610000000
0!
0%
#382615000000
1!
1%
#382620000000
0!
0%
#382625000000
1!
1%
#382630000000
0!
0%
#382635000000
1!
1%
#382640000000
0!
0%
#382645000000
1!
1%
#382650000000
0!
0%
#382655000000
1!
1%
#382660000000
0!
0%
#382665000000
1!
1%
#382670000000
0!
0%
#382675000000
1!
1%
#382680000000
0!
0%
#382685000000
1!
1%
#382690000000
0!
0%
#382695000000
1!
1%
#382700000000
0!
0%
#382705000000
1!
1%
#382710000000
0!
0%
#382715000000
1!
1%
#382720000000
0!
0%
#382725000000
1!
1%
#382730000000
0!
0%
#382735000000
1!
1%
#382740000000
0!
0%
#382745000000
1!
1%
#382750000000
0!
0%
#382755000000
1!
1%
#382760000000
0!
0%
#382765000000
1!
1%
#382770000000
0!
0%
#382775000000
1!
1%
#382780000000
0!
0%
#382785000000
1!
1%
#382790000000
0!
0%
#382795000000
1!
1%
#382800000000
0!
0%
#382805000000
1!
1%
#382810000000
0!
0%
#382815000000
1!
1%
#382820000000
0!
0%
#382825000000
1!
1%
#382830000000
0!
0%
#382835000000
1!
1%
#382840000000
0!
0%
#382845000000
1!
1%
#382850000000
0!
0%
#382855000000
1!
1%
#382860000000
0!
0%
#382865000000
1!
1%
#382870000000
0!
0%
#382875000000
1!
1%
#382880000000
0!
0%
#382885000000
1!
1%
#382890000000
0!
0%
#382895000000
1!
1%
#382900000000
0!
0%
#382905000000
1!
1%
#382910000000
0!
0%
#382915000000
1!
1%
#382920000000
0!
0%
#382925000000
1!
1%
#382930000000
0!
0%
#382935000000
1!
1%
#382940000000
0!
0%
#382945000000
1!
1%
#382950000000
0!
0%
#382955000000
1!
1%
#382960000000
0!
0%
#382965000000
1!
1%
#382970000000
0!
0%
#382975000000
1!
1%
#382980000000
0!
0%
#382985000000
1!
1%
#382990000000
0!
0%
#382995000000
1!
1%
#383000000000
0!
0%
#383005000000
1!
1%
#383010000000
0!
0%
#383015000000
1!
1%
#383020000000
0!
0%
#383025000000
1!
1%
#383030000000
0!
0%
#383035000000
1!
1%
#383040000000
0!
0%
#383045000000
1!
1%
#383050000000
0!
0%
#383055000000
1!
1%
#383060000000
0!
0%
#383065000000
1!
1%
#383070000000
0!
0%
#383075000000
1!
1%
#383080000000
0!
0%
#383085000000
1!
1%
#383090000000
0!
0%
#383095000000
1!
1%
#383100000000
0!
0%
#383105000000
1!
1%
#383110000000
0!
0%
#383115000000
1!
1%
#383120000000
0!
0%
#383125000000
1!
1%
#383130000000
0!
0%
#383135000000
1!
1%
#383140000000
0!
0%
#383145000000
1!
1%
#383150000000
0!
0%
#383155000000
1!
1%
#383160000000
0!
0%
#383165000000
1!
1%
#383170000000
0!
0%
#383175000000
1!
1%
#383180000000
0!
0%
#383185000000
1!
1%
#383190000000
0!
0%
#383195000000
1!
1%
#383200000000
0!
0%
#383205000000
1!
1%
#383210000000
0!
0%
#383215000000
1!
1%
#383220000000
0!
0%
#383225000000
1!
1%
#383230000000
0!
0%
#383235000000
1!
1%
#383240000000
0!
0%
#383245000000
1!
1%
#383250000000
0!
0%
#383255000000
1!
1%
#383260000000
0!
0%
#383265000000
1!
1%
#383270000000
0!
0%
#383275000000
1!
1%
#383280000000
0!
0%
#383285000000
1!
1%
#383290000000
0!
0%
#383295000000
1!
1%
#383300000000
0!
0%
#383305000000
1!
1%
#383310000000
0!
0%
#383315000000
1!
1%
#383320000000
0!
0%
#383325000000
1!
1%
#383330000000
0!
0%
#383335000000
1!
1%
#383340000000
0!
0%
#383345000000
1!
1%
#383350000000
0!
0%
#383355000000
1!
1%
#383360000000
0!
0%
#383365000000
1!
1%
#383370000000
0!
0%
#383375000000
1!
1%
#383380000000
0!
0%
#383385000000
1!
1%
#383390000000
0!
0%
#383395000000
1!
1%
#383400000000
0!
0%
#383405000000
1!
1%
#383410000000
0!
0%
#383415000000
1!
1%
#383420000000
0!
0%
#383425000000
1!
1%
#383430000000
0!
0%
#383435000000
1!
1%
#383440000000
0!
0%
#383445000000
1!
1%
#383450000000
0!
0%
#383455000000
1!
1%
#383460000000
0!
0%
#383465000000
1!
1%
#383470000000
0!
0%
#383475000000
1!
1%
#383480000000
0!
0%
#383485000000
1!
1%
#383490000000
0!
0%
#383495000000
1!
1%
#383500000000
0!
0%
#383505000000
1!
1%
#383510000000
0!
0%
#383515000000
1!
1%
#383520000000
0!
0%
#383525000000
1!
1%
#383530000000
0!
0%
#383535000000
1!
1%
#383540000000
0!
0%
#383545000000
1!
1%
#383550000000
0!
0%
#383555000000
1!
1%
#383560000000
0!
0%
#383565000000
1!
1%
#383570000000
0!
0%
#383575000000
1!
1%
#383580000000
0!
0%
#383585000000
1!
1%
#383590000000
0!
0%
#383595000000
1!
1%
#383600000000
0!
0%
#383605000000
1!
1%
#383610000000
0!
0%
#383615000000
1!
1%
#383620000000
0!
0%
#383625000000
1!
1%
#383630000000
0!
0%
#383635000000
1!
1%
#383640000000
0!
0%
#383645000000
1!
1%
#383650000000
0!
0%
#383655000000
1!
1%
#383660000000
0!
0%
#383665000000
1!
1%
#383670000000
0!
0%
#383675000000
1!
1%
#383680000000
0!
0%
#383685000000
1!
1%
#383690000000
0!
0%
#383695000000
1!
1%
#383700000000
0!
0%
#383705000000
1!
1%
#383710000000
0!
0%
#383715000000
1!
1%
#383720000000
0!
0%
#383725000000
1!
1%
#383730000000
0!
0%
#383735000000
1!
1%
#383740000000
0!
0%
#383745000000
1!
1%
#383750000000
0!
0%
#383755000000
1!
1%
#383760000000
0!
0%
#383765000000
1!
1%
#383770000000
0!
0%
#383775000000
1!
1%
#383780000000
0!
0%
#383785000000
1!
1%
#383790000000
0!
0%
#383795000000
1!
1%
#383800000000
0!
0%
#383805000000
1!
1%
#383810000000
0!
0%
#383815000000
1!
1%
#383820000000
0!
0%
#383825000000
1!
1%
#383830000000
0!
0%
#383835000000
1!
1%
#383840000000
0!
0%
#383845000000
1!
1%
#383850000000
0!
0%
#383855000000
1!
1%
#383860000000
0!
0%
#383865000000
1!
1%
#383870000000
0!
0%
#383875000000
1!
1%
#383880000000
0!
0%
#383885000000
1!
1%
#383890000000
0!
0%
#383895000000
1!
1%
#383900000000
0!
0%
#383905000000
1!
1%
#383910000000
0!
0%
#383915000000
1!
1%
#383920000000
0!
0%
#383925000000
1!
1%
#383930000000
0!
0%
#383935000000
1!
1%
#383940000000
0!
0%
#383945000000
1!
1%
#383950000000
0!
0%
#383955000000
1!
1%
#383960000000
0!
0%
#383965000000
1!
1%
#383970000000
0!
0%
#383975000000
1!
1%
#383980000000
0!
0%
#383985000000
1!
1%
#383990000000
0!
0%
#383995000000
1!
1%
#384000000000
0!
0%
#384005000000
1!
1%
#384010000000
0!
0%
#384015000000
1!
1%
#384020000000
0!
0%
#384025000000
1!
1%
#384030000000
0!
0%
#384035000000
1!
1%
#384040000000
0!
0%
#384045000000
1!
1%
#384050000000
0!
0%
#384055000000
1!
1%
#384060000000
0!
0%
#384065000000
1!
1%
#384070000000
0!
0%
#384075000000
1!
1%
#384080000000
0!
0%
#384085000000
1!
1%
#384090000000
0!
0%
#384095000000
1!
1%
#384100000000
0!
0%
#384105000000
1!
1%
#384110000000
0!
0%
#384115000000
1!
1%
#384120000000
0!
0%
#384125000000
1!
1%
#384130000000
0!
0%
#384135000000
1!
1%
#384140000000
0!
0%
#384145000000
1!
1%
#384150000000
0!
0%
#384155000000
1!
1%
#384160000000
0!
0%
#384165000000
1!
1%
#384170000000
0!
0%
#384175000000
1!
1%
#384180000000
0!
0%
#384185000000
1!
1%
#384190000000
0!
0%
#384195000000
1!
1%
#384200000000
0!
0%
#384205000000
1!
1%
#384210000000
0!
0%
#384215000000
1!
1%
#384220000000
0!
0%
#384225000000
1!
1%
#384230000000
0!
0%
#384235000000
1!
1%
#384240000000
0!
0%
#384245000000
1!
1%
#384250000000
0!
0%
#384255000000
1!
1%
#384260000000
0!
0%
#384265000000
1!
1%
#384270000000
0!
0%
#384275000000
1!
1%
#384280000000
0!
0%
#384285000000
1!
1%
#384290000000
0!
0%
#384295000000
1!
1%
#384300000000
0!
0%
#384305000000
1!
1%
#384310000000
0!
0%
#384315000000
1!
1%
#384320000000
0!
0%
#384325000000
1!
1%
#384330000000
0!
0%
#384335000000
1!
1%
#384340000000
0!
0%
#384345000000
1!
1%
#384350000000
0!
0%
#384355000000
1!
1%
#384360000000
0!
0%
#384365000000
1!
1%
#384370000000
0!
0%
#384375000000
1!
1%
#384380000000
0!
0%
#384385000000
1!
1%
#384390000000
0!
0%
#384395000000
1!
1%
#384400000000
0!
0%
#384405000000
1!
1%
#384410000000
0!
0%
#384415000000
1!
1%
#384420000000
0!
0%
#384425000000
1!
1%
#384430000000
0!
0%
#384435000000
1!
1%
#384440000000
0!
0%
#384445000000
1!
1%
#384450000000
0!
0%
#384455000000
1!
1%
#384460000000
0!
0%
#384465000000
1!
1%
#384470000000
0!
0%
#384475000000
1!
1%
#384480000000
0!
0%
#384485000000
1!
1%
#384490000000
0!
0%
#384495000000
1!
1%
#384500000000
0!
0%
#384505000000
1!
1%
#384510000000
0!
0%
#384515000000
1!
1%
#384520000000
0!
0%
#384525000000
1!
1%
#384530000000
0!
0%
#384535000000
1!
1%
#384540000000
0!
0%
#384545000000
1!
1%
#384550000000
0!
0%
#384555000000
1!
1%
#384560000000
0!
0%
#384565000000
1!
1%
#384570000000
0!
0%
#384575000000
1!
1%
#384580000000
0!
0%
#384585000000
1!
1%
#384590000000
0!
0%
#384595000000
1!
1%
#384600000000
0!
0%
#384605000000
1!
1%
#384610000000
0!
0%
#384615000000
1!
1%
#384620000000
0!
0%
#384625000000
1!
1%
#384630000000
0!
0%
#384635000000
1!
1%
#384640000000
0!
0%
#384645000000
1!
1%
#384650000000
0!
0%
#384655000000
1!
1%
#384660000000
0!
0%
#384665000000
1!
1%
#384670000000
0!
0%
#384675000000
1!
1%
#384680000000
0!
0%
#384685000000
1!
1%
#384690000000
0!
0%
#384695000000
1!
1%
#384700000000
0!
0%
#384705000000
1!
1%
#384710000000
0!
0%
#384715000000
1!
1%
#384720000000
0!
0%
#384725000000
1!
1%
#384730000000
0!
0%
#384735000000
1!
1%
#384740000000
0!
0%
#384745000000
1!
1%
#384750000000
0!
0%
#384755000000
1!
1%
#384760000000
0!
0%
#384765000000
1!
1%
#384770000000
0!
0%
#384775000000
1!
1%
#384780000000
0!
0%
#384785000000
1!
1%
#384790000000
0!
0%
#384795000000
1!
1%
#384800000000
0!
0%
#384805000000
1!
1%
#384810000000
0!
0%
#384815000000
1!
1%
#384820000000
0!
0%
#384825000000
1!
1%
#384830000000
0!
0%
#384835000000
1!
1%
#384840000000
0!
0%
#384845000000
1!
1%
#384850000000
0!
0%
#384855000000
1!
1%
#384860000000
0!
0%
#384865000000
1!
1%
#384870000000
0!
0%
#384875000000
1!
1%
#384880000000
0!
0%
#384885000000
1!
1%
#384890000000
0!
0%
#384895000000
1!
1%
#384900000000
0!
0%
#384905000000
1!
1%
#384910000000
0!
0%
#384915000000
1!
1%
#384920000000
0!
0%
#384925000000
1!
1%
#384930000000
0!
0%
#384935000000
1!
1%
#384940000000
0!
0%
#384945000000
1!
1%
#384950000000
0!
0%
#384955000000
1!
1%
#384960000000
0!
0%
#384965000000
1!
1%
#384970000000
0!
0%
#384975000000
1!
1%
#384980000000
0!
0%
#384985000000
1!
1%
#384990000000
0!
0%
#384995000000
1!
1%
#385000000000
0!
0%
#385005000000
1!
1%
#385010000000
0!
0%
#385015000000
1!
1%
#385020000000
0!
0%
#385025000000
1!
1%
#385030000000
0!
0%
#385035000000
1!
1%
#385040000000
0!
0%
#385045000000
1!
1%
#385050000000
0!
0%
#385055000000
1!
1%
#385060000000
0!
0%
#385065000000
1!
1%
#385070000000
0!
0%
#385075000000
1!
1%
#385080000000
0!
0%
#385085000000
1!
1%
#385090000000
0!
0%
#385095000000
1!
1%
#385100000000
0!
0%
#385105000000
1!
1%
#385110000000
0!
0%
#385115000000
1!
1%
#385120000000
0!
0%
#385125000000
1!
1%
#385130000000
0!
0%
#385135000000
1!
1%
#385140000000
0!
0%
#385145000000
1!
1%
#385150000000
0!
0%
#385155000000
1!
1%
#385160000000
0!
0%
#385165000000
1!
1%
#385170000000
0!
0%
#385175000000
1!
1%
#385180000000
0!
0%
#385185000000
1!
1%
#385190000000
0!
0%
#385195000000
1!
1%
#385200000000
0!
0%
#385205000000
1!
1%
#385210000000
0!
0%
#385215000000
1!
1%
#385220000000
0!
0%
#385225000000
1!
1%
#385230000000
0!
0%
#385235000000
1!
1%
#385240000000
0!
0%
#385245000000
1!
1%
#385250000000
0!
0%
#385255000000
1!
1%
#385260000000
0!
0%
#385265000000
1!
1%
#385270000000
0!
0%
#385275000000
1!
1%
#385280000000
0!
0%
#385285000000
1!
1%
#385290000000
0!
0%
#385295000000
1!
1%
#385300000000
0!
0%
#385305000000
1!
1%
#385310000000
0!
0%
#385315000000
1!
1%
#385320000000
0!
0%
#385325000000
1!
1%
#385330000000
0!
0%
#385335000000
1!
1%
#385340000000
0!
0%
#385345000000
1!
1%
#385350000000
0!
0%
#385355000000
1!
1%
#385360000000
0!
0%
#385365000000
1!
1%
#385370000000
0!
0%
#385375000000
1!
1%
#385380000000
0!
0%
#385385000000
1!
1%
#385390000000
0!
0%
#385395000000
1!
1%
#385400000000
0!
0%
#385405000000
1!
1%
#385410000000
0!
0%
#385415000000
1!
1%
#385420000000
0!
0%
#385425000000
1!
1%
#385430000000
0!
0%
#385435000000
1!
1%
#385440000000
0!
0%
#385445000000
1!
1%
#385450000000
0!
0%
#385455000000
1!
1%
#385460000000
0!
0%
#385465000000
1!
1%
#385470000000
0!
0%
#385475000000
1!
1%
#385480000000
0!
0%
#385485000000
1!
1%
#385490000000
0!
0%
#385495000000
1!
1%
#385500000000
0!
0%
#385505000000
1!
1%
#385510000000
0!
0%
#385515000000
1!
1%
#385520000000
0!
0%
#385525000000
1!
1%
#385530000000
0!
0%
#385535000000
1!
1%
#385540000000
0!
0%
#385545000000
1!
1%
#385550000000
0!
0%
#385555000000
1!
1%
#385560000000
0!
0%
#385565000000
1!
1%
#385570000000
0!
0%
#385575000000
1!
1%
#385580000000
0!
0%
#385585000000
1!
1%
#385590000000
0!
0%
#385595000000
1!
1%
#385600000000
0!
0%
#385605000000
1!
1%
#385610000000
0!
0%
#385615000000
1!
1%
#385620000000
0!
0%
#385625000000
1!
1%
#385630000000
0!
0%
#385635000000
1!
1%
#385640000000
0!
0%
#385645000000
1!
1%
#385650000000
0!
0%
#385655000000
1!
1%
#385660000000
0!
0%
#385665000000
1!
1%
#385670000000
0!
0%
#385675000000
1!
1%
#385680000000
0!
0%
#385685000000
1!
1%
#385690000000
0!
0%
#385695000000
1!
1%
#385700000000
0!
0%
#385705000000
1!
1%
#385710000000
0!
0%
#385715000000
1!
1%
#385720000000
0!
0%
#385725000000
1!
1%
#385730000000
0!
0%
#385735000000
1!
1%
#385740000000
0!
0%
#385745000000
1!
1%
#385750000000
0!
0%
#385755000000
1!
1%
#385760000000
0!
0%
#385765000000
1!
1%
#385770000000
0!
0%
#385775000000
1!
1%
#385780000000
0!
0%
#385785000000
1!
1%
#385790000000
0!
0%
#385795000000
1!
1%
#385800000000
0!
0%
#385805000000
1!
1%
#385810000000
0!
0%
#385815000000
1!
1%
#385820000000
0!
0%
#385825000000
1!
1%
#385830000000
0!
0%
#385835000000
1!
1%
#385840000000
0!
0%
#385845000000
1!
1%
#385850000000
0!
0%
#385855000000
1!
1%
#385860000000
0!
0%
#385865000000
1!
1%
#385870000000
0!
0%
#385875000000
1!
1%
#385880000000
0!
0%
#385885000000
1!
1%
#385890000000
0!
0%
#385895000000
1!
1%
#385900000000
0!
0%
#385905000000
1!
1%
#385910000000
0!
0%
#385915000000
1!
1%
#385920000000
0!
0%
#385925000000
1!
1%
#385930000000
0!
0%
#385935000000
1!
1%
#385940000000
0!
0%
#385945000000
1!
1%
#385950000000
0!
0%
#385955000000
1!
1%
#385960000000
0!
0%
#385965000000
1!
1%
#385970000000
0!
0%
#385975000000
1!
1%
#385980000000
0!
0%
#385985000000
1!
1%
#385990000000
0!
0%
#385995000000
1!
1%
#386000000000
0!
0%
#386005000000
1!
1%
#386010000000
0!
0%
#386015000000
1!
1%
#386020000000
0!
0%
#386025000000
1!
1%
#386030000000
0!
0%
#386035000000
1!
1%
#386040000000
0!
0%
#386045000000
1!
1%
#386050000000
0!
0%
#386055000000
1!
1%
#386060000000
0!
0%
#386065000000
1!
1%
#386070000000
0!
0%
#386075000000
1!
1%
#386080000000
0!
0%
#386085000000
1!
1%
#386090000000
0!
0%
#386095000000
1!
1%
#386100000000
0!
0%
#386105000000
1!
1%
#386110000000
0!
0%
#386115000000
1!
1%
#386120000000
0!
0%
#386125000000
1!
1%
#386130000000
0!
0%
#386135000000
1!
1%
#386140000000
0!
0%
#386145000000
1!
1%
#386150000000
0!
0%
#386155000000
1!
1%
#386160000000
0!
0%
#386165000000
1!
1%
#386170000000
0!
0%
#386175000000
1!
1%
#386180000000
0!
0%
#386185000000
1!
1%
#386190000000
0!
0%
#386195000000
1!
1%
#386200000000
0!
0%
#386205000000
1!
1%
#386210000000
0!
0%
#386215000000
1!
1%
#386220000000
0!
0%
#386225000000
1!
1%
#386230000000
0!
0%
#386235000000
1!
1%
#386240000000
0!
0%
#386245000000
1!
1%
#386250000000
0!
0%
#386255000000
1!
1%
#386260000000
0!
0%
#386265000000
1!
1%
#386270000000
0!
0%
#386275000000
1!
1%
#386280000000
0!
0%
#386285000000
1!
1%
#386290000000
0!
0%
#386295000000
1!
1%
#386300000000
0!
0%
#386305000000
1!
1%
#386310000000
0!
0%
#386315000000
1!
1%
#386320000000
0!
0%
#386325000000
1!
1%
#386330000000
0!
0%
#386335000000
1!
1%
#386340000000
0!
0%
#386345000000
1!
1%
#386350000000
0!
0%
#386355000000
1!
1%
#386360000000
0!
0%
#386365000000
1!
1%
#386370000000
0!
0%
#386375000000
1!
1%
#386380000000
0!
0%
#386385000000
1!
1%
#386390000000
0!
0%
#386395000000
1!
1%
#386400000000
0!
0%
#386405000000
1!
1%
#386410000000
0!
0%
#386415000000
1!
1%
#386420000000
0!
0%
#386425000000
1!
1%
#386430000000
0!
0%
#386435000000
1!
1%
#386440000000
0!
0%
#386445000000
1!
1%
#386450000000
0!
0%
#386455000000
1!
1%
#386460000000
0!
0%
#386465000000
1!
1%
#386470000000
0!
0%
#386475000000
1!
1%
#386480000000
0!
0%
#386485000000
1!
1%
#386490000000
0!
0%
#386495000000
1!
1%
#386500000000
0!
0%
#386505000000
1!
1%
#386510000000
0!
0%
#386515000000
1!
1%
#386520000000
0!
0%
#386525000000
1!
1%
#386530000000
0!
0%
#386535000000
1!
1%
#386540000000
0!
0%
#386545000000
1!
1%
#386550000000
0!
0%
#386555000000
1!
1%
#386560000000
0!
0%
#386565000000
1!
1%
#386570000000
0!
0%
#386575000000
1!
1%
#386580000000
0!
0%
#386585000000
1!
1%
#386590000000
0!
0%
#386595000000
1!
1%
#386600000000
0!
0%
#386605000000
1!
1%
#386610000000
0!
0%
#386615000000
1!
1%
#386620000000
0!
0%
#386625000000
1!
1%
#386630000000
0!
0%
#386635000000
1!
1%
#386640000000
0!
0%
#386645000000
1!
1%
#386650000000
0!
0%
#386655000000
1!
1%
#386660000000
0!
0%
#386665000000
1!
1%
#386670000000
0!
0%
#386675000000
1!
1%
#386680000000
0!
0%
#386685000000
1!
1%
#386690000000
0!
0%
#386695000000
1!
1%
#386700000000
0!
0%
#386705000000
1!
1%
#386710000000
0!
0%
#386715000000
1!
1%
#386720000000
0!
0%
#386725000000
1!
1%
#386730000000
0!
0%
#386735000000
1!
1%
#386740000000
0!
0%
#386745000000
1!
1%
#386750000000
0!
0%
#386755000000
1!
1%
#386760000000
0!
0%
#386765000000
1!
1%
#386770000000
0!
0%
#386775000000
1!
1%
#386780000000
0!
0%
#386785000000
1!
1%
#386790000000
0!
0%
#386795000000
1!
1%
#386800000000
0!
0%
#386805000000
1!
1%
#386810000000
0!
0%
#386815000000
1!
1%
#386820000000
0!
0%
#386825000000
1!
1%
#386830000000
0!
0%
#386835000000
1!
1%
#386840000000
0!
0%
#386845000000
1!
1%
#386850000000
0!
0%
#386855000000
1!
1%
#386860000000
0!
0%
#386865000000
1!
1%
#386870000000
0!
0%
#386875000000
1!
1%
#386880000000
0!
0%
#386885000000
1!
1%
#386890000000
0!
0%
#386895000000
1!
1%
#386900000000
0!
0%
#386905000000
1!
1%
#386910000000
0!
0%
#386915000000
1!
1%
#386920000000
0!
0%
#386925000000
1!
1%
#386930000000
0!
0%
#386935000000
1!
1%
#386940000000
0!
0%
#386945000000
1!
1%
#386950000000
0!
0%
#386955000000
1!
1%
#386960000000
0!
0%
#386965000000
1!
1%
#386970000000
0!
0%
#386975000000
1!
1%
#386980000000
0!
0%
#386985000000
1!
1%
#386990000000
0!
0%
#386995000000
1!
1%
#387000000000
0!
0%
#387005000000
1!
1%
#387010000000
0!
0%
#387015000000
1!
1%
#387020000000
0!
0%
#387025000000
1!
1%
#387030000000
0!
0%
#387035000000
1!
1%
#387040000000
0!
0%
#387045000000
1!
1%
#387050000000
0!
0%
#387055000000
1!
1%
#387060000000
0!
0%
#387065000000
1!
1%
#387070000000
0!
0%
#387075000000
1!
1%
#387080000000
0!
0%
#387085000000
1!
1%
#387090000000
0!
0%
#387095000000
1!
1%
#387100000000
0!
0%
#387105000000
1!
1%
#387110000000
0!
0%
#387115000000
1!
1%
#387120000000
0!
0%
#387125000000
1!
1%
#387130000000
0!
0%
#387135000000
1!
1%
#387140000000
0!
0%
#387145000000
1!
1%
#387150000000
0!
0%
#387155000000
1!
1%
#387160000000
0!
0%
#387165000000
1!
1%
#387170000000
0!
0%
#387175000000
1!
1%
#387180000000
0!
0%
#387185000000
1!
1%
#387190000000
0!
0%
#387195000000
1!
1%
#387200000000
0!
0%
#387205000000
1!
1%
#387210000000
0!
0%
#387215000000
1!
1%
#387220000000
0!
0%
#387225000000
1!
1%
#387230000000
0!
0%
#387235000000
1!
1%
#387240000000
0!
0%
#387245000000
1!
1%
#387250000000
0!
0%
#387255000000
1!
1%
#387260000000
0!
0%
#387265000000
1!
1%
#387270000000
0!
0%
#387275000000
1!
1%
#387280000000
0!
0%
#387285000000
1!
1%
#387290000000
0!
0%
#387295000000
1!
1%
#387300000000
0!
0%
#387305000000
1!
1%
#387310000000
0!
0%
#387315000000
1!
1%
#387320000000
0!
0%
#387325000000
1!
1%
#387330000000
0!
0%
#387335000000
1!
1%
#387340000000
0!
0%
#387345000000
1!
1%
#387350000000
0!
0%
#387355000000
1!
1%
#387360000000
0!
0%
#387365000000
1!
1%
#387370000000
0!
0%
#387375000000
1!
1%
#387380000000
0!
0%
#387385000000
1!
1%
#387390000000
0!
0%
#387395000000
1!
1%
#387400000000
0!
0%
#387405000000
1!
1%
#387410000000
0!
0%
#387415000000
1!
1%
#387420000000
0!
0%
#387425000000
1!
1%
#387430000000
0!
0%
#387435000000
1!
1%
#387440000000
0!
0%
#387445000000
1!
1%
#387450000000
0!
0%
#387455000000
1!
1%
#387460000000
0!
0%
#387465000000
1!
1%
#387470000000
0!
0%
#387475000000
1!
1%
#387480000000
0!
0%
#387485000000
1!
1%
#387490000000
0!
0%
#387495000000
1!
1%
#387500000000
0!
0%
#387505000000
1!
1%
#387510000000
0!
0%
#387515000000
1!
1%
#387520000000
0!
0%
#387525000000
1!
1%
#387530000000
0!
0%
#387535000000
1!
1%
#387540000000
0!
0%
#387545000000
1!
1%
#387550000000
0!
0%
#387555000000
1!
1%
#387560000000
0!
0%
#387565000000
1!
1%
#387570000000
0!
0%
#387575000000
1!
1%
#387580000000
0!
0%
#387585000000
1!
1%
#387590000000
0!
0%
#387595000000
1!
1%
#387600000000
0!
0%
#387605000000
1!
1%
#387610000000
0!
0%
#387615000000
1!
1%
#387620000000
0!
0%
#387625000000
1!
1%
#387630000000
0!
0%
#387635000000
1!
1%
#387640000000
0!
0%
#387645000000
1!
1%
#387650000000
0!
0%
#387655000000
1!
1%
#387660000000
0!
0%
#387665000000
1!
1%
#387670000000
0!
0%
#387675000000
1!
1%
#387680000000
0!
0%
#387685000000
1!
1%
#387690000000
0!
0%
#387695000000
1!
1%
#387700000000
0!
0%
#387705000000
1!
1%
#387710000000
0!
0%
#387715000000
1!
1%
#387720000000
0!
0%
#387725000000
1!
1%
#387730000000
0!
0%
#387735000000
1!
1%
#387740000000
0!
0%
#387745000000
1!
1%
#387750000000
0!
0%
#387755000000
1!
1%
#387760000000
0!
0%
#387765000000
1!
1%
#387770000000
0!
0%
#387775000000
1!
1%
#387780000000
0!
0%
#387785000000
1!
1%
#387790000000
0!
0%
#387795000000
1!
1%
#387800000000
0!
0%
#387805000000
1!
1%
#387810000000
0!
0%
#387815000000
1!
1%
#387820000000
0!
0%
#387825000000
1!
1%
#387830000000
0!
0%
#387835000000
1!
1%
#387840000000
0!
0%
#387845000000
1!
1%
#387850000000
0!
0%
#387855000000
1!
1%
#387860000000
0!
0%
#387865000000
1!
1%
#387870000000
0!
0%
#387875000000
1!
1%
#387880000000
0!
0%
#387885000000
1!
1%
#387890000000
0!
0%
#387895000000
1!
1%
#387900000000
0!
0%
#387905000000
1!
1%
#387910000000
0!
0%
#387915000000
1!
1%
#387920000000
0!
0%
#387925000000
1!
1%
#387930000000
0!
0%
#387935000000
1!
1%
#387940000000
0!
0%
#387945000000
1!
1%
#387950000000
0!
0%
#387955000000
1!
1%
#387960000000
0!
0%
#387965000000
1!
1%
#387970000000
0!
0%
#387975000000
1!
1%
#387980000000
0!
0%
#387985000000
1!
1%
#387990000000
0!
0%
#387995000000
1!
1%
#388000000000
0!
0%
#388005000000
1!
1%
#388010000000
0!
0%
#388015000000
1!
1%
#388020000000
0!
0%
#388025000000
1!
1%
#388030000000
0!
0%
#388035000000
1!
1%
#388040000000
0!
0%
#388045000000
1!
1%
#388050000000
0!
0%
#388055000000
1!
1%
#388060000000
0!
0%
#388065000000
1!
1%
#388070000000
0!
0%
#388075000000
1!
1%
#388080000000
0!
0%
#388085000000
1!
1%
#388090000000
0!
0%
#388095000000
1!
1%
#388100000000
0!
0%
#388105000000
1!
1%
#388110000000
0!
0%
#388115000000
1!
1%
#388120000000
0!
0%
#388125000000
1!
1%
#388130000000
0!
0%
#388135000000
1!
1%
#388140000000
0!
0%
#388145000000
1!
1%
#388150000000
0!
0%
#388155000000
1!
1%
#388160000000
0!
0%
#388165000000
1!
1%
#388170000000
0!
0%
#388175000000
1!
1%
#388180000000
0!
0%
#388185000000
1!
1%
#388190000000
0!
0%
#388195000000
1!
1%
#388200000000
0!
0%
#388205000000
1!
1%
#388210000000
0!
0%
#388215000000
1!
1%
#388220000000
0!
0%
#388225000000
1!
1%
#388230000000
0!
0%
#388235000000
1!
1%
#388240000000
0!
0%
#388245000000
1!
1%
#388250000000
0!
0%
#388255000000
1!
1%
#388260000000
0!
0%
#388265000000
1!
1%
#388270000000
0!
0%
#388275000000
1!
1%
#388280000000
0!
0%
#388285000000
1!
1%
#388290000000
0!
0%
#388295000000
1!
1%
#388300000000
0!
0%
#388305000000
1!
1%
#388310000000
0!
0%
#388315000000
1!
1%
#388320000000
0!
0%
#388325000000
1!
1%
#388330000000
0!
0%
#388335000000
1!
1%
#388340000000
0!
0%
#388345000000
1!
1%
#388350000000
0!
0%
#388355000000
1!
1%
#388360000000
0!
0%
#388365000000
1!
1%
#388370000000
0!
0%
#388375000000
1!
1%
#388380000000
0!
0%
#388385000000
1!
1%
#388390000000
0!
0%
#388395000000
1!
1%
#388400000000
0!
0%
#388405000000
1!
1%
#388410000000
0!
0%
#388415000000
1!
1%
#388420000000
0!
0%
#388425000000
1!
1%
#388430000000
0!
0%
#388435000000
1!
1%
#388440000000
0!
0%
#388445000000
1!
1%
#388450000000
0!
0%
#388455000000
1!
1%
#388460000000
0!
0%
#388465000000
1!
1%
#388470000000
0!
0%
#388475000000
1!
1%
#388480000000
0!
0%
#388485000000
1!
1%
#388490000000
0!
0%
#388495000000
1!
1%
#388500000000
0!
0%
#388505000000
1!
1%
#388510000000
0!
0%
#388515000000
1!
1%
#388520000000
0!
0%
#388525000000
1!
1%
#388530000000
0!
0%
#388535000000
1!
1%
#388540000000
0!
0%
#388545000000
1!
1%
#388550000000
0!
0%
#388555000000
1!
1%
#388560000000
0!
0%
#388565000000
1!
1%
#388570000000
0!
0%
#388575000000
1!
1%
#388580000000
0!
0%
#388585000000
1!
1%
#388590000000
0!
0%
#388595000000
1!
1%
#388600000000
0!
0%
#388605000000
1!
1%
#388610000000
0!
0%
#388615000000
1!
1%
#388620000000
0!
0%
#388625000000
1!
1%
#388630000000
0!
0%
#388635000000
1!
1%
#388640000000
0!
0%
#388645000000
1!
1%
#388650000000
0!
0%
#388655000000
1!
1%
#388660000000
0!
0%
#388665000000
1!
1%
#388670000000
0!
0%
#388675000000
1!
1%
#388680000000
0!
0%
#388685000000
1!
1%
#388690000000
0!
0%
#388695000000
1!
1%
#388700000000
0!
0%
#388705000000
1!
1%
#388710000000
0!
0%
#388715000000
1!
1%
#388720000000
0!
0%
#388725000000
1!
1%
#388730000000
0!
0%
#388735000000
1!
1%
#388740000000
0!
0%
#388745000000
1!
1%
#388750000000
0!
0%
#388755000000
1!
1%
#388760000000
0!
0%
#388765000000
1!
1%
#388770000000
0!
0%
#388775000000
1!
1%
#388780000000
0!
0%
#388785000000
1!
1%
#388790000000
0!
0%
#388795000000
1!
1%
#388800000000
0!
0%
#388805000000
1!
1%
#388810000000
0!
0%
#388815000000
1!
1%
#388820000000
0!
0%
#388825000000
1!
1%
#388830000000
0!
0%
#388835000000
1!
1%
#388840000000
0!
0%
#388845000000
1!
1%
#388850000000
0!
0%
#388855000000
1!
1%
#388860000000
0!
0%
#388865000000
1!
1%
#388870000000
0!
0%
#388875000000
1!
1%
#388880000000
0!
0%
#388885000000
1!
1%
#388890000000
0!
0%
#388895000000
1!
1%
#388900000000
0!
0%
#388905000000
1!
1%
#388910000000
0!
0%
#388915000000
1!
1%
#388920000000
0!
0%
#388925000000
1!
1%
#388930000000
0!
0%
#388935000000
1!
1%
#388940000000
0!
0%
#388945000000
1!
1%
#388950000000
0!
0%
#388955000000
1!
1%
#388960000000
0!
0%
#388965000000
1!
1%
#388970000000
0!
0%
#388975000000
1!
1%
#388980000000
0!
0%
#388985000000
1!
1%
#388990000000
0!
0%
#388995000000
1!
1%
#389000000000
0!
0%
#389005000000
1!
1%
#389010000000
0!
0%
#389015000000
1!
1%
#389020000000
0!
0%
#389025000000
1!
1%
#389030000000
0!
0%
#389035000000
1!
1%
#389040000000
0!
0%
#389045000000
1!
1%
#389050000000
0!
0%
#389055000000
1!
1%
#389060000000
0!
0%
#389065000000
1!
1%
#389070000000
0!
0%
#389075000000
1!
1%
#389080000000
0!
0%
#389085000000
1!
1%
#389090000000
0!
0%
#389095000000
1!
1%
#389100000000
0!
0%
#389105000000
1!
1%
#389110000000
0!
0%
#389115000000
1!
1%
#389120000000
0!
0%
#389125000000
1!
1%
#389130000000
0!
0%
#389135000000
1!
1%
#389140000000
0!
0%
#389145000000
1!
1%
#389150000000
0!
0%
#389155000000
1!
1%
#389160000000
0!
0%
#389165000000
1!
1%
#389170000000
0!
0%
#389175000000
1!
1%
#389180000000
0!
0%
#389185000000
1!
1%
#389190000000
0!
0%
#389195000000
1!
1%
#389200000000
0!
0%
#389205000000
1!
1%
#389210000000
0!
0%
#389215000000
1!
1%
#389220000000
0!
0%
#389225000000
1!
1%
#389230000000
0!
0%
#389235000000
1!
1%
#389240000000
0!
0%
#389245000000
1!
1%
#389250000000
0!
0%
#389255000000
1!
1%
#389260000000
0!
0%
#389265000000
1!
1%
#389270000000
0!
0%
#389275000000
1!
1%
#389280000000
0!
0%
#389285000000
1!
1%
#389290000000
0!
0%
#389295000000
1!
1%
#389300000000
0!
0%
#389305000000
1!
1%
#389310000000
0!
0%
#389315000000
1!
1%
#389320000000
0!
0%
#389325000000
1!
1%
#389330000000
0!
0%
#389335000000
1!
1%
#389340000000
0!
0%
#389345000000
1!
1%
#389350000000
0!
0%
#389355000000
1!
1%
#389360000000
0!
0%
#389365000000
1!
1%
#389370000000
0!
0%
#389375000000
1!
1%
#389380000000
0!
0%
#389385000000
1!
1%
#389390000000
0!
0%
#389395000000
1!
1%
#389400000000
0!
0%
#389405000000
1!
1%
#389410000000
0!
0%
#389415000000
1!
1%
#389420000000
0!
0%
#389425000000
1!
1%
#389430000000
0!
0%
#389435000000
1!
1%
#389440000000
0!
0%
#389445000000
1!
1%
#389450000000
0!
0%
#389455000000
1!
1%
#389460000000
0!
0%
#389465000000
1!
1%
#389470000000
0!
0%
#389475000000
1!
1%
#389480000000
0!
0%
#389485000000
1!
1%
#389490000000
0!
0%
#389495000000
1!
1%
#389500000000
0!
0%
#389505000000
1!
1%
#389510000000
0!
0%
#389515000000
1!
1%
#389520000000
0!
0%
#389525000000
1!
1%
#389530000000
0!
0%
#389535000000
1!
1%
#389540000000
0!
0%
#389545000000
1!
1%
#389550000000
0!
0%
#389555000000
1!
1%
#389560000000
0!
0%
#389565000000
1!
1%
#389570000000
0!
0%
#389575000000
1!
1%
#389580000000
0!
0%
#389585000000
1!
1%
#389590000000
0!
0%
#389595000000
1!
1%
#389600000000
0!
0%
#389605000000
1!
1%
#389610000000
0!
0%
#389615000000
1!
1%
#389620000000
0!
0%
#389625000000
1!
1%
#389630000000
0!
0%
#389635000000
1!
1%
#389640000000
0!
0%
#389645000000
1!
1%
#389650000000
0!
0%
#389655000000
1!
1%
#389660000000
0!
0%
#389665000000
1!
1%
#389670000000
0!
0%
#389675000000
1!
1%
#389680000000
0!
0%
#389685000000
1!
1%
#389690000000
0!
0%
#389695000000
1!
1%
#389700000000
0!
0%
#389705000000
1!
1%
#389710000000
0!
0%
#389715000000
1!
1%
#389720000000
0!
0%
#389725000000
1!
1%
#389730000000
0!
0%
#389735000000
1!
1%
#389740000000
0!
0%
#389745000000
1!
1%
#389750000000
0!
0%
#389755000000
1!
1%
#389760000000
0!
0%
#389765000000
1!
1%
#389770000000
0!
0%
#389775000000
1!
1%
#389780000000
0!
0%
#389785000000
1!
1%
#389790000000
0!
0%
#389795000000
1!
1%
#389800000000
0!
0%
#389805000000
1!
1%
#389810000000
0!
0%
#389815000000
1!
1%
#389820000000
0!
0%
#389825000000
1!
1%
#389830000000
0!
0%
#389835000000
1!
1%
#389840000000
0!
0%
#389845000000
1!
1%
#389850000000
0!
0%
#389855000000
1!
1%
#389860000000
0!
0%
#389865000000
1!
1%
#389870000000
0!
0%
#389875000000
1!
1%
#389880000000
0!
0%
#389885000000
1!
1%
#389890000000
0!
0%
#389895000000
1!
1%
#389900000000
0!
0%
#389905000000
1!
1%
#389910000000
0!
0%
#389915000000
1!
1%
#389920000000
0!
0%
#389925000000
1!
1%
#389930000000
0!
0%
#389935000000
1!
1%
#389940000000
0!
0%
#389945000000
1!
1%
#389950000000
0!
0%
#389955000000
1!
1%
#389960000000
0!
0%
#389965000000
1!
1%
#389970000000
0!
0%
#389975000000
1!
1%
#389980000000
0!
0%
#389985000000
1!
1%
#389990000000
0!
0%
#389995000000
1!
1%
#390000000000
0!
0%
#390005000000
1!
1%
#390010000000
0!
0%
#390015000000
1!
1%
#390020000000
0!
0%
#390025000000
1!
1%
#390030000000
0!
0%
#390035000000
1!
1%
#390040000000
0!
0%
#390045000000
1!
1%
#390050000000
0!
0%
#390055000000
1!
1%
#390060000000
0!
0%
#390065000000
1!
1%
#390070000000
0!
0%
#390075000000
1!
1%
#390080000000
0!
0%
#390085000000
1!
1%
#390090000000
0!
0%
#390095000000
1!
1%
#390100000000
0!
0%
#390105000000
1!
1%
#390110000000
0!
0%
#390115000000
1!
1%
#390120000000
0!
0%
#390125000000
1!
1%
#390130000000
0!
0%
#390135000000
1!
1%
#390140000000
0!
0%
#390145000000
1!
1%
#390150000000
0!
0%
#390155000000
1!
1%
#390160000000
0!
0%
#390165000000
1!
1%
#390170000000
0!
0%
#390175000000
1!
1%
#390180000000
0!
0%
#390185000000
1!
1%
#390190000000
0!
0%
#390195000000
1!
1%
#390200000000
0!
0%
#390205000000
1!
1%
#390210000000
0!
0%
#390215000000
1!
1%
#390220000000
0!
0%
#390225000000
1!
1%
#390230000000
0!
0%
#390235000000
1!
1%
#390240000000
0!
0%
#390245000000
1!
1%
#390250000000
0!
0%
#390255000000
1!
1%
#390260000000
0!
0%
#390265000000
1!
1%
#390270000000
0!
0%
#390275000000
1!
1%
#390280000000
0!
0%
#390285000000
1!
1%
#390290000000
0!
0%
#390295000000
1!
1%
#390300000000
0!
0%
#390305000000
1!
1%
#390310000000
0!
0%
#390315000000
1!
1%
#390320000000
0!
0%
#390325000000
1!
1%
#390330000000
0!
0%
#390335000000
1!
1%
#390340000000
0!
0%
#390345000000
1!
1%
#390350000000
0!
0%
#390355000000
1!
1%
#390360000000
0!
0%
#390365000000
1!
1%
#390370000000
0!
0%
#390375000000
1!
1%
#390380000000
0!
0%
#390385000000
1!
1%
#390390000000
0!
0%
#390395000000
1!
1%
#390400000000
0!
0%
#390405000000
1!
1%
#390410000000
0!
0%
#390415000000
1!
1%
#390420000000
0!
0%
#390425000000
1!
1%
#390430000000
0!
0%
#390435000000
1!
1%
#390440000000
0!
0%
#390445000000
1!
1%
#390450000000
0!
0%
#390455000000
1!
1%
#390460000000
0!
0%
#390465000000
1!
1%
#390470000000
0!
0%
#390475000000
1!
1%
#390480000000
0!
0%
#390485000000
1!
1%
#390490000000
0!
0%
#390495000000
1!
1%
#390500000000
0!
0%
#390505000000
1!
1%
#390510000000
0!
0%
#390515000000
1!
1%
#390520000000
0!
0%
#390525000000
1!
1%
#390530000000
0!
0%
#390535000000
1!
1%
#390540000000
0!
0%
#390545000000
1!
1%
#390550000000
0!
0%
#390555000000
1!
1%
#390560000000
0!
0%
#390565000000
1!
1%
#390570000000
0!
0%
#390575000000
1!
1%
#390580000000
0!
0%
#390585000000
1!
1%
#390590000000
0!
0%
#390595000000
1!
1%
#390600000000
0!
0%
#390605000000
1!
1%
#390610000000
0!
0%
#390615000000
1!
1%
#390620000000
0!
0%
#390625000000
1!
1%
#390630000000
0!
0%
#390635000000
1!
1%
#390640000000
0!
0%
#390645000000
1!
1%
#390650000000
0!
0%
#390655000000
1!
1%
#390660000000
0!
0%
#390665000000
1!
1%
#390670000000
0!
0%
#390675000000
1!
1%
#390680000000
0!
0%
#390685000000
1!
1%
#390690000000
0!
0%
#390695000000
1!
1%
#390700000000
0!
0%
#390705000000
1!
1%
#390710000000
0!
0%
#390715000000
1!
1%
#390720000000
0!
0%
#390725000000
1!
1%
#390730000000
0!
0%
#390735000000
1!
1%
#390740000000
0!
0%
#390745000000
1!
1%
#390750000000
0!
0%
#390755000000
1!
1%
#390760000000
0!
0%
#390765000000
1!
1%
#390770000000
0!
0%
#390775000000
1!
1%
#390780000000
0!
0%
#390785000000
1!
1%
#390790000000
0!
0%
#390795000000
1!
1%
#390800000000
0!
0%
#390805000000
1!
1%
#390810000000
0!
0%
#390815000000
1!
1%
#390820000000
0!
0%
#390825000000
1!
1%
#390830000000
0!
0%
#390835000000
1!
1%
#390840000000
0!
0%
#390845000000
1!
1%
#390850000000
0!
0%
#390855000000
1!
1%
#390860000000
0!
0%
#390865000000
1!
1%
#390870000000
0!
0%
#390875000000
1!
1%
#390880000000
0!
0%
#390885000000
1!
1%
#390890000000
0!
0%
#390895000000
1!
1%
#390900000000
0!
0%
#390905000000
1!
1%
#390910000000
0!
0%
#390915000000
1!
1%
#390920000000
0!
0%
#390925000000
1!
1%
#390930000000
0!
0%
#390935000000
1!
1%
#390940000000
0!
0%
#390945000000
1!
1%
#390950000000
0!
0%
#390955000000
1!
1%
#390960000000
0!
0%
#390965000000
1!
1%
#390970000000
0!
0%
#390975000000
1!
1%
#390980000000
0!
0%
#390985000000
1!
1%
#390990000000
0!
0%
#390995000000
1!
1%
#391000000000
0!
0%
#391005000000
1!
1%
#391010000000
0!
0%
#391015000000
1!
1%
#391020000000
0!
0%
#391025000000
1!
1%
#391030000000
0!
0%
#391035000000
1!
1%
#391040000000
0!
0%
#391045000000
1!
1%
#391050000000
0!
0%
#391055000000
1!
1%
#391060000000
0!
0%
#391065000000
1!
1%
#391070000000
0!
0%
#391075000000
1!
1%
#391080000000
0!
0%
#391085000000
1!
1%
#391090000000
0!
0%
#391095000000
1!
1%
#391100000000
0!
0%
#391105000000
1!
1%
#391110000000
0!
0%
#391115000000
1!
1%
#391120000000
0!
0%
#391125000000
1!
1%
#391130000000
0!
0%
#391135000000
1!
1%
#391140000000
0!
0%
#391145000000
1!
1%
#391150000000
0!
0%
#391155000000
1!
1%
#391160000000
0!
0%
#391165000000
1!
1%
#391170000000
0!
0%
#391175000000
1!
1%
#391180000000
0!
0%
#391185000000
1!
1%
#391190000000
0!
0%
#391195000000
1!
1%
#391200000000
0!
0%
#391205000000
1!
1%
#391210000000
0!
0%
#391215000000
1!
1%
#391220000000
0!
0%
#391225000000
1!
1%
#391230000000
0!
0%
#391235000000
1!
1%
#391240000000
0!
0%
#391245000000
1!
1%
#391250000000
0!
0%
#391255000000
1!
1%
#391260000000
0!
0%
#391265000000
1!
1%
#391270000000
0!
0%
#391275000000
1!
1%
#391280000000
0!
0%
#391285000000
1!
1%
#391290000000
0!
0%
#391295000000
1!
1%
#391300000000
0!
0%
#391305000000
1!
1%
#391310000000
0!
0%
#391315000000
1!
1%
#391320000000
0!
0%
#391325000000
1!
1%
#391330000000
0!
0%
#391335000000
1!
1%
#391340000000
0!
0%
#391345000000
1!
1%
#391350000000
0!
0%
#391355000000
1!
1%
#391360000000
0!
0%
#391365000000
1!
1%
#391370000000
0!
0%
#391375000000
1!
1%
#391380000000
0!
0%
#391385000000
1!
1%
#391390000000
0!
0%
#391395000000
1!
1%
#391400000000
0!
0%
#391405000000
1!
1%
#391410000000
0!
0%
#391415000000
1!
1%
#391420000000
0!
0%
#391425000000
1!
1%
#391430000000
0!
0%
#391435000000
1!
1%
#391440000000
0!
0%
#391445000000
1!
1%
#391450000000
0!
0%
#391455000000
1!
1%
#391460000000
0!
0%
#391465000000
1!
1%
#391470000000
0!
0%
#391475000000
1!
1%
#391480000000
0!
0%
#391485000000
1!
1%
#391490000000
0!
0%
#391495000000
1!
1%
#391500000000
0!
0%
#391505000000
1!
1%
#391510000000
0!
0%
#391515000000
1!
1%
#391520000000
0!
0%
#391525000000
1!
1%
#391530000000
0!
0%
#391535000000
1!
1%
#391540000000
0!
0%
#391545000000
1!
1%
#391550000000
0!
0%
#391555000000
1!
1%
#391560000000
0!
0%
#391565000000
1!
1%
#391570000000
0!
0%
#391575000000
1!
1%
#391580000000
0!
0%
#391585000000
1!
1%
#391590000000
0!
0%
#391595000000
1!
1%
#391600000000
0!
0%
#391605000000
1!
1%
#391610000000
0!
0%
#391615000000
1!
1%
#391620000000
0!
0%
#391625000000
1!
1%
#391630000000
0!
0%
#391635000000
1!
1%
#391640000000
0!
0%
#391645000000
1!
1%
#391650000000
0!
0%
#391655000000
1!
1%
#391660000000
0!
0%
#391665000000
1!
1%
#391670000000
0!
0%
#391675000000
1!
1%
#391680000000
0!
0%
#391685000000
1!
1%
#391690000000
0!
0%
#391695000000
1!
1%
#391700000000
0!
0%
#391705000000
1!
1%
#391710000000
0!
0%
#391715000000
1!
1%
#391720000000
0!
0%
#391725000000
1!
1%
#391730000000
0!
0%
#391735000000
1!
1%
#391740000000
0!
0%
#391745000000
1!
1%
#391750000000
0!
0%
#391755000000
1!
1%
#391760000000
0!
0%
#391765000000
1!
1%
#391770000000
0!
0%
#391775000000
1!
1%
#391780000000
0!
0%
#391785000000
1!
1%
#391790000000
0!
0%
#391795000000
1!
1%
#391800000000
0!
0%
#391805000000
1!
1%
#391810000000
0!
0%
#391815000000
1!
1%
#391820000000
0!
0%
#391825000000
1!
1%
#391830000000
0!
0%
#391835000000
1!
1%
#391840000000
0!
0%
#391845000000
1!
1%
#391850000000
0!
0%
#391855000000
1!
1%
#391860000000
0!
0%
#391865000000
1!
1%
#391870000000
0!
0%
#391875000000
1!
1%
#391880000000
0!
0%
#391885000000
1!
1%
#391890000000
0!
0%
#391895000000
1!
1%
#391900000000
0!
0%
#391905000000
1!
1%
#391910000000
0!
0%
#391915000000
1!
1%
#391920000000
0!
0%
#391925000000
1!
1%
#391930000000
0!
0%
#391935000000
1!
1%
#391940000000
0!
0%
#391945000000
1!
1%
#391950000000
0!
0%
#391955000000
1!
1%
#391960000000
0!
0%
#391965000000
1!
1%
#391970000000
0!
0%
#391975000000
1!
1%
#391980000000
0!
0%
#391985000000
1!
1%
#391990000000
0!
0%
#391995000000
1!
1%
#392000000000
0!
0%
#392005000000
1!
1%
#392010000000
0!
0%
#392015000000
1!
1%
#392020000000
0!
0%
#392025000000
1!
1%
#392030000000
0!
0%
#392035000000
1!
1%
#392040000000
0!
0%
#392045000000
1!
1%
#392050000000
0!
0%
#392055000000
1!
1%
#392060000000
0!
0%
#392065000000
1!
1%
#392070000000
0!
0%
#392075000000
1!
1%
#392080000000
0!
0%
#392085000000
1!
1%
#392090000000
0!
0%
#392095000000
1!
1%
#392100000000
0!
0%
#392105000000
1!
1%
#392110000000
0!
0%
#392115000000
1!
1%
#392120000000
0!
0%
#392125000000
1!
1%
#392130000000
0!
0%
#392135000000
1!
1%
#392140000000
0!
0%
#392145000000
1!
1%
#392150000000
0!
0%
#392155000000
1!
1%
#392160000000
0!
0%
#392165000000
1!
1%
#392170000000
0!
0%
#392175000000
1!
1%
#392180000000
0!
0%
#392185000000
1!
1%
#392190000000
0!
0%
#392195000000
1!
1%
#392200000000
0!
0%
#392205000000
1!
1%
#392210000000
0!
0%
#392215000000
1!
1%
#392220000000
0!
0%
#392225000000
1!
1%
#392230000000
0!
0%
#392235000000
1!
1%
#392240000000
0!
0%
#392245000000
1!
1%
#392250000000
0!
0%
#392255000000
1!
1%
#392260000000
0!
0%
#392265000000
1!
1%
#392270000000
0!
0%
#392275000000
1!
1%
#392280000000
0!
0%
#392285000000
1!
1%
#392290000000
0!
0%
#392295000000
1!
1%
#392300000000
0!
0%
#392305000000
1!
1%
#392310000000
0!
0%
#392315000000
1!
1%
#392320000000
0!
0%
#392325000000
1!
1%
#392330000000
0!
0%
#392335000000
1!
1%
#392340000000
0!
0%
#392345000000
1!
1%
#392350000000
0!
0%
#392355000000
1!
1%
#392360000000
0!
0%
#392365000000
1!
1%
#392370000000
0!
0%
#392375000000
1!
1%
#392380000000
0!
0%
#392385000000
1!
1%
#392390000000
0!
0%
#392395000000
1!
1%
#392400000000
0!
0%
#392405000000
1!
1%
#392410000000
0!
0%
#392415000000
1!
1%
#392420000000
0!
0%
#392425000000
1!
1%
#392430000000
0!
0%
#392435000000
1!
1%
#392440000000
0!
0%
#392445000000
1!
1%
#392450000000
0!
0%
#392455000000
1!
1%
#392460000000
0!
0%
#392465000000
1!
1%
#392470000000
0!
0%
#392475000000
1!
1%
#392480000000
0!
0%
#392485000000
1!
1%
#392490000000
0!
0%
#392495000000
1!
1%
#392500000000
0!
0%
#392505000000
1!
1%
#392510000000
0!
0%
#392515000000
1!
1%
#392520000000
0!
0%
#392525000000
1!
1%
#392530000000
0!
0%
#392535000000
1!
1%
#392540000000
0!
0%
#392545000000
1!
1%
#392550000000
0!
0%
#392555000000
1!
1%
#392560000000
0!
0%
#392565000000
1!
1%
#392570000000
0!
0%
#392575000000
1!
1%
#392580000000
0!
0%
#392585000000
1!
1%
#392590000000
0!
0%
#392595000000
1!
1%
#392600000000
0!
0%
#392605000000
1!
1%
#392610000000
0!
0%
#392615000000
1!
1%
#392620000000
0!
0%
#392625000000
1!
1%
#392630000000
0!
0%
#392635000000
1!
1%
#392640000000
0!
0%
#392645000000
1!
1%
#392650000000
0!
0%
#392655000000
1!
1%
#392660000000
0!
0%
#392665000000
1!
1%
#392670000000
0!
0%
#392675000000
1!
1%
#392680000000
0!
0%
#392685000000
1!
1%
#392690000000
0!
0%
#392695000000
1!
1%
#392700000000
0!
0%
#392705000000
1!
1%
#392710000000
0!
0%
#392715000000
1!
1%
#392720000000
0!
0%
#392725000000
1!
1%
#392730000000
0!
0%
#392735000000
1!
1%
#392740000000
0!
0%
#392745000000
1!
1%
#392750000000
0!
0%
#392755000000
1!
1%
#392760000000
0!
0%
#392765000000
1!
1%
#392770000000
0!
0%
#392775000000
1!
1%
#392780000000
0!
0%
#392785000000
1!
1%
#392790000000
0!
0%
#392795000000
1!
1%
#392800000000
0!
0%
#392805000000
1!
1%
#392810000000
0!
0%
#392815000000
1!
1%
#392820000000
0!
0%
#392825000000
1!
1%
#392830000000
0!
0%
#392835000000
1!
1%
#392840000000
0!
0%
#392845000000
1!
1%
#392850000000
0!
0%
#392855000000
1!
1%
#392860000000
0!
0%
#392865000000
1!
1%
#392870000000
0!
0%
#392875000000
1!
1%
#392880000000
0!
0%
#392885000000
1!
1%
#392890000000
0!
0%
#392895000000
1!
1%
#392900000000
0!
0%
#392905000000
1!
1%
#392910000000
0!
0%
#392915000000
1!
1%
#392920000000
0!
0%
#392925000000
1!
1%
#392930000000
0!
0%
#392935000000
1!
1%
#392940000000
0!
0%
#392945000000
1!
1%
#392950000000
0!
0%
#392955000000
1!
1%
#392960000000
0!
0%
#392965000000
1!
1%
#392970000000
0!
0%
#392975000000
1!
1%
#392980000000
0!
0%
#392985000000
1!
1%
#392990000000
0!
0%
#392995000000
1!
1%
#393000000000
0!
0%
#393005000000
1!
1%
#393010000000
0!
0%
#393015000000
1!
1%
#393020000000
0!
0%
#393025000000
1!
1%
#393030000000
0!
0%
#393035000000
1!
1%
#393040000000
0!
0%
#393045000000
1!
1%
#393050000000
0!
0%
#393055000000
1!
1%
#393060000000
0!
0%
#393065000000
1!
1%
#393070000000
0!
0%
#393075000000
1!
1%
#393080000000
0!
0%
#393085000000
1!
1%
#393090000000
0!
0%
#393095000000
1!
1%
#393100000000
0!
0%
#393105000000
1!
1%
#393110000000
0!
0%
#393115000000
1!
1%
#393120000000
0!
0%
#393125000000
1!
1%
#393130000000
0!
0%
#393135000000
1!
1%
#393140000000
0!
0%
#393145000000
1!
1%
#393150000000
0!
0%
#393155000000
1!
1%
#393160000000
0!
0%
#393165000000
1!
1%
#393170000000
0!
0%
#393175000000
1!
1%
#393180000000
0!
0%
#393185000000
1!
1%
#393190000000
0!
0%
#393195000000
1!
1%
#393200000000
0!
0%
#393205000000
1!
1%
#393210000000
0!
0%
#393215000000
1!
1%
#393220000000
0!
0%
#393225000000
1!
1%
#393230000000
0!
0%
#393235000000
1!
1%
#393240000000
0!
0%
#393245000000
1!
1%
#393250000000
0!
0%
#393255000000
1!
1%
#393260000000
0!
0%
#393265000000
1!
1%
#393270000000
0!
0%
#393275000000
1!
1%
#393280000000
0!
0%
#393285000000
1!
1%
#393290000000
0!
0%
#393295000000
1!
1%
#393300000000
0!
0%
#393305000000
1!
1%
#393310000000
0!
0%
#393315000000
1!
1%
#393320000000
0!
0%
#393325000000
1!
1%
#393330000000
0!
0%
#393335000000
1!
1%
#393340000000
0!
0%
#393345000000
1!
1%
#393350000000
0!
0%
#393355000000
1!
1%
#393360000000
0!
0%
#393365000000
1!
1%
#393370000000
0!
0%
#393375000000
1!
1%
#393380000000
0!
0%
#393385000000
1!
1%
#393390000000
0!
0%
#393395000000
1!
1%
#393400000000
0!
0%
#393405000000
1!
1%
#393410000000
0!
0%
#393415000000
1!
1%
#393420000000
0!
0%
#393425000000
1!
1%
#393430000000
0!
0%
#393435000000
1!
1%
#393440000000
0!
0%
#393445000000
1!
1%
#393450000000
0!
0%
#393455000000
1!
1%
#393460000000
0!
0%
#393465000000
1!
1%
#393470000000
0!
0%
#393475000000
1!
1%
#393480000000
0!
0%
#393485000000
1!
1%
#393490000000
0!
0%
#393495000000
1!
1%
#393500000000
0!
0%
#393505000000
1!
1%
#393510000000
0!
0%
#393515000000
1!
1%
#393520000000
0!
0%
#393525000000
1!
1%
#393530000000
0!
0%
#393535000000
1!
1%
#393540000000
0!
0%
#393545000000
1!
1%
#393550000000
0!
0%
#393555000000
1!
1%
#393560000000
0!
0%
#393565000000
1!
1%
#393570000000
0!
0%
#393575000000
1!
1%
#393580000000
0!
0%
#393585000000
1!
1%
#393590000000
0!
0%
#393595000000
1!
1%
#393600000000
0!
0%
#393605000000
1!
1%
#393610000000
0!
0%
#393615000000
1!
1%
#393620000000
0!
0%
#393625000000
1!
1%
#393630000000
0!
0%
#393635000000
1!
1%
#393640000000
0!
0%
#393645000000
1!
1%
#393650000000
0!
0%
#393655000000
1!
1%
#393660000000
0!
0%
#393665000000
1!
1%
#393670000000
0!
0%
#393675000000
1!
1%
#393680000000
0!
0%
#393685000000
1!
1%
#393690000000
0!
0%
#393695000000
1!
1%
#393700000000
0!
0%
#393705000000
1!
1%
#393710000000
0!
0%
#393715000000
1!
1%
#393720000000
0!
0%
#393725000000
1!
1%
#393730000000
0!
0%
#393735000000
1!
1%
#393740000000
0!
0%
#393745000000
1!
1%
#393750000000
0!
0%
#393755000000
1!
1%
#393760000000
0!
0%
#393765000000
1!
1%
#393770000000
0!
0%
#393775000000
1!
1%
#393780000000
0!
0%
#393785000000
1!
1%
#393790000000
0!
0%
#393795000000
1!
1%
#393800000000
0!
0%
#393805000000
1!
1%
#393810000000
0!
0%
#393815000000
1!
1%
#393820000000
0!
0%
#393825000000
1!
1%
#393830000000
0!
0%
#393835000000
1!
1%
#393840000000
0!
0%
#393845000000
1!
1%
#393850000000
0!
0%
#393855000000
1!
1%
#393860000000
0!
0%
#393865000000
1!
1%
#393870000000
0!
0%
#393875000000
1!
1%
#393880000000
0!
0%
#393885000000
1!
1%
#393890000000
0!
0%
#393895000000
1!
1%
#393900000000
0!
0%
#393905000000
1!
1%
#393910000000
0!
0%
#393915000000
1!
1%
#393920000000
0!
0%
#393925000000
1!
1%
#393930000000
0!
0%
#393935000000
1!
1%
#393940000000
0!
0%
#393945000000
1!
1%
#393950000000
0!
0%
#393955000000
1!
1%
#393960000000
0!
0%
#393965000000
1!
1%
#393970000000
0!
0%
#393975000000
1!
1%
#393980000000
0!
0%
#393985000000
1!
1%
#393990000000
0!
0%
#393995000000
1!
1%
#394000000000
0!
0%
#394005000000
1!
1%
#394010000000
0!
0%
#394015000000
1!
1%
#394020000000
0!
0%
#394025000000
1!
1%
#394030000000
0!
0%
#394035000000
1!
1%
#394040000000
0!
0%
#394045000000
1!
1%
#394050000000
0!
0%
#394055000000
1!
1%
#394060000000
0!
0%
#394065000000
1!
1%
#394070000000
0!
0%
#394075000000
1!
1%
#394080000000
0!
0%
#394085000000
1!
1%
#394090000000
0!
0%
#394095000000
1!
1%
#394100000000
0!
0%
#394105000000
1!
1%
#394110000000
0!
0%
#394115000000
1!
1%
#394120000000
0!
0%
#394125000000
1!
1%
#394130000000
0!
0%
#394135000000
1!
1%
#394140000000
0!
0%
#394145000000
1!
1%
#394150000000
0!
0%
#394155000000
1!
1%
#394160000000
0!
0%
#394165000000
1!
1%
#394170000000
0!
0%
#394175000000
1!
1%
#394180000000
0!
0%
#394185000000
1!
1%
#394190000000
0!
0%
#394195000000
1!
1%
#394200000000
0!
0%
#394205000000
1!
1%
#394210000000
0!
0%
#394215000000
1!
1%
#394220000000
0!
0%
#394225000000
1!
1%
#394230000000
0!
0%
#394235000000
1!
1%
#394240000000
0!
0%
#394245000000
1!
1%
#394250000000
0!
0%
#394255000000
1!
1%
#394260000000
0!
0%
#394265000000
1!
1%
#394270000000
0!
0%
#394275000000
1!
1%
#394280000000
0!
0%
#394285000000
1!
1%
#394290000000
0!
0%
#394295000000
1!
1%
#394300000000
0!
0%
#394305000000
1!
1%
#394310000000
0!
0%
#394315000000
1!
1%
#394320000000
0!
0%
#394325000000
1!
1%
#394330000000
0!
0%
#394335000000
1!
1%
#394340000000
0!
0%
#394345000000
1!
1%
#394350000000
0!
0%
#394355000000
1!
1%
#394360000000
0!
0%
#394365000000
1!
1%
#394370000000
0!
0%
#394375000000
1!
1%
#394380000000
0!
0%
#394385000000
1!
1%
#394390000000
0!
0%
#394395000000
1!
1%
#394400000000
0!
0%
#394405000000
1!
1%
#394410000000
0!
0%
#394415000000
1!
1%
#394420000000
0!
0%
#394425000000
1!
1%
#394430000000
0!
0%
#394435000000
1!
1%
#394440000000
0!
0%
#394445000000
1!
1%
#394450000000
0!
0%
#394455000000
1!
1%
#394460000000
0!
0%
#394465000000
1!
1%
#394470000000
0!
0%
#394475000000
1!
1%
#394480000000
0!
0%
#394485000000
1!
1%
#394490000000
0!
0%
#394495000000
1!
1%
#394500000000
0!
0%
#394505000000
1!
1%
#394510000000
0!
0%
#394515000000
1!
1%
#394520000000
0!
0%
#394525000000
1!
1%
#394530000000
0!
0%
#394535000000
1!
1%
#394540000000
0!
0%
#394545000000
1!
1%
#394550000000
0!
0%
#394555000000
1!
1%
#394560000000
0!
0%
#394565000000
1!
1%
#394570000000
0!
0%
#394575000000
1!
1%
#394580000000
0!
0%
#394585000000
1!
1%
#394590000000
0!
0%
#394595000000
1!
1%
#394600000000
0!
0%
#394605000000
1!
1%
#394610000000
0!
0%
#394615000000
1!
1%
#394620000000
0!
0%
#394625000000
1!
1%
#394630000000
0!
0%
#394635000000
1!
1%
#394640000000
0!
0%
#394645000000
1!
1%
#394650000000
0!
0%
#394655000000
1!
1%
#394660000000
0!
0%
#394665000000
1!
1%
#394670000000
0!
0%
#394675000000
1!
1%
#394680000000
0!
0%
#394685000000
1!
1%
#394690000000
0!
0%
#394695000000
1!
1%
#394700000000
0!
0%
#394705000000
1!
1%
#394710000000
0!
0%
#394715000000
1!
1%
#394720000000
0!
0%
#394725000000
1!
1%
#394730000000
0!
0%
#394735000000
1!
1%
#394740000000
0!
0%
#394745000000
1!
1%
#394750000000
0!
0%
#394755000000
1!
1%
#394760000000
0!
0%
#394765000000
1!
1%
#394770000000
0!
0%
#394775000000
1!
1%
#394780000000
0!
0%
#394785000000
1!
1%
#394790000000
0!
0%
#394795000000
1!
1%
#394800000000
0!
0%
#394805000000
1!
1%
#394810000000
0!
0%
#394815000000
1!
1%
#394820000000
0!
0%
#394825000000
1!
1%
#394830000000
0!
0%
#394835000000
1!
1%
#394840000000
0!
0%
#394845000000
1!
1%
#394850000000
0!
0%
#394855000000
1!
1%
#394860000000
0!
0%
#394865000000
1!
1%
#394870000000
0!
0%
#394875000000
1!
1%
#394880000000
0!
0%
#394885000000
1!
1%
#394890000000
0!
0%
#394895000000
1!
1%
#394900000000
0!
0%
#394905000000
1!
1%
#394910000000
0!
0%
#394915000000
1!
1%
#394920000000
0!
0%
#394925000000
1!
1%
#394930000000
0!
0%
#394935000000
1!
1%
#394940000000
0!
0%
#394945000000
1!
1%
#394950000000
0!
0%
#394955000000
1!
1%
#394960000000
0!
0%
#394965000000
1!
1%
#394970000000
0!
0%
#394975000000
1!
1%
#394980000000
0!
0%
#394985000000
1!
1%
#394990000000
0!
0%
#394995000000
1!
1%
#395000000000
0!
0%
#395005000000
1!
1%
#395010000000
0!
0%
#395015000000
1!
1%
#395020000000
0!
0%
#395025000000
1!
1%
#395030000000
0!
0%
#395035000000
1!
1%
#395040000000
0!
0%
#395045000000
1!
1%
#395050000000
0!
0%
#395055000000
1!
1%
#395060000000
0!
0%
#395065000000
1!
1%
#395070000000
0!
0%
#395075000000
1!
1%
#395080000000
0!
0%
#395085000000
1!
1%
#395090000000
0!
0%
#395095000000
1!
1%
#395100000000
0!
0%
#395105000000
1!
1%
#395110000000
0!
0%
#395115000000
1!
1%
#395120000000
0!
0%
#395125000000
1!
1%
#395130000000
0!
0%
#395135000000
1!
1%
#395140000000
0!
0%
#395145000000
1!
1%
#395150000000
0!
0%
#395155000000
1!
1%
#395160000000
0!
0%
#395165000000
1!
1%
#395170000000
0!
0%
#395175000000
1!
1%
#395180000000
0!
0%
#395185000000
1!
1%
#395190000000
0!
0%
#395195000000
1!
1%
#395200000000
0!
0%
#395205000000
1!
1%
#395210000000
0!
0%
#395215000000
1!
1%
#395220000000
0!
0%
#395225000000
1!
1%
#395230000000
0!
0%
#395235000000
1!
1%
#395240000000
0!
0%
#395245000000
1!
1%
#395250000000
0!
0%
#395255000000
1!
1%
#395260000000
0!
0%
#395265000000
1!
1%
#395270000000
0!
0%
#395275000000
1!
1%
#395280000000
0!
0%
#395285000000
1!
1%
#395290000000
0!
0%
#395295000000
1!
1%
#395300000000
0!
0%
#395305000000
1!
1%
#395310000000
0!
0%
#395315000000
1!
1%
#395320000000
0!
0%
#395325000000
1!
1%
#395330000000
0!
0%
#395335000000
1!
1%
#395340000000
0!
0%
#395345000000
1!
1%
#395350000000
0!
0%
#395355000000
1!
1%
#395360000000
0!
0%
#395365000000
1!
1%
#395370000000
0!
0%
#395375000000
1!
1%
#395380000000
0!
0%
#395385000000
1!
1%
#395390000000
0!
0%
#395395000000
1!
1%
#395400000000
0!
0%
#395405000000
1!
1%
#395410000000
0!
0%
#395415000000
1!
1%
#395420000000
0!
0%
#395425000000
1!
1%
#395430000000
0!
0%
#395435000000
1!
1%
#395440000000
0!
0%
#395445000000
1!
1%
#395450000000
0!
0%
#395455000000
1!
1%
#395460000000
0!
0%
#395465000000
1!
1%
#395470000000
0!
0%
#395475000000
1!
1%
#395480000000
0!
0%
#395485000000
1!
1%
#395490000000
0!
0%
#395495000000
1!
1%
#395500000000
0!
0%
#395505000000
1!
1%
#395510000000
0!
0%
#395515000000
1!
1%
#395520000000
0!
0%
#395525000000
1!
1%
#395530000000
0!
0%
#395535000000
1!
1%
#395540000000
0!
0%
#395545000000
1!
1%
#395550000000
0!
0%
#395555000000
1!
1%
#395560000000
0!
0%
#395565000000
1!
1%
#395570000000
0!
0%
#395575000000
1!
1%
#395580000000
0!
0%
#395585000000
1!
1%
#395590000000
0!
0%
#395595000000
1!
1%
#395600000000
0!
0%
#395605000000
1!
1%
#395610000000
0!
0%
#395615000000
1!
1%
#395620000000
0!
0%
#395625000000
1!
1%
#395630000000
0!
0%
#395635000000
1!
1%
#395640000000
0!
0%
#395645000000
1!
1%
#395650000000
0!
0%
#395655000000
1!
1%
#395660000000
0!
0%
#395665000000
1!
1%
#395670000000
0!
0%
#395675000000
1!
1%
#395680000000
0!
0%
#395685000000
1!
1%
#395690000000
0!
0%
#395695000000
1!
1%
#395700000000
0!
0%
#395705000000
1!
1%
#395710000000
0!
0%
#395715000000
1!
1%
#395720000000
0!
0%
#395725000000
1!
1%
#395730000000
0!
0%
#395735000000
1!
1%
#395740000000
0!
0%
#395745000000
1!
1%
#395750000000
0!
0%
#395755000000
1!
1%
#395760000000
0!
0%
#395765000000
1!
1%
#395770000000
0!
0%
#395775000000
1!
1%
#395780000000
0!
0%
#395785000000
1!
1%
#395790000000
0!
0%
#395795000000
1!
1%
#395800000000
0!
0%
#395805000000
1!
1%
#395810000000
0!
0%
#395815000000
1!
1%
#395820000000
0!
0%
#395825000000
1!
1%
#395830000000
0!
0%
#395835000000
1!
1%
#395840000000
0!
0%
#395845000000
1!
1%
#395850000000
0!
0%
#395855000000
1!
1%
#395860000000
0!
0%
#395865000000
1!
1%
#395870000000
0!
0%
#395875000000
1!
1%
#395880000000
0!
0%
#395885000000
1!
1%
#395890000000
0!
0%
#395895000000
1!
1%
#395900000000
0!
0%
#395905000000
1!
1%
#395910000000
0!
0%
#395915000000
1!
1%
#395920000000
0!
0%
#395925000000
1!
1%
#395930000000
0!
0%
#395935000000
1!
1%
#395940000000
0!
0%
#395945000000
1!
1%
#395950000000
0!
0%
#395955000000
1!
1%
#395960000000
0!
0%
#395965000000
1!
1%
#395970000000
0!
0%
#395975000000
1!
1%
#395980000000
0!
0%
#395985000000
1!
1%
#395990000000
0!
0%
#395995000000
1!
1%
#396000000000
0!
0%
#396005000000
1!
1%
#396010000000
0!
0%
#396015000000
1!
1%
#396020000000
0!
0%
#396025000000
1!
1%
#396030000000
0!
0%
#396035000000
1!
1%
#396040000000
0!
0%
#396045000000
1!
1%
#396050000000
0!
0%
#396055000000
1!
1%
#396060000000
0!
0%
#396065000000
1!
1%
#396070000000
0!
0%
#396075000000
1!
1%
#396080000000
0!
0%
#396085000000
1!
1%
#396090000000
0!
0%
#396095000000
1!
1%
#396100000000
0!
0%
#396105000000
1!
1%
#396110000000
0!
0%
#396115000000
1!
1%
#396120000000
0!
0%
#396125000000
1!
1%
#396130000000
0!
0%
#396135000000
1!
1%
#396140000000
0!
0%
#396145000000
1!
1%
#396150000000
0!
0%
#396155000000
1!
1%
#396160000000
0!
0%
#396165000000
1!
1%
#396170000000
0!
0%
#396175000000
1!
1%
#396180000000
0!
0%
#396185000000
1!
1%
#396190000000
0!
0%
#396195000000
1!
1%
#396200000000
0!
0%
#396205000000
1!
1%
#396210000000
0!
0%
#396215000000
1!
1%
#396220000000
0!
0%
#396225000000
1!
1%
#396230000000
0!
0%
#396235000000
1!
1%
#396240000000
0!
0%
#396245000000
1!
1%
#396250000000
0!
0%
#396255000000
1!
1%
#396260000000
0!
0%
#396265000000
1!
1%
#396270000000
0!
0%
#396275000000
1!
1%
#396280000000
0!
0%
#396285000000
1!
1%
#396290000000
0!
0%
#396295000000
1!
1%
#396300000000
0!
0%
#396305000000
1!
1%
#396310000000
0!
0%
#396315000000
1!
1%
#396320000000
0!
0%
#396325000000
1!
1%
#396330000000
0!
0%
#396335000000
1!
1%
#396340000000
0!
0%
#396345000000
1!
1%
#396350000000
0!
0%
#396355000000
1!
1%
#396360000000
0!
0%
#396365000000
1!
1%
#396370000000
0!
0%
#396375000000
1!
1%
#396380000000
0!
0%
#396385000000
1!
1%
#396390000000
0!
0%
#396395000000
1!
1%
#396400000000
0!
0%
#396405000000
1!
1%
#396410000000
0!
0%
#396415000000
1!
1%
#396420000000
0!
0%
#396425000000
1!
1%
#396430000000
0!
0%
#396435000000
1!
1%
#396440000000
0!
0%
#396445000000
1!
1%
#396450000000
0!
0%
#396455000000
1!
1%
#396460000000
0!
0%
#396465000000
1!
1%
#396470000000
0!
0%
#396475000000
1!
1%
#396480000000
0!
0%
#396485000000
1!
1%
#396490000000
0!
0%
#396495000000
1!
1%
#396500000000
0!
0%
#396505000000
1!
1%
#396510000000
0!
0%
#396515000000
1!
1%
#396520000000
0!
0%
#396525000000
1!
1%
#396530000000
0!
0%
#396535000000
1!
1%
#396540000000
0!
0%
#396545000000
1!
1%
#396550000000
0!
0%
#396555000000
1!
1%
#396560000000
0!
0%
#396565000000
1!
1%
#396570000000
0!
0%
#396575000000
1!
1%
#396580000000
0!
0%
#396585000000
1!
1%
#396590000000
0!
0%
#396595000000
1!
1%
#396600000000
0!
0%
#396605000000
1!
1%
#396610000000
0!
0%
#396615000000
1!
1%
#396620000000
0!
0%
#396625000000
1!
1%
#396630000000
0!
0%
#396635000000
1!
1%
#396640000000
0!
0%
#396645000000
1!
1%
#396650000000
0!
0%
#396655000000
1!
1%
#396660000000
0!
0%
#396665000000
1!
1%
#396670000000
0!
0%
#396675000000
1!
1%
#396680000000
0!
0%
#396685000000
1!
1%
#396690000000
0!
0%
#396695000000
1!
1%
#396700000000
0!
0%
#396705000000
1!
1%
#396710000000
0!
0%
#396715000000
1!
1%
#396720000000
0!
0%
#396725000000
1!
1%
#396730000000
0!
0%
#396735000000
1!
1%
#396740000000
0!
0%
#396745000000
1!
1%
#396750000000
0!
0%
#396755000000
1!
1%
#396760000000
0!
0%
#396765000000
1!
1%
#396770000000
0!
0%
#396775000000
1!
1%
#396780000000
0!
0%
#396785000000
1!
1%
#396790000000
0!
0%
#396795000000
1!
1%
#396800000000
0!
0%
#396805000000
1!
1%
#396810000000
0!
0%
#396815000000
1!
1%
#396820000000
0!
0%
#396825000000
1!
1%
#396830000000
0!
0%
#396835000000
1!
1%
#396840000000
0!
0%
#396845000000
1!
1%
#396850000000
0!
0%
#396855000000
1!
1%
#396860000000
0!
0%
#396865000000
1!
1%
#396870000000
0!
0%
#396875000000
1!
1%
#396880000000
0!
0%
#396885000000
1!
1%
#396890000000
0!
0%
#396895000000
1!
1%
#396900000000
0!
0%
#396905000000
1!
1%
#396910000000
0!
0%
#396915000000
1!
1%
#396920000000
0!
0%
#396925000000
1!
1%
#396930000000
0!
0%
#396935000000
1!
1%
#396940000000
0!
0%
#396945000000
1!
1%
#396950000000
0!
0%
#396955000000
1!
1%
#396960000000
0!
0%
#396965000000
1!
1%
#396970000000
0!
0%
#396975000000
1!
1%
#396980000000
0!
0%
#396985000000
1!
1%
#396990000000
0!
0%
#396995000000
1!
1%
#397000000000
0!
0%
#397005000000
1!
1%
#397010000000
0!
0%
#397015000000
1!
1%
#397020000000
0!
0%
#397025000000
1!
1%
#397030000000
0!
0%
#397035000000
1!
1%
#397040000000
0!
0%
#397045000000
1!
1%
#397050000000
0!
0%
#397055000000
1!
1%
#397060000000
0!
0%
#397065000000
1!
1%
#397070000000
0!
0%
#397075000000
1!
1%
#397080000000
0!
0%
#397085000000
1!
1%
#397090000000
0!
0%
#397095000000
1!
1%
#397100000000
0!
0%
#397105000000
1!
1%
#397110000000
0!
0%
#397115000000
1!
1%
#397120000000
0!
0%
#397125000000
1!
1%
#397130000000
0!
0%
#397135000000
1!
1%
#397140000000
0!
0%
#397145000000
1!
1%
#397150000000
0!
0%
#397155000000
1!
1%
#397160000000
0!
0%
#397165000000
1!
1%
#397170000000
0!
0%
#397175000000
1!
1%
#397180000000
0!
0%
#397185000000
1!
1%
#397190000000
0!
0%
#397195000000
1!
1%
#397200000000
0!
0%
#397205000000
1!
1%
#397210000000
0!
0%
#397215000000
1!
1%
#397220000000
0!
0%
#397225000000
1!
1%
#397230000000
0!
0%
#397235000000
1!
1%
#397240000000
0!
0%
#397245000000
1!
1%
#397250000000
0!
0%
#397255000000
1!
1%
#397260000000
0!
0%
#397265000000
1!
1%
#397270000000
0!
0%
#397275000000
1!
1%
#397280000000
0!
0%
#397285000000
1!
1%
#397290000000
0!
0%
#397295000000
1!
1%
#397300000000
0!
0%
#397305000000
1!
1%
#397310000000
0!
0%
#397315000000
1!
1%
#397320000000
0!
0%
#397325000000
1!
1%
#397330000000
0!
0%
#397335000000
1!
1%
#397340000000
0!
0%
#397345000000
1!
1%
#397350000000
0!
0%
#397355000000
1!
1%
#397360000000
0!
0%
#397365000000
1!
1%
#397370000000
0!
0%
#397375000000
1!
1%
#397380000000
0!
0%
#397385000000
1!
1%
#397390000000
0!
0%
#397395000000
1!
1%
#397400000000
0!
0%
#397405000000
1!
1%
#397410000000
0!
0%
#397415000000
1!
1%
#397420000000
0!
0%
#397425000000
1!
1%
#397430000000
0!
0%
#397435000000
1!
1%
#397440000000
0!
0%
#397445000000
1!
1%
#397450000000
0!
0%
#397455000000
1!
1%
#397460000000
0!
0%
#397465000000
1!
1%
#397470000000
0!
0%
#397475000000
1!
1%
#397480000000
0!
0%
#397485000000
1!
1%
#397490000000
0!
0%
#397495000000
1!
1%
#397500000000
0!
0%
#397505000000
1!
1%
#397510000000
0!
0%
#397515000000
1!
1%
#397520000000
0!
0%
#397525000000
1!
1%
#397530000000
0!
0%
#397535000000
1!
1%
#397540000000
0!
0%
#397545000000
1!
1%
#397550000000
0!
0%
#397555000000
1!
1%
#397560000000
0!
0%
#397565000000
1!
1%
#397570000000
0!
0%
#397575000000
1!
1%
#397580000000
0!
0%
#397585000000
1!
1%
#397590000000
0!
0%
#397595000000
1!
1%
#397600000000
0!
0%
#397605000000
1!
1%
#397610000000
0!
0%
#397615000000
1!
1%
#397620000000
0!
0%
#397625000000
1!
1%
#397630000000
0!
0%
#397635000000
1!
1%
#397640000000
0!
0%
#397645000000
1!
1%
#397650000000
0!
0%
#397655000000
1!
1%
#397660000000
0!
0%
#397665000000
1!
1%
#397670000000
0!
0%
#397675000000
1!
1%
#397680000000
0!
0%
#397685000000
1!
1%
#397690000000
0!
0%
#397695000000
1!
1%
#397700000000
0!
0%
#397705000000
1!
1%
#397710000000
0!
0%
#397715000000
1!
1%
#397720000000
0!
0%
#397725000000
1!
1%
#397730000000
0!
0%
#397735000000
1!
1%
#397740000000
0!
0%
#397745000000
1!
1%
#397750000000
0!
0%
#397755000000
1!
1%
#397760000000
0!
0%
#397765000000
1!
1%
#397770000000
0!
0%
#397775000000
1!
1%
#397780000000
0!
0%
#397785000000
1!
1%
#397790000000
0!
0%
#397795000000
1!
1%
#397800000000
0!
0%
#397805000000
1!
1%
#397810000000
0!
0%
#397815000000
1!
1%
#397820000000
0!
0%
#397825000000
1!
1%
#397830000000
0!
0%
#397835000000
1!
1%
#397840000000
0!
0%
#397845000000
1!
1%
#397850000000
0!
0%
#397855000000
1!
1%
#397860000000
0!
0%
#397865000000
1!
1%
#397870000000
0!
0%
#397875000000
1!
1%
#397880000000
0!
0%
#397885000000
1!
1%
#397890000000
0!
0%
#397895000000
1!
1%
#397900000000
0!
0%
#397905000000
1!
1%
#397910000000
0!
0%
#397915000000
1!
1%
#397920000000
0!
0%
#397925000000
1!
1%
#397930000000
0!
0%
#397935000000
1!
1%
#397940000000
0!
0%
#397945000000
1!
1%
#397950000000
0!
0%
#397955000000
1!
1%
#397960000000
0!
0%
#397965000000
1!
1%
#397970000000
0!
0%
#397975000000
1!
1%
#397980000000
0!
0%
#397985000000
1!
1%
#397990000000
0!
0%
#397995000000
1!
1%
#398000000000
0!
0%
#398005000000
1!
1%
#398010000000
0!
0%
#398015000000
1!
1%
#398020000000
0!
0%
#398025000000
1!
1%
#398030000000
0!
0%
#398035000000
1!
1%
#398040000000
0!
0%
#398045000000
1!
1%
#398050000000
0!
0%
#398055000000
1!
1%
#398060000000
0!
0%
#398065000000
1!
1%
#398070000000
0!
0%
#398075000000
1!
1%
#398080000000
0!
0%
#398085000000
1!
1%
#398090000000
0!
0%
#398095000000
1!
1%
#398100000000
0!
0%
#398105000000
1!
1%
#398110000000
0!
0%
#398115000000
1!
1%
#398120000000
0!
0%
#398125000000
1!
1%
#398130000000
0!
0%
#398135000000
1!
1%
#398140000000
0!
0%
#398145000000
1!
1%
#398150000000
0!
0%
#398155000000
1!
1%
#398160000000
0!
0%
#398165000000
1!
1%
#398170000000
0!
0%
#398175000000
1!
1%
#398180000000
0!
0%
#398185000000
1!
1%
#398190000000
0!
0%
#398195000000
1!
1%
#398200000000
0!
0%
#398205000000
1!
1%
#398210000000
0!
0%
#398215000000
1!
1%
#398220000000
0!
0%
#398225000000
1!
1%
#398230000000
0!
0%
#398235000000
1!
1%
#398240000000
0!
0%
#398245000000
1!
1%
#398250000000
0!
0%
#398255000000
1!
1%
#398260000000
0!
0%
#398265000000
1!
1%
#398270000000
0!
0%
#398275000000
1!
1%
#398280000000
0!
0%
#398285000000
1!
1%
#398290000000
0!
0%
#398295000000
1!
1%
#398300000000
0!
0%
#398305000000
1!
1%
#398310000000
0!
0%
#398315000000
1!
1%
#398320000000
0!
0%
#398325000000
1!
1%
#398330000000
0!
0%
#398335000000
1!
1%
#398340000000
0!
0%
#398345000000
1!
1%
#398350000000
0!
0%
#398355000000
1!
1%
#398360000000
0!
0%
#398365000000
1!
1%
#398370000000
0!
0%
#398375000000
1!
1%
#398380000000
0!
0%
#398385000000
1!
1%
#398390000000
0!
0%
#398395000000
1!
1%
#398400000000
0!
0%
#398405000000
1!
1%
#398410000000
0!
0%
#398415000000
1!
1%
#398420000000
0!
0%
#398425000000
1!
1%
#398430000000
0!
0%
#398435000000
1!
1%
#398440000000
0!
0%
#398445000000
1!
1%
#398450000000
0!
0%
#398455000000
1!
1%
#398460000000
0!
0%
#398465000000
1!
1%
#398470000000
0!
0%
#398475000000
1!
1%
#398480000000
0!
0%
#398485000000
1!
1%
#398490000000
0!
0%
#398495000000
1!
1%
#398500000000
0!
0%
#398505000000
1!
1%
#398510000000
0!
0%
#398515000000
1!
1%
#398520000000
0!
0%
#398525000000
1!
1%
#398530000000
0!
0%
#398535000000
1!
1%
#398540000000
0!
0%
#398545000000
1!
1%
#398550000000
0!
0%
#398555000000
1!
1%
#398560000000
0!
0%
#398565000000
1!
1%
#398570000000
0!
0%
#398575000000
1!
1%
#398580000000
0!
0%
#398585000000
1!
1%
#398590000000
0!
0%
#398595000000
1!
1%
#398600000000
0!
0%
#398605000000
1!
1%
#398610000000
0!
0%
#398615000000
1!
1%
#398620000000
0!
0%
#398625000000
1!
1%
#398630000000
0!
0%
#398635000000
1!
1%
#398640000000
0!
0%
#398645000000
1!
1%
#398650000000
0!
0%
#398655000000
1!
1%
#398660000000
0!
0%
#398665000000
1!
1%
#398670000000
0!
0%
#398675000000
1!
1%
#398680000000
0!
0%
#398685000000
1!
1%
#398690000000
0!
0%
#398695000000
1!
1%
#398700000000
0!
0%
#398705000000
1!
1%
#398710000000
0!
0%
#398715000000
1!
1%
#398720000000
0!
0%
#398725000000
1!
1%
#398730000000
0!
0%
#398735000000
1!
1%
#398740000000
0!
0%
#398745000000
1!
1%
#398750000000
0!
0%
#398755000000
1!
1%
#398760000000
0!
0%
#398765000000
1!
1%
#398770000000
0!
0%
#398775000000
1!
1%
#398780000000
0!
0%
#398785000000
1!
1%
#398790000000
0!
0%
#398795000000
1!
1%
#398800000000
0!
0%
#398805000000
1!
1%
#398810000000
0!
0%
#398815000000
1!
1%
#398820000000
0!
0%
#398825000000
1!
1%
#398830000000
0!
0%
#398835000000
1!
1%
#398840000000
0!
0%
#398845000000
1!
1%
#398850000000
0!
0%
#398855000000
1!
1%
#398860000000
0!
0%
#398865000000
1!
1%
#398870000000
0!
0%
#398875000000
1!
1%
#398880000000
0!
0%
#398885000000
1!
1%
#398890000000
0!
0%
#398895000000
1!
1%
#398900000000
0!
0%
#398905000000
1!
1%
#398910000000
0!
0%
#398915000000
1!
1%
#398920000000
0!
0%
#398925000000
1!
1%
#398930000000
0!
0%
#398935000000
1!
1%
#398940000000
0!
0%
#398945000000
1!
1%
#398950000000
0!
0%
#398955000000
1!
1%
#398960000000
0!
0%
#398965000000
1!
1%
#398970000000
0!
0%
#398975000000
1!
1%
#398980000000
0!
0%
#398985000000
1!
1%
#398990000000
0!
0%
#398995000000
1!
1%
#399000000000
0!
0%
#399005000000
1!
1%
#399010000000
0!
0%
#399015000000
1!
1%
#399020000000
0!
0%
#399025000000
1!
1%
#399030000000
0!
0%
#399035000000
1!
1%
#399040000000
0!
0%
#399045000000
1!
1%
#399050000000
0!
0%
#399055000000
1!
1%
#399060000000
0!
0%
#399065000000
1!
1%
#399070000000
0!
0%
#399075000000
1!
1%
#399080000000
0!
0%
#399085000000
1!
1%
#399090000000
0!
0%
#399095000000
1!
1%
#399100000000
0!
0%
#399105000000
1!
1%
#399110000000
0!
0%
#399115000000
1!
1%
#399120000000
0!
0%
#399125000000
1!
1%
#399130000000
0!
0%
#399135000000
1!
1%
#399140000000
0!
0%
#399145000000
1!
1%
#399150000000
0!
0%
#399155000000
1!
1%
#399160000000
0!
0%
#399165000000
1!
1%
#399170000000
0!
0%
#399175000000
1!
1%
#399180000000
0!
0%
#399185000000
1!
1%
#399190000000
0!
0%
#399195000000
1!
1%
#399200000000
0!
0%
#399205000000
1!
1%
#399210000000
0!
0%
#399215000000
1!
1%
#399220000000
0!
0%
#399225000000
1!
1%
#399230000000
0!
0%
#399235000000
1!
1%
#399240000000
0!
0%
#399245000000
1!
1%
#399250000000
0!
0%
#399255000000
1!
1%
#399260000000
0!
0%
#399265000000
1!
1%
#399270000000
0!
0%
#399275000000
1!
1%
#399280000000
0!
0%
#399285000000
1!
1%
#399290000000
0!
0%
#399295000000
1!
1%
#399300000000
0!
0%
#399305000000
1!
1%
#399310000000
0!
0%
#399315000000
1!
1%
#399320000000
0!
0%
#399325000000
1!
1%
#399330000000
0!
0%
#399335000000
1!
1%
#399340000000
0!
0%
#399345000000
1!
1%
#399350000000
0!
0%
#399355000000
1!
1%
#399360000000
0!
0%
#399365000000
1!
1%
#399370000000
0!
0%
#399375000000
1!
1%
#399380000000
0!
0%
#399385000000
1!
1%
#399390000000
0!
0%
#399395000000
1!
1%
#399400000000
0!
0%
#399405000000
1!
1%
#399410000000
0!
0%
#399415000000
1!
1%
#399420000000
0!
0%
#399425000000
1!
1%
#399430000000
0!
0%
#399435000000
1!
1%
#399440000000
0!
0%
#399445000000
1!
1%
#399450000000
0!
0%
#399455000000
1!
1%
#399460000000
0!
0%
#399465000000
1!
1%
#399470000000
0!
0%
#399475000000
1!
1%
#399480000000
0!
0%
#399485000000
1!
1%
#399490000000
0!
0%
#399495000000
1!
1%
#399500000000
0!
0%
#399505000000
1!
1%
#399510000000
0!
0%
#399515000000
1!
1%
#399520000000
0!
0%
#399525000000
1!
1%
#399530000000
0!
0%
#399535000000
1!
1%
#399540000000
0!
0%
#399545000000
1!
1%
#399550000000
0!
0%
#399555000000
1!
1%
#399560000000
0!
0%
#399565000000
1!
1%
#399570000000
0!
0%
#399575000000
1!
1%
#399580000000
0!
0%
#399585000000
1!
1%
#399590000000
0!
0%
#399595000000
1!
1%
#399600000000
0!
0%
#399605000000
1!
1%
#399610000000
0!
0%
#399615000000
1!
1%
#399620000000
0!
0%
#399625000000
1!
1%
#399630000000
0!
0%
#399635000000
1!
1%
#399640000000
0!
0%
#399645000000
1!
1%
#399650000000
0!
0%
#399655000000
1!
1%
#399660000000
0!
0%
#399665000000
1!
1%
#399670000000
0!
0%
#399675000000
1!
1%
#399680000000
0!
0%
#399685000000
1!
1%
#399690000000
0!
0%
#399695000000
1!
1%
#399700000000
0!
0%
#399705000000
1!
1%
#399710000000
0!
0%
#399715000000
1!
1%
#399720000000
0!
0%
#399725000000
1!
1%
#399730000000
0!
0%
#399735000000
1!
1%
#399740000000
0!
0%
#399745000000
1!
1%
#399750000000
0!
0%
#399755000000
1!
1%
#399760000000
0!
0%
#399765000000
1!
1%
#399770000000
0!
0%
#399775000000
1!
1%
#399780000000
0!
0%
#399785000000
1!
1%
#399790000000
0!
0%
#399795000000
1!
1%
#399800000000
0!
0%
#399805000000
1!
1%
#399810000000
0!
0%
#399815000000
1!
1%
#399820000000
0!
0%
#399825000000
1!
1%
#399830000000
0!
0%
#399835000000
1!
1%
#399840000000
0!
0%
#399845000000
1!
1%
#399850000000
0!
0%
#399855000000
1!
1%
#399860000000
0!
0%
#399865000000
1!
1%
#399870000000
0!
0%
#399875000000
1!
1%
#399880000000
0!
0%
#399885000000
1!
1%
#399890000000
0!
0%
#399895000000
1!
1%
#399900000000
0!
0%
#399905000000
1!
1%
#399910000000
0!
0%
#399915000000
1!
1%
#399920000000
0!
0%
#399925000000
1!
1%
#399930000000
0!
0%
#399935000000
1!
1%
#399940000000
0!
0%
#399945000000
1!
1%
#399950000000
0!
0%
#399955000000
1!
1%
#399960000000
0!
0%
#399965000000
1!
1%
#399970000000
0!
0%
#399975000000
1!
1%
#399980000000
0!
0%
#399985000000
1!
1%
#399990000000
0!
0%
#399995000000
1!
1%
#400000000000
0!
0%
#400005000000
1!
1%
#400010000000
0!
0%
#400015000000
1!
1%
#400020000000
0!
0%
#400025000000
1!
1%
#400030000000
0!
0%
#400035000000
1!
1%
#400040000000
0!
0%
#400045000000
1!
1%
#400050000000
0!
0%
#400055000000
1!
1%
#400060000000
0!
0%
#400065000000
1!
1%
#400070000000
0!
0%
#400075000000
1!
1%
#400080000000
0!
0%
#400085000000
1!
1%
#400090000000
0!
0%
#400095000000
1!
1%
#400100000000
0!
0%
#400105000000
1!
1%
#400110000000
0!
0%
#400115000000
1!
1%
#400120000000
0!
0%
#400125000000
1!
1%
#400130000000
0!
0%
#400135000000
1!
1%
#400140000000
0!
0%
#400145000000
1!
1%
#400150000000
0!
0%
#400155000000
1!
1%
#400160000000
0!
0%
#400165000000
1!
1%
#400170000000
0!
0%
#400175000000
1!
1%
#400180000000
0!
0%
#400185000000
1!
1%
#400190000000
0!
0%
#400195000000
1!
1%
#400200000000
0!
0%
#400205000000
1!
1%
#400210000000
0!
0%
#400215000000
1!
1%
#400220000000
0!
0%
#400225000000
1!
1%
#400230000000
0!
0%
#400235000000
1!
1%
#400240000000
0!
0%
#400245000000
1!
1%
#400250000000
0!
0%
#400255000000
1!
1%
#400260000000
0!
0%
#400265000000
1!
1%
#400270000000
0!
0%
#400275000000
1!
1%
#400280000000
0!
0%
#400285000000
1!
1%
#400290000000
0!
0%
#400295000000
1!
1%
#400300000000
0!
0%
#400305000000
1!
1%
#400310000000
0!
0%
#400315000000
1!
1%
#400320000000
0!
0%
#400325000000
1!
1%
#400330000000
0!
0%
#400335000000
1!
1%
#400340000000
0!
0%
#400345000000
1!
1%
#400350000000
0!
0%
#400355000000
1!
1%
#400360000000
0!
0%
#400365000000
1!
1%
#400370000000
0!
0%
#400375000000
1!
1%
#400380000000
0!
0%
#400385000000
1!
1%
#400390000000
0!
0%
#400395000000
1!
1%
#400400000000
0!
0%
#400405000000
1!
1%
#400410000000
0!
0%
#400415000000
1!
1%
#400420000000
0!
0%
#400425000000
1!
1%
#400430000000
0!
0%
#400435000000
1!
1%
#400440000000
0!
0%
#400445000000
1!
1%
#400450000000
0!
0%
#400455000000
1!
1%
#400460000000
0!
0%
#400465000000
1!
1%
#400470000000
0!
0%
#400475000000
1!
1%
#400480000000
0!
0%
#400485000000
1!
1%
#400490000000
0!
0%
#400495000000
1!
1%
#400500000000
0!
0%
#400505000000
1!
1%
#400510000000
0!
0%
#400515000000
1!
1%
#400520000000
0!
0%
#400525000000
1!
1%
#400530000000
0!
0%
#400535000000
1!
1%
#400540000000
0!
0%
#400545000000
1!
1%
#400550000000
0!
0%
#400555000000
1!
1%
#400560000000
0!
0%
#400565000000
1!
1%
#400570000000
0!
0%
#400575000000
1!
1%
#400580000000
0!
0%
#400585000000
1!
1%
#400590000000
0!
0%
#400595000000
1!
1%
#400600000000
0!
0%
#400605000000
1!
1%
#400610000000
0!
0%
#400615000000
1!
1%
#400620000000
0!
0%
#400625000000
1!
1%
#400630000000
0!
0%
#400635000000
1!
1%
#400640000000
0!
0%
#400645000000
1!
1%
#400650000000
0!
0%
#400655000000
1!
1%
#400660000000
0!
0%
#400665000000
1!
1%
#400670000000
0!
0%
#400675000000
1!
1%
#400680000000
0!
0%
#400685000000
1!
1%
#400690000000
0!
0%
#400695000000
1!
1%
#400700000000
0!
0%
#400705000000
1!
1%
#400710000000
0!
0%
#400715000000
1!
1%
#400720000000
0!
0%
#400725000000
1!
1%
#400730000000
0!
0%
#400735000000
1!
1%
#400740000000
0!
0%
#400745000000
1!
1%
#400750000000
0!
0%
#400755000000
1!
1%
#400760000000
0!
0%
#400765000000
1!
1%
#400770000000
0!
0%
#400775000000
1!
1%
#400780000000
0!
0%
#400785000000
1!
1%
#400790000000
0!
0%
#400795000000
1!
1%
#400800000000
0!
0%
#400805000000
1!
1%
#400810000000
0!
0%
#400815000000
1!
1%
#400820000000
0!
0%
#400825000000
1!
1%
#400830000000
0!
0%
#400835000000
1!
1%
#400840000000
0!
0%
#400845000000
1!
1%
#400850000000
0!
0%
#400855000000
1!
1%
#400860000000
0!
0%
#400865000000
1!
1%
#400870000000
0!
0%
#400875000000
1!
1%
#400880000000
0!
0%
#400885000000
1!
1%
#400890000000
0!
0%
#400895000000
1!
1%
#400900000000
0!
0%
#400905000000
1!
1%
#400910000000
0!
0%
#400915000000
1!
1%
#400920000000
0!
0%
#400925000000
1!
1%
#400930000000
0!
0%
#400935000000
1!
1%
#400940000000
0!
0%
#400945000000
1!
1%
#400950000000
0!
0%
#400955000000
1!
1%
#400960000000
0!
0%
#400965000000
1!
1%
#400970000000
0!
0%
#400975000000
1!
1%
#400980000000
0!
0%
#400985000000
1!
1%
#400990000000
0!
0%
#400995000000
1!
1%
#401000000000
0!
0%
#401005000000
1!
1%
#401010000000
0!
0%
#401015000000
1!
1%
#401020000000
0!
0%
#401025000000
1!
1%
#401030000000
0!
0%
#401035000000
1!
1%
#401040000000
0!
0%
#401045000000
1!
1%
#401050000000
0!
0%
#401055000000
1!
1%
#401060000000
0!
0%
#401065000000
1!
1%
#401070000000
0!
0%
#401075000000
1!
1%
#401080000000
0!
0%
#401085000000
1!
1%
#401090000000
0!
0%
#401095000000
1!
1%
#401100000000
0!
0%
#401105000000
1!
1%
#401110000000
0!
0%
#401115000000
1!
1%
#401120000000
0!
0%
#401125000000
1!
1%
#401130000000
0!
0%
#401135000000
1!
1%
#401140000000
0!
0%
#401145000000
1!
1%
#401150000000
0!
0%
#401155000000
1!
1%
#401160000000
0!
0%
#401165000000
1!
1%
#401170000000
0!
0%
#401175000000
1!
1%
#401180000000
0!
0%
#401185000000
1!
1%
#401190000000
0!
0%
#401195000000
1!
1%
#401200000000
0!
0%
#401205000000
1!
1%
#401210000000
0!
0%
#401215000000
1!
1%
#401220000000
0!
0%
#401225000000
1!
1%
#401230000000
0!
0%
#401235000000
1!
1%
#401240000000
0!
0%
#401245000000
1!
1%
#401250000000
0!
0%
#401255000000
1!
1%
#401260000000
0!
0%
#401265000000
1!
1%
#401270000000
0!
0%
#401275000000
1!
1%
#401280000000
0!
0%
#401285000000
1!
1%
#401290000000
0!
0%
#401295000000
1!
1%
#401300000000
0!
0%
#401305000000
1!
1%
#401310000000
0!
0%
#401315000000
1!
1%
#401320000000
0!
0%
#401325000000
1!
1%
#401330000000
0!
0%
#401335000000
1!
1%
#401340000000
0!
0%
#401345000000
1!
1%
#401350000000
0!
0%
#401355000000
1!
1%
#401360000000
0!
0%
#401365000000
1!
1%
#401370000000
0!
0%
#401375000000
1!
1%
#401380000000
0!
0%
#401385000000
1!
1%
#401390000000
0!
0%
#401395000000
1!
1%
#401400000000
0!
0%
#401405000000
1!
1%
#401410000000
0!
0%
#401415000000
1!
1%
#401420000000
0!
0%
#401425000000
1!
1%
#401430000000
0!
0%
#401435000000
1!
1%
#401440000000
0!
0%
#401445000000
1!
1%
#401450000000
0!
0%
#401455000000
1!
1%
#401460000000
0!
0%
#401465000000
1!
1%
#401470000000
0!
0%
#401475000000
1!
1%
#401480000000
0!
0%
#401485000000
1!
1%
#401490000000
0!
0%
#401495000000
1!
1%
#401500000000
0!
0%
#401505000000
1!
1%
#401510000000
0!
0%
#401515000000
1!
1%
#401520000000
0!
0%
#401525000000
1!
1%
#401530000000
0!
0%
#401535000000
1!
1%
#401540000000
0!
0%
#401545000000
1!
1%
#401550000000
0!
0%
#401555000000
1!
1%
#401560000000
0!
0%
#401565000000
1!
1%
#401570000000
0!
0%
#401575000000
1!
1%
#401580000000
0!
0%
#401585000000
1!
1%
#401590000000
0!
0%
#401595000000
1!
1%
#401600000000
0!
0%
#401605000000
1!
1%
#401610000000
0!
0%
#401615000000
1!
1%
#401620000000
0!
0%
#401625000000
1!
1%
#401630000000
0!
0%
#401635000000
1!
1%
#401640000000
0!
0%
#401645000000
1!
1%
#401650000000
0!
0%
#401655000000
1!
1%
#401660000000
0!
0%
#401665000000
1!
1%
#401670000000
0!
0%
#401675000000
1!
1%
#401680000000
0!
0%
#401685000000
1!
1%
#401690000000
0!
0%
#401695000000
1!
1%
#401700000000
0!
0%
#401705000000
1!
1%
#401710000000
0!
0%
#401715000000
1!
1%
#401720000000
0!
0%
#401725000000
1!
1%
#401730000000
0!
0%
#401735000000
1!
1%
#401740000000
0!
0%
#401745000000
1!
1%
#401750000000
0!
0%
#401755000000
1!
1%
#401760000000
0!
0%
#401765000000
1!
1%
#401770000000
0!
0%
#401775000000
1!
1%
#401780000000
0!
0%
#401785000000
1!
1%
#401790000000
0!
0%
#401795000000
1!
1%
#401800000000
0!
0%
#401805000000
1!
1%
#401810000000
0!
0%
#401815000000
1!
1%
#401820000000
0!
0%
#401825000000
1!
1%
#401830000000
0!
0%
#401835000000
1!
1%
#401840000000
0!
0%
#401845000000
1!
1%
#401850000000
0!
0%
#401855000000
1!
1%
#401860000000
0!
0%
#401865000000
1!
1%
#401870000000
0!
0%
#401875000000
1!
1%
#401880000000
0!
0%
#401885000000
1!
1%
#401890000000
0!
0%
#401895000000
1!
1%
#401900000000
0!
0%
#401905000000
1!
1%
#401910000000
0!
0%
#401915000000
1!
1%
#401920000000
0!
0%
#401925000000
1!
1%
#401930000000
0!
0%
#401935000000
1!
1%
#401940000000
0!
0%
#401945000000
1!
1%
#401950000000
0!
0%
#401955000000
1!
1%
#401960000000
0!
0%
#401965000000
1!
1%
#401970000000
0!
0%
#401975000000
1!
1%
#401980000000
0!
0%
#401985000000
1!
1%
#401990000000
0!
0%
#401995000000
1!
1%
#402000000000
0!
0%
#402005000000
1!
1%
#402010000000
0!
0%
#402015000000
1!
1%
#402020000000
0!
0%
#402025000000
1!
1%
#402030000000
0!
0%
#402035000000
1!
1%
#402040000000
0!
0%
#402045000000
1!
1%
#402050000000
0!
0%
#402055000000
1!
1%
#402060000000
0!
0%
#402065000000
1!
1%
#402070000000
0!
0%
#402075000000
1!
1%
#402080000000
0!
0%
#402085000000
1!
1%
#402090000000
0!
0%
#402095000000
1!
1%
#402100000000
0!
0%
#402105000000
1!
1%
#402110000000
0!
0%
#402115000000
1!
1%
#402120000000
0!
0%
#402125000000
1!
1%
#402130000000
0!
0%
#402135000000
1!
1%
#402140000000
0!
0%
#402145000000
1!
1%
#402150000000
0!
0%
#402155000000
1!
1%
#402160000000
0!
0%
#402165000000
1!
1%
#402170000000
0!
0%
#402175000000
1!
1%
#402180000000
0!
0%
#402185000000
1!
1%
#402190000000
0!
0%
#402195000000
1!
1%
#402200000000
0!
0%
#402205000000
1!
1%
#402210000000
0!
0%
#402215000000
1!
1%
#402220000000
0!
0%
#402225000000
1!
1%
#402230000000
0!
0%
#402235000000
1!
1%
#402240000000
0!
0%
#402245000000
1!
1%
#402250000000
0!
0%
#402255000000
1!
1%
#402260000000
0!
0%
#402265000000
1!
1%
#402270000000
0!
0%
#402275000000
1!
1%
#402280000000
0!
0%
#402285000000
1!
1%
#402290000000
0!
0%
#402295000000
1!
1%
#402300000000
0!
0%
#402305000000
1!
1%
#402310000000
0!
0%
#402315000000
1!
1%
#402320000000
0!
0%
#402325000000
1!
1%
#402330000000
0!
0%
#402335000000
1!
1%
#402340000000
0!
0%
#402345000000
1!
1%
#402350000000
0!
0%
#402355000000
1!
1%
#402360000000
0!
0%
#402365000000
1!
1%
#402370000000
0!
0%
#402375000000
1!
1%
#402380000000
0!
0%
#402385000000
1!
1%
#402390000000
0!
0%
#402395000000
1!
1%
#402400000000
0!
0%
#402405000000
1!
1%
#402410000000
0!
0%
#402415000000
1!
1%
#402420000000
0!
0%
#402425000000
1!
1%
#402430000000
0!
0%
#402435000000
1!
1%
#402440000000
0!
0%
#402445000000
1!
1%
#402450000000
0!
0%
#402455000000
1!
1%
#402460000000
0!
0%
#402465000000
1!
1%
#402470000000
0!
0%
#402475000000
1!
1%
#402480000000
0!
0%
#402485000000
1!
1%
#402490000000
0!
0%
#402495000000
1!
1%
#402500000000
0!
0%
#402505000000
1!
1%
#402510000000
0!
0%
#402515000000
1!
1%
#402520000000
0!
0%
#402525000000
1!
1%
#402530000000
0!
0%
#402535000000
1!
1%
#402540000000
0!
0%
#402545000000
1!
1%
#402550000000
0!
0%
#402555000000
1!
1%
#402560000000
0!
0%
#402565000000
1!
1%
#402570000000
0!
0%
#402575000000
1!
1%
#402580000000
0!
0%
#402585000000
1!
1%
#402590000000
0!
0%
#402595000000
1!
1%
#402600000000
0!
0%
#402605000000
1!
1%
#402610000000
0!
0%
#402615000000
1!
1%
#402620000000
0!
0%
#402625000000
1!
1%
#402630000000
0!
0%
#402635000000
1!
1%
#402640000000
0!
0%
#402645000000
1!
1%
#402650000000
0!
0%
#402655000000
1!
1%
#402660000000
0!
0%
#402665000000
1!
1%
#402670000000
0!
0%
#402675000000
1!
1%
#402680000000
0!
0%
#402685000000
1!
1%
#402690000000
0!
0%
#402695000000
1!
1%
#402700000000
0!
0%
#402705000000
1!
1%
#402710000000
0!
0%
#402715000000
1!
1%
#402720000000
0!
0%
#402725000000
1!
1%
#402730000000
0!
0%
#402735000000
1!
1%
#402740000000
0!
0%
#402745000000
1!
1%
#402750000000
0!
0%
#402755000000
1!
1%
#402760000000
0!
0%
#402765000000
1!
1%
#402770000000
0!
0%
#402775000000
1!
1%
#402780000000
0!
0%
#402785000000
1!
1%
#402790000000
0!
0%
#402795000000
1!
1%
#402800000000
0!
0%
#402805000000
1!
1%
#402810000000
0!
0%
#402815000000
1!
1%
#402820000000
0!
0%
#402825000000
1!
1%
#402830000000
0!
0%
#402835000000
1!
1%
#402840000000
0!
0%
#402845000000
1!
1%
#402850000000
0!
0%
#402855000000
1!
1%
#402860000000
0!
0%
#402865000000
1!
1%
#402870000000
0!
0%
#402875000000
1!
1%
#402880000000
0!
0%
#402885000000
1!
1%
#402890000000
0!
0%
#402895000000
1!
1%
#402900000000
0!
0%
#402905000000
1!
1%
#402910000000
0!
0%
#402915000000
1!
1%
#402920000000
0!
0%
#402925000000
1!
1%
#402930000000
0!
0%
#402935000000
1!
1%
#402940000000
0!
0%
#402945000000
1!
1%
#402950000000
0!
0%
#402955000000
1!
1%
#402960000000
0!
0%
#402965000000
1!
1%
#402970000000
0!
0%
#402975000000
1!
1%
#402980000000
0!
0%
#402985000000
1!
1%
#402990000000
0!
0%
#402995000000
1!
1%
#403000000000
0!
0%
#403005000000
1!
1%
#403010000000
0!
0%
#403015000000
1!
1%
#403020000000
0!
0%
#403025000000
1!
1%
#403030000000
0!
0%
#403035000000
1!
1%
#403040000000
0!
0%
#403045000000
1!
1%
#403050000000
0!
0%
#403055000000
1!
1%
#403060000000
0!
0%
#403065000000
1!
1%
#403070000000
0!
0%
#403075000000
1!
1%
#403080000000
0!
0%
#403085000000
1!
1%
#403090000000
0!
0%
#403095000000
1!
1%
#403100000000
0!
0%
#403105000000
1!
1%
#403110000000
0!
0%
#403115000000
1!
1%
#403120000000
0!
0%
#403125000000
1!
1%
#403130000000
0!
0%
#403135000000
1!
1%
#403140000000
0!
0%
#403145000000
1!
1%
#403150000000
0!
0%
#403155000000
1!
1%
#403160000000
0!
0%
#403165000000
1!
1%
#403170000000
0!
0%
#403175000000
1!
1%
#403180000000
0!
0%
#403185000000
1!
1%
#403190000000
0!
0%
#403195000000
1!
1%
#403200000000
0!
0%
#403205000000
1!
1%
#403210000000
0!
0%
#403215000000
1!
1%
#403220000000
0!
0%
#403225000000
1!
1%
#403230000000
0!
0%
#403235000000
1!
1%
#403240000000
0!
0%
#403245000000
1!
1%
#403250000000
0!
0%
#403255000000
1!
1%
#403260000000
0!
0%
#403265000000
1!
1%
#403270000000
0!
0%
#403275000000
1!
1%
#403280000000
0!
0%
#403285000000
1!
1%
#403290000000
0!
0%
#403295000000
1!
1%
#403300000000
0!
0%
#403305000000
1!
1%
#403310000000
0!
0%
#403315000000
1!
1%
#403320000000
0!
0%
#403325000000
1!
1%
#403330000000
0!
0%
#403335000000
1!
1%
#403340000000
0!
0%
#403345000000
1!
1%
#403350000000
0!
0%
#403355000000
1!
1%
#403360000000
0!
0%
#403365000000
1!
1%
#403370000000
0!
0%
#403375000000
1!
1%
#403380000000
0!
0%
#403385000000
1!
1%
#403390000000
0!
0%
#403395000000
1!
1%
#403400000000
0!
0%
#403405000000
1!
1%
#403410000000
0!
0%
#403415000000
1!
1%
#403420000000
0!
0%
#403425000000
1!
1%
#403430000000
0!
0%
#403435000000
1!
1%
#403440000000
0!
0%
#403445000000
1!
1%
#403450000000
0!
0%
#403455000000
1!
1%
#403460000000
0!
0%
#403465000000
1!
1%
#403470000000
0!
0%
#403475000000
1!
1%
#403480000000
0!
0%
#403485000000
1!
1%
#403490000000
0!
0%
#403495000000
1!
1%
#403500000000
0!
0%
#403505000000
1!
1%
#403510000000
0!
0%
#403515000000
1!
1%
#403520000000
0!
0%
#403525000000
1!
1%
#403530000000
0!
0%
#403535000000
1!
1%
#403540000000
0!
0%
#403545000000
1!
1%
#403550000000
0!
0%
#403555000000
1!
1%
#403560000000
0!
0%
#403565000000
1!
1%
#403570000000
0!
0%
#403575000000
1!
1%
#403580000000
0!
0%
#403585000000
1!
1%
#403590000000
0!
0%
#403595000000
1!
1%
#403600000000
0!
0%
#403605000000
1!
1%
#403610000000
0!
0%
#403615000000
1!
1%
#403620000000
0!
0%
#403625000000
1!
1%
#403630000000
0!
0%
#403635000000
1!
1%
#403640000000
0!
0%
#403645000000
1!
1%
#403650000000
0!
0%
#403655000000
1!
1%
#403660000000
0!
0%
#403665000000
1!
1%
#403670000000
0!
0%
#403675000000
1!
1%
#403680000000
0!
0%
#403685000000
1!
1%
#403690000000
0!
0%
#403695000000
1!
1%
#403700000000
0!
0%
#403705000000
1!
1%
#403710000000
0!
0%
#403715000000
1!
1%
#403720000000
0!
0%
#403725000000
1!
1%
#403730000000
0!
0%
#403735000000
1!
1%
#403740000000
0!
0%
#403745000000
1!
1%
#403750000000
0!
0%
#403755000000
1!
1%
#403760000000
0!
0%
#403765000000
1!
1%
#403770000000
0!
0%
#403775000000
1!
1%
#403780000000
0!
0%
#403785000000
1!
1%
#403790000000
0!
0%
#403795000000
1!
1%
#403800000000
0!
0%
#403805000000
1!
1%
#403810000000
0!
0%
#403815000000
1!
1%
#403820000000
0!
0%
#403825000000
1!
1%
#403830000000
0!
0%
#403835000000
1!
1%
#403840000000
0!
0%
#403845000000
1!
1%
#403850000000
0!
0%
#403855000000
1!
1%
#403860000000
0!
0%
#403865000000
1!
1%
#403870000000
0!
0%
#403875000000
1!
1%
#403880000000
0!
0%
#403885000000
1!
1%
#403890000000
0!
0%
#403895000000
1!
1%
#403900000000
0!
0%
#403905000000
1!
1%
#403910000000
0!
0%
#403915000000
1!
1%
#403920000000
0!
0%
#403925000000
1!
1%
#403930000000
0!
0%
#403935000000
1!
1%
#403940000000
0!
0%
#403945000000
1!
1%
#403950000000
0!
0%
#403955000000
1!
1%
#403960000000
0!
0%
#403965000000
1!
1%
#403970000000
0!
0%
#403975000000
1!
1%
#403980000000
0!
0%
#403985000000
1!
1%
#403990000000
0!
0%
#403995000000
1!
1%
#404000000000
0!
0%
#404005000000
1!
1%
#404010000000
0!
0%
#404015000000
1!
1%
#404020000000
0!
0%
#404025000000
1!
1%
#404030000000
0!
0%
#404035000000
1!
1%
#404040000000
0!
0%
#404045000000
1!
1%
#404050000000
0!
0%
#404055000000
1!
1%
#404060000000
0!
0%
#404065000000
1!
1%
#404070000000
0!
0%
#404075000000
1!
1%
#404080000000
0!
0%
#404085000000
1!
1%
#404090000000
0!
0%
#404095000000
1!
1%
#404100000000
0!
0%
#404105000000
1!
1%
#404110000000
0!
0%
#404115000000
1!
1%
#404120000000
0!
0%
#404125000000
1!
1%
#404130000000
0!
0%
#404135000000
1!
1%
#404140000000
0!
0%
#404145000000
1!
1%
#404150000000
0!
0%
#404155000000
1!
1%
#404160000000
0!
0%
#404165000000
1!
1%
#404170000000
0!
0%
#404175000000
1!
1%
#404180000000
0!
0%
#404185000000
1!
1%
#404190000000
0!
0%
#404195000000
1!
1%
#404200000000
0!
0%
#404205000000
1!
1%
#404210000000
0!
0%
#404215000000
1!
1%
#404220000000
0!
0%
#404225000000
1!
1%
#404230000000
0!
0%
#404235000000
1!
1%
#404240000000
0!
0%
#404245000000
1!
1%
#404250000000
0!
0%
#404255000000
1!
1%
#404260000000
0!
0%
#404265000000
1!
1%
#404270000000
0!
0%
#404275000000
1!
1%
#404280000000
0!
0%
#404285000000
1!
1%
#404290000000
0!
0%
#404295000000
1!
1%
#404300000000
0!
0%
#404305000000
1!
1%
#404310000000
0!
0%
#404315000000
1!
1%
#404320000000
0!
0%
#404325000000
1!
1%
#404330000000
0!
0%
#404335000000
1!
1%
#404340000000
0!
0%
#404345000000
1!
1%
#404350000000
0!
0%
#404355000000
1!
1%
#404360000000
0!
0%
#404365000000
1!
1%
#404370000000
0!
0%
#404375000000
1!
1%
#404380000000
0!
0%
#404385000000
1!
1%
#404390000000
0!
0%
#404395000000
1!
1%
#404400000000
0!
0%
#404405000000
1!
1%
#404410000000
0!
0%
#404415000000
1!
1%
#404420000000
0!
0%
#404425000000
1!
1%
#404430000000
0!
0%
#404435000000
1!
1%
#404440000000
0!
0%
#404445000000
1!
1%
#404450000000
0!
0%
#404455000000
1!
1%
#404460000000
0!
0%
#404465000000
1!
1%
#404470000000
0!
0%
#404475000000
1!
1%
#404480000000
0!
0%
#404485000000
1!
1%
#404490000000
0!
0%
#404495000000
1!
1%
#404500000000
0!
0%
#404505000000
1!
1%
#404510000000
0!
0%
#404515000000
1!
1%
#404520000000
0!
0%
#404525000000
1!
1%
#404530000000
0!
0%
#404535000000
1!
1%
#404540000000
0!
0%
#404545000000
1!
1%
#404550000000
0!
0%
#404555000000
1!
1%
#404560000000
0!
0%
#404565000000
1!
1%
#404570000000
0!
0%
#404575000000
1!
1%
#404580000000
0!
0%
#404585000000
1!
1%
#404590000000
0!
0%
#404595000000
1!
1%
#404600000000
0!
0%
#404605000000
1!
1%
#404610000000
0!
0%
#404615000000
1!
1%
#404620000000
0!
0%
#404625000000
1!
1%
#404630000000
0!
0%
#404635000000
1!
1%
#404640000000
0!
0%
#404645000000
1!
1%
#404650000000
0!
0%
#404655000000
1!
1%
#404660000000
0!
0%
#404665000000
1!
1%
#404670000000
0!
0%
#404675000000
1!
1%
#404680000000
0!
0%
#404685000000
1!
1%
#404690000000
0!
0%
#404695000000
1!
1%
#404700000000
0!
0%
#404705000000
1!
1%
#404710000000
0!
0%
#404715000000
1!
1%
#404720000000
0!
0%
#404725000000
1!
1%
#404730000000
0!
0%
#404735000000
1!
1%
#404740000000
0!
0%
#404745000000
1!
1%
#404750000000
0!
0%
#404755000000
1!
1%
#404760000000
0!
0%
#404765000000
1!
1%
#404770000000
0!
0%
#404775000000
1!
1%
#404780000000
0!
0%
#404785000000
1!
1%
#404790000000
0!
0%
#404795000000
1!
1%
#404800000000
0!
0%
#404805000000
1!
1%
#404810000000
0!
0%
#404815000000
1!
1%
#404820000000
0!
0%
#404825000000
1!
1%
#404830000000
0!
0%
#404835000000
1!
1%
#404840000000
0!
0%
#404845000000
1!
1%
#404850000000
0!
0%
#404855000000
1!
1%
#404860000000
0!
0%
#404865000000
1!
1%
#404870000000
0!
0%
#404875000000
1!
1%
#404880000000
0!
0%
#404885000000
1!
1%
#404890000000
0!
0%
#404895000000
1!
1%
#404900000000
0!
0%
#404905000000
1!
1%
#404910000000
0!
0%
#404915000000
1!
1%
#404920000000
0!
0%
#404925000000
1!
1%
#404930000000
0!
0%
#404935000000
1!
1%
#404940000000
0!
0%
#404945000000
1!
1%
#404950000000
0!
0%
#404955000000
1!
1%
#404960000000
0!
0%
#404965000000
1!
1%
#404970000000
0!
0%
#404975000000
1!
1%
#404980000000
0!
0%
#404985000000
1!
1%
#404990000000
0!
0%
#404995000000
1!
1%
#405000000000
0!
0%
#405005000000
1!
1%
#405010000000
0!
0%
#405015000000
1!
1%
#405020000000
0!
0%
#405025000000
1!
1%
#405030000000
0!
0%
#405035000000
1!
1%
#405040000000
0!
0%
#405045000000
1!
1%
#405050000000
0!
0%
#405055000000
1!
1%
#405060000000
0!
0%
#405065000000
1!
1%
#405070000000
0!
0%
#405075000000
1!
1%
#405080000000
0!
0%
#405085000000
1!
1%
#405090000000
0!
0%
#405095000000
1!
1%
#405100000000
0!
0%
#405105000000
1!
1%
#405110000000
0!
0%
#405115000000
1!
1%
#405120000000
0!
0%
#405125000000
1!
1%
#405130000000
0!
0%
#405135000000
1!
1%
#405140000000
0!
0%
#405145000000
1!
1%
#405150000000
0!
0%
#405155000000
1!
1%
#405160000000
0!
0%
#405165000000
1!
1%
#405170000000
0!
0%
#405175000000
1!
1%
#405180000000
0!
0%
#405185000000
1!
1%
#405190000000
0!
0%
#405195000000
1!
1%
#405200000000
0!
0%
#405205000000
1!
1%
#405210000000
0!
0%
#405215000000
1!
1%
#405220000000
0!
0%
#405225000000
1!
1%
#405230000000
0!
0%
#405235000000
1!
1%
#405240000000
0!
0%
#405245000000
1!
1%
#405250000000
0!
0%
#405255000000
1!
1%
#405260000000
0!
0%
#405265000000
1!
1%
#405270000000
0!
0%
#405275000000
1!
1%
#405280000000
0!
0%
#405285000000
1!
1%
#405290000000
0!
0%
#405295000000
1!
1%
#405300000000
0!
0%
#405305000000
1!
1%
#405310000000
0!
0%
#405315000000
1!
1%
#405320000000
0!
0%
#405325000000
1!
1%
#405330000000
0!
0%
#405335000000
1!
1%
#405340000000
0!
0%
#405345000000
1!
1%
#405350000000
0!
0%
#405355000000
1!
1%
#405360000000
0!
0%
#405365000000
1!
1%
#405370000000
0!
0%
#405375000000
1!
1%
#405380000000
0!
0%
#405385000000
1!
1%
#405390000000
0!
0%
#405395000000
1!
1%
#405400000000
0!
0%
#405405000000
1!
1%
#405410000000
0!
0%
#405415000000
1!
1%
#405420000000
0!
0%
#405425000000
1!
1%
#405430000000
0!
0%
#405435000000
1!
1%
#405440000000
0!
0%
#405445000000
1!
1%
#405450000000
0!
0%
#405455000000
1!
1%
#405460000000
0!
0%
#405465000000
1!
1%
#405470000000
0!
0%
#405475000000
1!
1%
#405480000000
0!
0%
#405485000000
1!
1%
#405490000000
0!
0%
#405495000000
1!
1%
#405500000000
0!
0%
#405505000000
1!
1%
#405510000000
0!
0%
#405515000000
1!
1%
#405520000000
0!
0%
#405525000000
1!
1%
#405530000000
0!
0%
#405535000000
1!
1%
#405540000000
0!
0%
#405545000000
1!
1%
#405550000000
0!
0%
#405555000000
1!
1%
#405560000000
0!
0%
#405565000000
1!
1%
#405570000000
0!
0%
#405575000000
1!
1%
#405580000000
0!
0%
#405585000000
1!
1%
#405590000000
0!
0%
#405595000000
1!
1%
#405600000000
0!
0%
#405605000000
1!
1%
#405610000000
0!
0%
#405615000000
1!
1%
#405620000000
0!
0%
#405625000000
1!
1%
#405630000000
0!
0%
#405635000000
1!
1%
#405640000000
0!
0%
#405645000000
1!
1%
#405650000000
0!
0%
#405655000000
1!
1%
#405660000000
0!
0%
#405665000000
1!
1%
#405670000000
0!
0%
#405675000000
1!
1%
#405680000000
0!
0%
#405685000000
1!
1%
#405690000000
0!
0%
#405695000000
1!
1%
#405700000000
0!
0%
#405705000000
1!
1%
#405710000000
0!
0%
#405715000000
1!
1%
#405720000000
0!
0%
#405725000000
1!
1%
#405730000000
0!
0%
#405735000000
1!
1%
#405740000000
0!
0%
#405745000000
1!
1%
#405750000000
0!
0%
#405755000000
1!
1%
#405760000000
0!
0%
#405765000000
1!
1%
#405770000000
0!
0%
#405775000000
1!
1%
#405780000000
0!
0%
#405785000000
1!
1%
#405790000000
0!
0%
#405795000000
1!
1%
#405800000000
0!
0%
#405805000000
1!
1%
#405810000000
0!
0%
#405815000000
1!
1%
#405820000000
0!
0%
#405825000000
1!
1%
#405830000000
0!
0%
#405835000000
1!
1%
#405840000000
0!
0%
#405845000000
1!
1%
#405850000000
0!
0%
#405855000000
1!
1%
#405860000000
0!
0%
#405865000000
1!
1%
#405870000000
0!
0%
#405875000000
1!
1%
#405880000000
0!
0%
#405885000000
1!
1%
#405890000000
0!
0%
#405895000000
1!
1%
#405900000000
0!
0%
#405905000000
1!
1%
#405910000000
0!
0%
#405915000000
1!
1%
#405920000000
0!
0%
#405925000000
1!
1%
#405930000000
0!
0%
#405935000000
1!
1%
#405940000000
0!
0%
#405945000000
1!
1%
#405950000000
0!
0%
#405955000000
1!
1%
#405960000000
0!
0%
#405965000000
1!
1%
#405970000000
0!
0%
#405975000000
1!
1%
#405980000000
0!
0%
#405985000000
1!
1%
#405990000000
0!
0%
#405995000000
1!
1%
#406000000000
0!
0%
#406005000000
1!
1%
#406010000000
0!
0%
#406015000000
1!
1%
#406020000000
0!
0%
#406025000000
1!
1%
#406030000000
0!
0%
#406035000000
1!
1%
#406040000000
0!
0%
#406045000000
1!
1%
#406050000000
0!
0%
#406055000000
1!
1%
#406060000000
0!
0%
#406065000000
1!
1%
#406070000000
0!
0%
#406075000000
1!
1%
#406080000000
0!
0%
#406085000000
1!
1%
#406090000000
0!
0%
#406095000000
1!
1%
#406100000000
0!
0%
#406105000000
1!
1%
#406110000000
0!
0%
#406115000000
1!
1%
#406120000000
0!
0%
#406125000000
1!
1%
#406130000000
0!
0%
#406135000000
1!
1%
#406140000000
0!
0%
#406145000000
1!
1%
#406150000000
0!
0%
#406155000000
1!
1%
#406160000000
0!
0%
#406165000000
1!
1%
#406170000000
0!
0%
#406175000000
1!
1%
#406180000000
0!
0%
#406185000000
1!
1%
#406190000000
0!
0%
#406195000000
1!
1%
#406200000000
0!
0%
#406205000000
1!
1%
#406210000000
0!
0%
#406215000000
1!
1%
#406220000000
0!
0%
#406225000000
1!
1%
#406230000000
0!
0%
#406235000000
1!
1%
#406240000000
0!
0%
#406245000000
1!
1%
#406250000000
0!
0%
#406255000000
1!
1%
#406260000000
0!
0%
#406265000000
1!
1%
#406270000000
0!
0%
#406275000000
1!
1%
#406280000000
0!
0%
#406285000000
1!
1%
#406290000000
0!
0%
#406295000000
1!
1%
#406300000000
0!
0%
#406305000000
1!
1%
#406310000000
0!
0%
#406315000000
1!
1%
#406320000000
0!
0%
#406325000000
1!
1%
#406330000000
0!
0%
#406335000000
1!
1%
#406340000000
0!
0%
#406345000000
1!
1%
#406350000000
0!
0%
#406355000000
1!
1%
#406360000000
0!
0%
#406365000000
1!
1%
#406370000000
0!
0%
#406375000000
1!
1%
#406380000000
0!
0%
#406385000000
1!
1%
#406390000000
0!
0%
#406395000000
1!
1%
#406400000000
0!
0%
#406405000000
1!
1%
#406410000000
0!
0%
#406415000000
1!
1%
#406420000000
0!
0%
#406425000000
1!
1%
#406430000000
0!
0%
#406435000000
1!
1%
#406440000000
0!
0%
#406445000000
1!
1%
#406450000000
0!
0%
#406455000000
1!
1%
#406460000000
0!
0%
#406465000000
1!
1%
#406470000000
0!
0%
#406475000000
1!
1%
#406480000000
0!
0%
#406485000000
1!
1%
#406490000000
0!
0%
#406495000000
1!
1%
#406500000000
0!
0%
#406505000000
1!
1%
#406510000000
0!
0%
#406515000000
1!
1%
#406520000000
0!
0%
#406525000000
1!
1%
#406530000000
0!
0%
#406535000000
1!
1%
#406540000000
0!
0%
#406545000000
1!
1%
#406550000000
0!
0%
#406555000000
1!
1%
#406560000000
0!
0%
#406565000000
1!
1%
#406570000000
0!
0%
#406575000000
1!
1%
#406580000000
0!
0%
#406585000000
1!
1%
#406590000000
0!
0%
#406595000000
1!
1%
#406600000000
0!
0%
#406605000000
1!
1%
#406610000000
0!
0%
#406615000000
1!
1%
#406620000000
0!
0%
#406625000000
1!
1%
#406630000000
0!
0%
#406635000000
1!
1%
#406640000000
0!
0%
#406645000000
1!
1%
#406650000000
0!
0%
#406655000000
1!
1%
#406660000000
0!
0%
#406665000000
1!
1%
#406670000000
0!
0%
#406675000000
1!
1%
#406680000000
0!
0%
#406685000000
1!
1%
#406690000000
0!
0%
#406695000000
1!
1%
#406700000000
0!
0%
#406705000000
1!
1%
#406710000000
0!
0%
#406715000000
1!
1%
#406720000000
0!
0%
#406725000000
1!
1%
#406730000000
0!
0%
#406735000000
1!
1%
#406740000000
0!
0%
#406745000000
1!
1%
#406750000000
0!
0%
#406755000000
1!
1%
#406760000000
0!
0%
#406765000000
1!
1%
#406770000000
0!
0%
#406775000000
1!
1%
#406780000000
0!
0%
#406785000000
1!
1%
#406790000000
0!
0%
#406795000000
1!
1%
#406800000000
0!
0%
#406805000000
1!
1%
#406810000000
0!
0%
#406815000000
1!
1%
#406820000000
0!
0%
#406825000000
1!
1%
#406830000000
0!
0%
#406835000000
1!
1%
#406840000000
0!
0%
#406845000000
1!
1%
#406850000000
0!
0%
#406855000000
1!
1%
#406860000000
0!
0%
#406865000000
1!
1%
#406870000000
0!
0%
#406875000000
1!
1%
#406880000000
0!
0%
#406885000000
1!
1%
#406890000000
0!
0%
#406895000000
1!
1%
#406900000000
0!
0%
#406905000000
1!
1%
#406910000000
0!
0%
#406915000000
1!
1%
#406920000000
0!
0%
#406925000000
1!
1%
#406930000000
0!
0%
#406935000000
1!
1%
#406940000000
0!
0%
#406945000000
1!
1%
#406950000000
0!
0%
#406955000000
1!
1%
#406960000000
0!
0%
#406965000000
1!
1%
#406970000000
0!
0%
#406975000000
1!
1%
#406980000000
0!
0%
#406985000000
1!
1%
#406990000000
0!
0%
#406995000000
1!
1%
#407000000000
0!
0%
#407005000000
1!
1%
#407010000000
0!
0%
#407015000000
1!
1%
#407020000000
0!
0%
#407025000000
1!
1%
#407030000000
0!
0%
#407035000000
1!
1%
#407040000000
0!
0%
#407045000000
1!
1%
#407050000000
0!
0%
#407055000000
1!
1%
#407060000000
0!
0%
#407065000000
1!
1%
#407070000000
0!
0%
#407075000000
1!
1%
#407080000000
0!
0%
#407085000000
1!
1%
#407090000000
0!
0%
#407095000000
1!
1%
#407100000000
0!
0%
#407105000000
1!
1%
#407110000000
0!
0%
#407115000000
1!
1%
#407120000000
0!
0%
#407125000000
1!
1%
#407130000000
0!
0%
#407135000000
1!
1%
#407140000000
0!
0%
#407145000000
1!
1%
#407150000000
0!
0%
#407155000000
1!
1%
#407160000000
0!
0%
#407165000000
1!
1%
#407170000000
0!
0%
#407175000000
1!
1%
#407180000000
0!
0%
#407185000000
1!
1%
#407190000000
0!
0%
#407195000000
1!
1%
#407200000000
0!
0%
#407205000000
1!
1%
#407210000000
0!
0%
#407215000000
1!
1%
#407220000000
0!
0%
#407225000000
1!
1%
#407230000000
0!
0%
#407235000000
1!
1%
#407240000000
0!
0%
#407245000000
1!
1%
#407250000000
0!
0%
#407255000000
1!
1%
#407260000000
0!
0%
#407265000000
1!
1%
#407270000000
0!
0%
#407275000000
1!
1%
#407280000000
0!
0%
#407285000000
1!
1%
#407290000000
0!
0%
#407295000000
1!
1%
#407300000000
0!
0%
#407305000000
1!
1%
#407310000000
0!
0%
#407315000000
1!
1%
#407320000000
0!
0%
#407325000000
1!
1%
#407330000000
0!
0%
#407335000000
1!
1%
#407340000000
0!
0%
#407345000000
1!
1%
#407350000000
0!
0%
#407355000000
1!
1%
#407360000000
0!
0%
#407365000000
1!
1%
#407370000000
0!
0%
#407375000000
1!
1%
#407380000000
0!
0%
#407385000000
1!
1%
#407390000000
0!
0%
#407395000000
1!
1%
#407400000000
0!
0%
#407405000000
1!
1%
#407410000000
0!
0%
#407415000000
1!
1%
#407420000000
0!
0%
#407425000000
1!
1%
#407430000000
0!
0%
#407435000000
1!
1%
#407440000000
0!
0%
#407445000000
1!
1%
#407450000000
0!
0%
#407455000000
1!
1%
#407460000000
0!
0%
#407465000000
1!
1%
#407470000000
0!
0%
#407475000000
1!
1%
#407480000000
0!
0%
#407485000000
1!
1%
#407490000000
0!
0%
#407495000000
1!
1%
#407500000000
0!
0%
#407505000000
1!
1%
#407510000000
0!
0%
#407515000000
1!
1%
#407520000000
0!
0%
#407525000000
1!
1%
#407530000000
0!
0%
#407535000000
1!
1%
#407540000000
0!
0%
#407545000000
1!
1%
#407550000000
0!
0%
#407555000000
1!
1%
#407560000000
0!
0%
#407565000000
1!
1%
#407570000000
0!
0%
#407575000000
1!
1%
#407580000000
0!
0%
#407585000000
1!
1%
#407590000000
0!
0%
#407595000000
1!
1%
#407600000000
0!
0%
#407605000000
1!
1%
#407610000000
0!
0%
#407615000000
1!
1%
#407620000000
0!
0%
#407625000000
1!
1%
#407630000000
0!
0%
#407635000000
1!
1%
#407640000000
0!
0%
#407645000000
1!
1%
#407650000000
0!
0%
#407655000000
1!
1%
#407660000000
0!
0%
#407665000000
1!
1%
#407670000000
0!
0%
#407675000000
1!
1%
#407680000000
0!
0%
#407685000000
1!
1%
#407690000000
0!
0%
#407695000000
1!
1%
#407700000000
0!
0%
#407705000000
1!
1%
#407710000000
0!
0%
#407715000000
1!
1%
#407720000000
0!
0%
#407725000000
1!
1%
#407730000000
0!
0%
#407735000000
1!
1%
#407740000000
0!
0%
#407745000000
1!
1%
#407750000000
0!
0%
#407755000000
1!
1%
#407760000000
0!
0%
#407765000000
1!
1%
#407770000000
0!
0%
#407775000000
1!
1%
#407780000000
0!
0%
#407785000000
1!
1%
#407790000000
0!
0%
#407795000000
1!
1%
#407800000000
0!
0%
#407805000000
1!
1%
#407810000000
0!
0%
#407815000000
1!
1%
#407820000000
0!
0%
#407825000000
1!
1%
#407830000000
0!
0%
#407835000000
1!
1%
#407840000000
0!
0%
#407845000000
1!
1%
#407850000000
0!
0%
#407855000000
1!
1%
#407860000000
0!
0%
#407865000000
1!
1%
#407870000000
0!
0%
#407875000000
1!
1%
#407880000000
0!
0%
#407885000000
1!
1%
#407890000000
0!
0%
#407895000000
1!
1%
#407900000000
0!
0%
#407905000000
1!
1%
#407910000000
0!
0%
#407915000000
1!
1%
#407920000000
0!
0%
#407925000000
1!
1%
#407930000000
0!
0%
#407935000000
1!
1%
#407940000000
0!
0%
#407945000000
1!
1%
#407950000000
0!
0%
#407955000000
1!
1%
#407960000000
0!
0%
#407965000000
1!
1%
#407970000000
0!
0%
#407975000000
1!
1%
#407980000000
0!
0%
#407985000000
1!
1%
#407990000000
0!
0%
#407995000000
1!
1%
#408000000000
0!
0%
#408005000000
1!
1%
#408010000000
0!
0%
#408015000000
1!
1%
#408020000000
0!
0%
#408025000000
1!
1%
#408030000000
0!
0%
#408035000000
1!
1%
#408040000000
0!
0%
#408045000000
1!
1%
#408050000000
0!
0%
#408055000000
1!
1%
#408060000000
0!
0%
#408065000000
1!
1%
#408070000000
0!
0%
#408075000000
1!
1%
#408080000000
0!
0%
#408085000000
1!
1%
#408090000000
0!
0%
#408095000000
1!
1%
#408100000000
0!
0%
#408105000000
1!
1%
#408110000000
0!
0%
#408115000000
1!
1%
#408120000000
0!
0%
#408125000000
1!
1%
#408130000000
0!
0%
#408135000000
1!
1%
#408140000000
0!
0%
#408145000000
1!
1%
#408150000000
0!
0%
#408155000000
1!
1%
#408160000000
0!
0%
#408165000000
1!
1%
#408170000000
0!
0%
#408175000000
1!
1%
#408180000000
0!
0%
#408185000000
1!
1%
#408190000000
0!
0%
#408195000000
1!
1%
#408200000000
0!
0%
#408205000000
1!
1%
#408210000000
0!
0%
#408215000000
1!
1%
#408220000000
0!
0%
#408225000000
1!
1%
#408230000000
0!
0%
#408235000000
1!
1%
#408240000000
0!
0%
#408245000000
1!
1%
#408250000000
0!
0%
#408255000000
1!
1%
#408260000000
0!
0%
#408265000000
1!
1%
#408270000000
0!
0%
#408275000000
1!
1%
#408280000000
0!
0%
#408285000000
1!
1%
#408290000000
0!
0%
#408295000000
1!
1%
#408300000000
0!
0%
#408305000000
1!
1%
#408310000000
0!
0%
#408315000000
1!
1%
#408320000000
0!
0%
#408325000000
1!
1%
#408330000000
0!
0%
#408335000000
1!
1%
#408340000000
0!
0%
#408345000000
1!
1%
#408350000000
0!
0%
#408355000000
1!
1%
#408360000000
0!
0%
#408365000000
1!
1%
#408370000000
0!
0%
#408375000000
1!
1%
#408380000000
0!
0%
#408385000000
1!
1%
#408390000000
0!
0%
#408395000000
1!
1%
#408400000000
0!
0%
#408405000000
1!
1%
#408410000000
0!
0%
#408415000000
1!
1%
#408420000000
0!
0%
#408425000000
1!
1%
#408430000000
0!
0%
#408435000000
1!
1%
#408440000000
0!
0%
#408445000000
1!
1%
#408450000000
0!
0%
#408455000000
1!
1%
#408460000000
0!
0%
#408465000000
1!
1%
#408470000000
0!
0%
#408475000000
1!
1%
#408480000000
0!
0%
#408485000000
1!
1%
#408490000000
0!
0%
#408495000000
1!
1%
#408500000000
0!
0%
#408505000000
1!
1%
#408510000000
0!
0%
#408515000000
1!
1%
#408520000000
0!
0%
#408525000000
1!
1%
#408530000000
0!
0%
#408535000000
1!
1%
#408540000000
0!
0%
#408545000000
1!
1%
#408550000000
0!
0%
#408555000000
1!
1%
#408560000000
0!
0%
#408565000000
1!
1%
#408570000000
0!
0%
#408575000000
1!
1%
#408580000000
0!
0%
#408585000000
1!
1%
#408590000000
0!
0%
#408595000000
1!
1%
#408600000000
0!
0%
#408605000000
1!
1%
#408610000000
0!
0%
#408615000000
1!
1%
#408620000000
0!
0%
#408625000000
1!
1%
#408630000000
0!
0%
#408635000000
1!
1%
#408640000000
0!
0%
#408645000000
1!
1%
#408650000000
0!
0%
#408655000000
1!
1%
#408660000000
0!
0%
#408665000000
1!
1%
#408670000000
0!
0%
#408675000000
1!
1%
#408680000000
0!
0%
#408685000000
1!
1%
#408690000000
0!
0%
#408695000000
1!
1%
#408700000000
0!
0%
#408705000000
1!
1%
#408710000000
0!
0%
#408715000000
1!
1%
#408720000000
0!
0%
#408725000000
1!
1%
#408730000000
0!
0%
#408735000000
1!
1%
#408740000000
0!
0%
#408745000000
1!
1%
#408750000000
0!
0%
#408755000000
1!
1%
#408760000000
0!
0%
#408765000000
1!
1%
#408770000000
0!
0%
#408775000000
1!
1%
#408780000000
0!
0%
#408785000000
1!
1%
#408790000000
0!
0%
#408795000000
1!
1%
#408800000000
0!
0%
#408805000000
1!
1%
#408810000000
0!
0%
#408815000000
1!
1%
#408820000000
0!
0%
#408825000000
1!
1%
#408830000000
0!
0%
#408835000000
1!
1%
#408840000000
0!
0%
#408845000000
1!
1%
#408850000000
0!
0%
#408855000000
1!
1%
#408860000000
0!
0%
#408865000000
1!
1%
#408870000000
0!
0%
#408875000000
1!
1%
#408880000000
0!
0%
#408885000000
1!
1%
#408890000000
0!
0%
#408895000000
1!
1%
#408900000000
0!
0%
#408905000000
1!
1%
#408910000000
0!
0%
#408915000000
1!
1%
#408920000000
0!
0%
#408925000000
1!
1%
#408930000000
0!
0%
#408935000000
1!
1%
#408940000000
0!
0%
#408945000000
1!
1%
#408950000000
0!
0%
#408955000000
1!
1%
#408960000000
0!
0%
#408965000000
1!
1%
#408970000000
0!
0%
#408975000000
1!
1%
#408980000000
0!
0%
#408985000000
1!
1%
#408990000000
0!
0%
#408995000000
1!
1%
#409000000000
0!
0%
#409005000000
1!
1%
#409010000000
0!
0%
#409015000000
1!
1%
#409020000000
0!
0%
#409025000000
1!
1%
#409030000000
0!
0%
#409035000000
1!
1%
#409040000000
0!
0%
#409045000000
1!
1%
#409050000000
0!
0%
#409055000000
1!
1%
#409060000000
0!
0%
#409065000000
1!
1%
#409070000000
0!
0%
#409075000000
1!
1%
#409080000000
0!
0%
#409085000000
1!
1%
#409090000000
0!
0%
#409095000000
1!
1%
#409100000000
0!
0%
#409105000000
1!
1%
#409110000000
0!
0%
#409115000000
1!
1%
#409120000000
0!
0%
#409125000000
1!
1%
#409130000000
0!
0%
#409135000000
1!
1%
#409140000000
0!
0%
#409145000000
1!
1%
#409150000000
0!
0%
#409155000000
1!
1%
#409160000000
0!
0%
#409165000000
1!
1%
#409170000000
0!
0%
#409175000000
1!
1%
#409180000000
0!
0%
#409185000000
1!
1%
#409190000000
0!
0%
#409195000000
1!
1%
#409200000000
0!
0%
#409205000000
1!
1%
#409210000000
0!
0%
#409215000000
1!
1%
#409220000000
0!
0%
#409225000000
1!
1%
#409230000000
0!
0%
#409235000000
1!
1%
#409240000000
0!
0%
#409245000000
1!
1%
#409250000000
0!
0%
#409255000000
1!
1%
#409260000000
0!
0%
#409265000000
1!
1%
#409270000000
0!
0%
#409275000000
1!
1%
#409280000000
0!
0%
#409285000000
1!
1%
#409290000000
0!
0%
#409295000000
1!
1%
#409300000000
0!
0%
#409305000000
1!
1%
#409310000000
0!
0%
#409315000000
1!
1%
#409320000000
0!
0%
#409325000000
1!
1%
#409330000000
0!
0%
#409335000000
1!
1%
#409340000000
0!
0%
#409345000000
1!
1%
#409350000000
0!
0%
#409355000000
1!
1%
#409360000000
0!
0%
#409365000000
1!
1%
#409370000000
0!
0%
#409375000000
1!
1%
#409380000000
0!
0%
#409385000000
1!
1%
#409390000000
0!
0%
#409395000000
1!
1%
#409400000000
0!
0%
#409405000000
1!
1%
#409410000000
0!
0%
#409415000000
1!
1%
#409420000000
0!
0%
#409425000000
1!
1%
#409430000000
0!
0%
#409435000000
1!
1%
#409440000000
0!
0%
#409445000000
1!
1%
#409450000000
0!
0%
#409455000000
1!
1%
#409460000000
0!
0%
#409465000000
1!
1%
#409470000000
0!
0%
#409475000000
1!
1%
#409480000000
0!
0%
#409485000000
1!
1%
#409490000000
0!
0%
#409495000000
1!
1%
#409500000000
0!
0%
#409505000000
1!
1%
#409510000000
0!
0%
#409515000000
1!
1%
#409520000000
0!
0%
#409525000000
1!
1%
#409530000000
0!
0%
#409535000000
1!
1%
#409540000000
0!
0%
#409545000000
1!
1%
#409550000000
0!
0%
#409555000000
1!
1%
#409560000000
0!
0%
#409565000000
1!
1%
#409570000000
0!
0%
#409575000000
1!
1%
#409580000000
0!
0%
#409585000000
1!
1%
#409590000000
0!
0%
#409595000000
1!
1%
#409600000000
0!
0%
#409605000000
1!
1%
#409610000000
0!
0%
#409615000000
1!
1%
#409620000000
0!
0%
#409625000000
1!
1%
#409630000000
0!
0%
#409635000000
1!
1%
#409640000000
0!
0%
#409645000000
1!
1%
#409650000000
0!
0%
#409655000000
1!
1%
#409660000000
0!
0%
#409665000000
1!
1%
#409670000000
0!
0%
#409675000000
1!
1%
#409680000000
0!
0%
#409685000000
1!
1%
#409690000000
0!
0%
#409695000000
1!
1%
#409700000000
0!
0%
#409705000000
1!
1%
#409710000000
0!
0%
#409715000000
1!
1%
#409720000000
0!
0%
#409725000000
1!
1%
#409730000000
0!
0%
#409735000000
1!
1%
#409740000000
0!
0%
#409745000000
1!
1%
#409750000000
0!
0%
#409755000000
1!
1%
#409760000000
0!
0%
#409765000000
1!
1%
#409770000000
0!
0%
#409775000000
1!
1%
#409780000000
0!
0%
#409785000000
1!
1%
#409790000000
0!
0%
#409795000000
1!
1%
#409800000000
0!
0%
#409805000000
1!
1%
#409810000000
0!
0%
#409815000000
1!
1%
#409820000000
0!
0%
#409825000000
1!
1%
#409830000000
0!
0%
#409835000000
1!
1%
#409840000000
0!
0%
#409845000000
1!
1%
#409850000000
0!
0%
#409855000000
1!
1%
#409860000000
0!
0%
#409865000000
1!
1%
#409870000000
0!
0%
#409875000000
1!
1%
#409880000000
0!
0%
#409885000000
1!
1%
#409890000000
0!
0%
#409895000000
1!
1%
#409900000000
0!
0%
#409905000000
1!
1%
#409910000000
0!
0%
#409915000000
1!
1%
#409920000000
0!
0%
#409925000000
1!
1%
#409930000000
0!
0%
#409935000000
1!
1%
#409940000000
0!
0%
#409945000000
1!
1%
#409950000000
0!
0%
#409955000000
1!
1%
#409960000000
0!
0%
#409965000000
1!
1%
#409970000000
0!
0%
#409975000000
1!
1%
#409980000000
0!
0%
#409985000000
1!
1%
#409990000000
0!
0%
#409995000000
1!
1%
#410000000000
0!
0%
#410005000000
1!
1%
#410010000000
0!
0%
#410015000000
1!
1%
#410020000000
0!
0%
#410025000000
1!
1%
#410030000000
0!
0%
#410035000000
1!
1%
#410040000000
0!
0%
#410045000000
1!
1%
#410050000000
0!
0%
#410055000000
1!
1%
#410060000000
0!
0%
#410065000000
1!
1%
#410070000000
0!
0%
#410075000000
1!
1%
#410080000000
0!
0%
#410085000000
1!
1%
#410090000000
0!
0%
#410095000000
1!
1%
#410100000000
0!
0%
#410105000000
1!
1%
#410110000000
0!
0%
#410115000000
1!
1%
#410120000000
0!
0%
#410125000000
1!
1%
#410130000000
0!
0%
#410135000000
1!
1%
#410140000000
0!
0%
#410145000000
1!
1%
#410150000000
0!
0%
#410155000000
1!
1%
#410160000000
0!
0%
#410165000000
1!
1%
#410170000000
0!
0%
#410175000000
1!
1%
#410180000000
0!
0%
#410185000000
1!
1%
#410190000000
0!
0%
#410195000000
1!
1%
#410200000000
0!
0%
#410205000000
1!
1%
#410210000000
0!
0%
#410215000000
1!
1%
#410220000000
0!
0%
#410225000000
1!
1%
#410230000000
0!
0%
#410235000000
1!
1%
#410240000000
0!
0%
#410245000000
1!
1%
#410250000000
0!
0%
#410255000000
1!
1%
#410260000000
0!
0%
#410265000000
1!
1%
#410270000000
0!
0%
#410275000000
1!
1%
#410280000000
0!
0%
#410285000000
1!
1%
#410290000000
0!
0%
#410295000000
1!
1%
#410300000000
0!
0%
#410305000000
1!
1%
#410310000000
0!
0%
#410315000000
1!
1%
#410320000000
0!
0%
#410325000000
1!
1%
#410330000000
0!
0%
#410335000000
1!
1%
#410340000000
0!
0%
#410345000000
1!
1%
#410350000000
0!
0%
#410355000000
1!
1%
#410360000000
0!
0%
#410365000000
1!
1%
#410370000000
0!
0%
#410375000000
1!
1%
#410380000000
0!
0%
#410385000000
1!
1%
#410390000000
0!
0%
#410395000000
1!
1%
#410400000000
0!
0%
#410405000000
1!
1%
#410410000000
0!
0%
#410415000000
1!
1%
#410420000000
0!
0%
#410425000000
1!
1%
#410430000000
0!
0%
#410435000000
1!
1%
#410440000000
0!
0%
#410445000000
1!
1%
#410450000000
0!
0%
#410455000000
1!
1%
#410460000000
0!
0%
#410465000000
1!
1%
#410470000000
0!
0%
#410475000000
1!
1%
#410480000000
0!
0%
#410485000000
1!
1%
#410490000000
0!
0%
#410495000000
1!
1%
#410500000000
0!
0%
#410505000000
1!
1%
#410510000000
0!
0%
#410515000000
1!
1%
#410520000000
0!
0%
#410525000000
1!
1%
#410530000000
0!
0%
#410535000000
1!
1%
#410540000000
0!
0%
#410545000000
1!
1%
#410550000000
0!
0%
#410555000000
1!
1%
#410560000000
0!
0%
#410565000000
1!
1%
#410570000000
0!
0%
#410575000000
1!
1%
#410580000000
0!
0%
#410585000000
1!
1%
#410590000000
0!
0%
#410595000000
1!
1%
#410600000000
0!
0%
#410605000000
1!
1%
#410610000000
0!
0%
#410615000000
1!
1%
#410620000000
0!
0%
#410625000000
1!
1%
#410630000000
0!
0%
#410635000000
1!
1%
#410640000000
0!
0%
#410645000000
1!
1%
#410650000000
0!
0%
#410655000000
1!
1%
#410660000000
0!
0%
#410665000000
1!
1%
#410670000000
0!
0%
#410675000000
1!
1%
#410680000000
0!
0%
#410685000000
1!
1%
#410690000000
0!
0%
#410695000000
1!
1%
#410700000000
0!
0%
#410705000000
1!
1%
#410710000000
0!
0%
#410715000000
1!
1%
#410720000000
0!
0%
#410725000000
1!
1%
#410730000000
0!
0%
#410735000000
1!
1%
#410740000000
0!
0%
#410745000000
1!
1%
#410750000000
0!
0%
#410755000000
1!
1%
#410760000000
0!
0%
#410765000000
1!
1%
#410770000000
0!
0%
#410775000000
1!
1%
#410780000000
0!
0%
#410785000000
1!
1%
#410790000000
0!
0%
#410795000000
1!
1%
#410800000000
0!
0%
#410805000000
1!
1%
#410810000000
0!
0%
#410815000000
1!
1%
#410820000000
0!
0%
#410825000000
1!
1%
#410830000000
0!
0%
#410835000000
1!
1%
#410840000000
0!
0%
#410845000000
1!
1%
#410850000000
0!
0%
#410855000000
1!
1%
#410860000000
0!
0%
#410865000000
1!
1%
#410870000000
0!
0%
#410875000000
1!
1%
#410880000000
0!
0%
#410885000000
1!
1%
#410890000000
0!
0%
#410895000000
1!
1%
#410900000000
0!
0%
#410905000000
1!
1%
#410910000000
0!
0%
#410915000000
1!
1%
#410920000000
0!
0%
#410925000000
1!
1%
#410930000000
0!
0%
#410935000000
1!
1%
#410940000000
0!
0%
#410945000000
1!
1%
#410950000000
0!
0%
#410955000000
1!
1%
#410960000000
0!
0%
#410965000000
1!
1%
#410970000000
0!
0%
#410975000000
1!
1%
#410980000000
0!
0%
#410985000000
1!
1%
#410990000000
0!
0%
#410995000000
1!
1%
#411000000000
0!
0%
#411005000000
1!
1%
#411010000000
0!
0%
#411015000000
1!
1%
#411020000000
0!
0%
#411025000000
1!
1%
#411030000000
0!
0%
#411035000000
1!
1%
#411040000000
0!
0%
#411045000000
1!
1%
#411050000000
0!
0%
#411055000000
1!
1%
#411060000000
0!
0%
#411065000000
1!
1%
#411070000000
0!
0%
#411075000000
1!
1%
#411080000000
0!
0%
#411085000000
1!
1%
#411090000000
0!
0%
#411095000000
1!
1%
#411100000000
0!
0%
#411105000000
1!
1%
#411110000000
0!
0%
#411115000000
1!
1%
#411120000000
0!
0%
#411125000000
1!
1%
#411130000000
0!
0%
#411135000000
1!
1%
#411140000000
0!
0%
#411145000000
1!
1%
#411150000000
0!
0%
#411155000000
1!
1%
#411160000000
0!
0%
#411165000000
1!
1%
#411170000000
0!
0%
#411175000000
1!
1%
#411180000000
0!
0%
#411185000000
1!
1%
#411190000000
0!
0%
#411195000000
1!
1%
#411200000000
0!
0%
#411205000000
1!
1%
#411210000000
0!
0%
#411215000000
1!
1%
#411220000000
0!
0%
#411225000000
1!
1%
#411230000000
0!
0%
#411235000000
1!
1%
#411240000000
0!
0%
#411245000000
1!
1%
#411250000000
0!
0%
#411255000000
1!
1%
#411260000000
0!
0%
#411265000000
1!
1%
#411270000000
0!
0%
#411275000000
1!
1%
#411280000000
0!
0%
#411285000000
1!
1%
#411290000000
0!
0%
#411295000000
1!
1%
#411300000000
0!
0%
#411305000000
1!
1%
#411310000000
0!
0%
#411315000000
1!
1%
#411320000000
0!
0%
#411325000000
1!
1%
#411330000000
0!
0%
#411335000000
1!
1%
#411340000000
0!
0%
#411345000000
1!
1%
#411350000000
0!
0%
#411355000000
1!
1%
#411360000000
0!
0%
#411365000000
1!
1%
#411370000000
0!
0%
#411375000000
1!
1%
#411380000000
0!
0%
#411385000000
1!
1%
#411390000000
0!
0%
#411395000000
1!
1%
#411400000000
0!
0%
#411405000000
1!
1%
#411410000000
0!
0%
#411415000000
1!
1%
#411420000000
0!
0%
#411425000000
1!
1%
#411430000000
0!
0%
#411435000000
1!
1%
#411440000000
0!
0%
#411445000000
1!
1%
#411450000000
0!
0%
#411455000000
1!
1%
#411460000000
0!
0%
#411465000000
1!
1%
#411470000000
0!
0%
#411475000000
1!
1%
#411480000000
0!
0%
#411485000000
1!
1%
#411490000000
0!
0%
#411495000000
1!
1%
#411500000000
0!
0%
#411505000000
1!
1%
#411510000000
0!
0%
#411515000000
1!
1%
#411520000000
0!
0%
#411525000000
1!
1%
#411530000000
0!
0%
#411535000000
1!
1%
#411540000000
0!
0%
#411545000000
1!
1%
#411550000000
0!
0%
#411555000000
1!
1%
#411560000000
0!
0%
#411565000000
1!
1%
#411570000000
0!
0%
#411575000000
1!
1%
#411580000000
0!
0%
#411585000000
1!
1%
#411590000000
0!
0%
#411595000000
1!
1%
#411600000000
0!
0%
#411605000000
1!
1%
#411610000000
0!
0%
#411615000000
1!
1%
#411620000000
0!
0%
#411625000000
1!
1%
#411630000000
0!
0%
#411635000000
1!
1%
#411640000000
0!
0%
#411645000000
1!
1%
#411650000000
0!
0%
#411655000000
1!
1%
#411660000000
0!
0%
#411665000000
1!
1%
#411670000000
0!
0%
#411675000000
1!
1%
#411680000000
0!
0%
#411685000000
1!
1%
#411690000000
0!
0%
#411695000000
1!
1%
#411700000000
0!
0%
#411705000000
1!
1%
#411710000000
0!
0%
#411715000000
1!
1%
#411720000000
0!
0%
#411725000000
1!
1%
#411730000000
0!
0%
#411735000000
1!
1%
#411740000000
0!
0%
#411745000000
1!
1%
#411750000000
0!
0%
#411755000000
1!
1%
#411760000000
0!
0%
#411765000000
1!
1%
#411770000000
0!
0%
#411775000000
1!
1%
#411780000000
0!
0%
#411785000000
1!
1%
#411790000000
0!
0%
#411795000000
1!
1%
#411800000000
0!
0%
#411805000000
1!
1%
#411810000000
0!
0%
#411815000000
1!
1%
#411820000000
0!
0%
#411825000000
1!
1%
#411830000000
0!
0%
#411835000000
1!
1%
#411840000000
0!
0%
#411845000000
1!
1%
#411850000000
0!
0%
#411855000000
1!
1%
#411860000000
0!
0%
#411865000000
1!
1%
#411870000000
0!
0%
#411875000000
1!
1%
#411880000000
0!
0%
#411885000000
1!
1%
#411890000000
0!
0%
#411895000000
1!
1%
#411900000000
0!
0%
#411905000000
1!
1%
#411910000000
0!
0%
#411915000000
1!
1%
#411920000000
0!
0%
#411925000000
1!
1%
#411930000000
0!
0%
#411935000000
1!
1%
#411940000000
0!
0%
#411945000000
1!
1%
#411950000000
0!
0%
#411955000000
1!
1%
#411960000000
0!
0%
#411965000000
1!
1%
#411970000000
0!
0%
#411975000000
1!
1%
#411980000000
0!
0%
#411985000000
1!
1%
#411990000000
0!
0%
#411995000000
1!
1%
#412000000000
0!
0%
#412005000000
1!
1%
#412010000000
0!
0%
#412015000000
1!
1%
#412020000000
0!
0%
#412025000000
1!
1%
#412030000000
0!
0%
#412035000000
1!
1%
#412040000000
0!
0%
#412045000000
1!
1%
#412050000000
0!
0%
#412055000000
1!
1%
#412060000000
0!
0%
#412065000000
1!
1%
#412070000000
0!
0%
#412075000000
1!
1%
#412080000000
0!
0%
#412085000000
1!
1%
#412090000000
0!
0%
#412095000000
1!
1%
#412100000000
0!
0%
#412105000000
1!
1%
#412110000000
0!
0%
#412115000000
1!
1%
#412120000000
0!
0%
#412125000000
1!
1%
#412130000000
0!
0%
#412135000000
1!
1%
#412140000000
0!
0%
#412145000000
1!
1%
#412150000000
0!
0%
#412155000000
1!
1%
#412160000000
0!
0%
#412165000000
1!
1%
#412170000000
0!
0%
#412175000000
1!
1%
#412180000000
0!
0%
#412185000000
1!
1%
#412190000000
0!
0%
#412195000000
1!
1%
#412200000000
0!
0%
#412205000000
1!
1%
#412210000000
0!
0%
#412215000000
1!
1%
#412220000000
0!
0%
#412225000000
1!
1%
#412230000000
0!
0%
#412235000000
1!
1%
#412240000000
0!
0%
#412245000000
1!
1%
#412250000000
0!
0%
#412255000000
1!
1%
#412260000000
0!
0%
#412265000000
1!
1%
#412270000000
0!
0%
#412275000000
1!
1%
#412280000000
0!
0%
#412285000000
1!
1%
#412290000000
0!
0%
#412295000000
1!
1%
#412300000000
0!
0%
#412305000000
1!
1%
#412310000000
0!
0%
#412315000000
1!
1%
#412320000000
0!
0%
#412325000000
1!
1%
#412330000000
0!
0%
#412335000000
1!
1%
#412340000000
0!
0%
#412345000000
1!
1%
#412350000000
0!
0%
#412355000000
1!
1%
#412360000000
0!
0%
#412365000000
1!
1%
#412370000000
0!
0%
#412375000000
1!
1%
#412380000000
0!
0%
#412385000000
1!
1%
#412390000000
0!
0%
#412395000000
1!
1%
#412400000000
0!
0%
#412405000000
1!
1%
#412410000000
0!
0%
#412415000000
1!
1%
#412420000000
0!
0%
#412425000000
1!
1%
#412430000000
0!
0%
#412435000000
1!
1%
#412440000000
0!
0%
#412445000000
1!
1%
#412450000000
0!
0%
#412455000000
1!
1%
#412460000000
0!
0%
#412465000000
1!
1%
#412470000000
0!
0%
#412475000000
1!
1%
#412480000000
0!
0%
#412485000000
1!
1%
#412490000000
0!
0%
#412495000000
1!
1%
#412500000000
0!
0%
#412505000000
1!
1%
#412510000000
0!
0%
#412515000000
1!
1%
#412520000000
0!
0%
#412525000000
1!
1%
#412530000000
0!
0%
#412535000000
1!
1%
#412540000000
0!
0%
#412545000000
1!
1%
#412550000000
0!
0%
#412555000000
1!
1%
#412560000000
0!
0%
#412565000000
1!
1%
#412570000000
0!
0%
#412575000000
1!
1%
#412580000000
0!
0%
#412585000000
1!
1%
#412590000000
0!
0%
#412595000000
1!
1%
#412600000000
0!
0%
#412605000000
1!
1%
#412610000000
0!
0%
#412615000000
1!
1%
#412620000000
0!
0%
#412625000000
1!
1%
#412630000000
0!
0%
#412635000000
1!
1%
#412640000000
0!
0%
#412645000000
1!
1%
#412650000000
0!
0%
#412655000000
1!
1%
#412660000000
0!
0%
#412665000000
1!
1%
#412670000000
0!
0%
#412675000000
1!
1%
#412680000000
0!
0%
#412685000000
1!
1%
#412690000000
0!
0%
#412695000000
1!
1%
#412700000000
0!
0%
#412705000000
1!
1%
#412710000000
0!
0%
#412715000000
1!
1%
#412720000000
0!
0%
#412725000000
1!
1%
#412730000000
0!
0%
#412735000000
1!
1%
#412740000000
0!
0%
#412745000000
1!
1%
#412750000000
0!
0%
#412755000000
1!
1%
#412760000000
0!
0%
#412765000000
1!
1%
#412770000000
0!
0%
#412775000000
1!
1%
#412780000000
0!
0%
#412785000000
1!
1%
#412790000000
0!
0%
#412795000000
1!
1%
#412800000000
0!
0%
#412805000000
1!
1%
#412810000000
0!
0%
#412815000000
1!
1%
#412820000000
0!
0%
#412825000000
1!
1%
#412830000000
0!
0%
#412835000000
1!
1%
#412840000000
0!
0%
#412845000000
1!
1%
#412850000000
0!
0%
#412855000000
1!
1%
#412860000000
0!
0%
#412865000000
1!
1%
#412870000000
0!
0%
#412875000000
1!
1%
#412880000000
0!
0%
#412885000000
1!
1%
#412890000000
0!
0%
#412895000000
1!
1%
#412900000000
0!
0%
#412905000000
1!
1%
#412910000000
0!
0%
#412915000000
1!
1%
#412920000000
0!
0%
#412925000000
1!
1%
#412930000000
0!
0%
#412935000000
1!
1%
#412940000000
0!
0%
#412945000000
1!
1%
#412950000000
0!
0%
#412955000000
1!
1%
#412960000000
0!
0%
#412965000000
1!
1%
#412970000000
0!
0%
#412975000000
1!
1%
#412980000000
0!
0%
#412985000000
1!
1%
#412990000000
0!
0%
#412995000000
1!
1%
#413000000000
0!
0%
#413005000000
1!
1%
#413010000000
0!
0%
#413015000000
1!
1%
#413020000000
0!
0%
#413025000000
1!
1%
#413030000000
0!
0%
#413035000000
1!
1%
#413040000000
0!
0%
#413045000000
1!
1%
#413050000000
0!
0%
#413055000000
1!
1%
#413060000000
0!
0%
#413065000000
1!
1%
#413070000000
0!
0%
#413075000000
1!
1%
#413080000000
0!
0%
#413085000000
1!
1%
#413090000000
0!
0%
#413095000000
1!
1%
#413100000000
0!
0%
#413105000000
1!
1%
#413110000000
0!
0%
#413115000000
1!
1%
#413120000000
0!
0%
#413125000000
1!
1%
#413130000000
0!
0%
#413135000000
1!
1%
#413140000000
0!
0%
#413145000000
1!
1%
#413150000000
0!
0%
#413155000000
1!
1%
#413160000000
0!
0%
#413165000000
1!
1%
#413170000000
0!
0%
#413175000000
1!
1%
#413180000000
0!
0%
#413185000000
1!
1%
#413190000000
0!
0%
#413195000000
1!
1%
#413200000000
0!
0%
#413205000000
1!
1%
#413210000000
0!
0%
#413215000000
1!
1%
#413220000000
0!
0%
#413225000000
1!
1%
#413230000000
0!
0%
#413235000000
1!
1%
#413240000000
0!
0%
#413245000000
1!
1%
#413250000000
0!
0%
#413255000000
1!
1%
#413260000000
0!
0%
#413265000000
1!
1%
#413270000000
0!
0%
#413275000000
1!
1%
#413280000000
0!
0%
#413285000000
1!
1%
#413290000000
0!
0%
#413295000000
1!
1%
#413300000000
0!
0%
#413305000000
1!
1%
#413310000000
0!
0%
#413315000000
1!
1%
#413320000000
0!
0%
#413325000000
1!
1%
#413330000000
0!
0%
#413335000000
1!
1%
#413340000000
0!
0%
#413345000000
1!
1%
#413350000000
0!
0%
#413355000000
1!
1%
#413360000000
0!
0%
#413365000000
1!
1%
#413370000000
0!
0%
#413375000000
1!
1%
#413380000000
0!
0%
#413385000000
1!
1%
#413390000000
0!
0%
#413395000000
1!
1%
#413400000000
0!
0%
#413405000000
1!
1%
#413410000000
0!
0%
#413415000000
1!
1%
#413420000000
0!
0%
#413425000000
1!
1%
#413430000000
0!
0%
#413435000000
1!
1%
#413440000000
0!
0%
#413445000000
1!
1%
#413450000000
0!
0%
#413455000000
1!
1%
#413460000000
0!
0%
#413465000000
1!
1%
#413470000000
0!
0%
#413475000000
1!
1%
#413480000000
0!
0%
#413485000000
1!
1%
#413490000000
0!
0%
#413495000000
1!
1%
#413500000000
0!
0%
#413505000000
1!
1%
#413510000000
0!
0%
#413515000000
1!
1%
#413520000000
0!
0%
#413525000000
1!
1%
#413530000000
0!
0%
#413535000000
1!
1%
#413540000000
0!
0%
#413545000000
1!
1%
#413550000000
0!
0%
#413555000000
1!
1%
#413560000000
0!
0%
#413565000000
1!
1%
#413570000000
0!
0%
#413575000000
1!
1%
#413580000000
0!
0%
#413585000000
1!
1%
#413590000000
0!
0%
#413595000000
1!
1%
#413600000000
0!
0%
#413605000000
1!
1%
#413610000000
0!
0%
#413615000000
1!
1%
#413620000000
0!
0%
#413625000000
1!
1%
#413630000000
0!
0%
#413635000000
1!
1%
#413640000000
0!
0%
#413645000000
1!
1%
#413650000000
0!
0%
#413655000000
1!
1%
#413660000000
0!
0%
#413665000000
1!
1%
#413670000000
0!
0%
#413675000000
1!
1%
#413680000000
0!
0%
#413685000000
1!
1%
#413690000000
0!
0%
#413695000000
1!
1%
#413700000000
0!
0%
#413705000000
1!
1%
#413710000000
0!
0%
#413715000000
1!
1%
#413720000000
0!
0%
#413725000000
1!
1%
#413730000000
0!
0%
#413735000000
1!
1%
#413740000000
0!
0%
#413745000000
1!
1%
#413750000000
0!
0%
#413755000000
1!
1%
#413760000000
0!
0%
#413765000000
1!
1%
#413770000000
0!
0%
#413775000000
1!
1%
#413780000000
0!
0%
#413785000000
1!
1%
#413790000000
0!
0%
#413795000000
1!
1%
#413800000000
0!
0%
#413805000000
1!
1%
#413810000000
0!
0%
#413815000000
1!
1%
#413820000000
0!
0%
#413825000000
1!
1%
#413830000000
0!
0%
#413835000000
1!
1%
#413840000000
0!
0%
#413845000000
1!
1%
#413850000000
0!
0%
#413855000000
1!
1%
#413860000000
0!
0%
#413865000000
1!
1%
#413870000000
0!
0%
#413875000000
1!
1%
#413880000000
0!
0%
#413885000000
1!
1%
#413890000000
0!
0%
#413895000000
1!
1%
#413900000000
0!
0%
#413905000000
1!
1%
#413910000000
0!
0%
#413915000000
1!
1%
#413920000000
0!
0%
#413925000000
1!
1%
#413930000000
0!
0%
#413935000000
1!
1%
#413940000000
0!
0%
#413945000000
1!
1%
#413950000000
0!
0%
#413955000000
1!
1%
#413960000000
0!
0%
#413965000000
1!
1%
#413970000000
0!
0%
#413975000000
1!
1%
#413980000000
0!
0%
#413985000000
1!
1%
#413990000000
0!
0%
#413995000000
1!
1%
#414000000000
0!
0%
#414005000000
1!
1%
#414010000000
0!
0%
#414015000000
1!
1%
#414020000000
0!
0%
#414025000000
1!
1%
#414030000000
0!
0%
#414035000000
1!
1%
#414040000000
0!
0%
#414045000000
1!
1%
#414050000000
0!
0%
#414055000000
1!
1%
#414060000000
0!
0%
#414065000000
1!
1%
#414070000000
0!
0%
#414075000000
1!
1%
#414080000000
0!
0%
#414085000000
1!
1%
#414090000000
0!
0%
#414095000000
1!
1%
#414100000000
0!
0%
#414105000000
1!
1%
#414110000000
0!
0%
#414115000000
1!
1%
#414120000000
0!
0%
#414125000000
1!
1%
#414130000000
0!
0%
#414135000000
1!
1%
#414140000000
0!
0%
#414145000000
1!
1%
#414150000000
0!
0%
#414155000000
1!
1%
#414160000000
0!
0%
#414165000000
1!
1%
#414170000000
0!
0%
#414175000000
1!
1%
#414180000000
0!
0%
#414185000000
1!
1%
#414190000000
0!
0%
#414195000000
1!
1%
#414200000000
0!
0%
#414205000000
1!
1%
#414210000000
0!
0%
#414215000000
1!
1%
#414220000000
0!
0%
#414225000000
1!
1%
#414230000000
0!
0%
#414235000000
1!
1%
#414240000000
0!
0%
#414245000000
1!
1%
#414250000000
0!
0%
#414255000000
1!
1%
#414260000000
0!
0%
#414265000000
1!
1%
#414270000000
0!
0%
#414275000000
1!
1%
#414280000000
0!
0%
#414285000000
1!
1%
#414290000000
0!
0%
#414295000000
1!
1%
#414300000000
0!
0%
#414305000000
1!
1%
#414310000000
0!
0%
#414315000000
1!
1%
#414320000000
0!
0%
#414325000000
1!
1%
#414330000000
0!
0%
#414335000000
1!
1%
#414340000000
0!
0%
#414345000000
1!
1%
#414350000000
0!
0%
#414355000000
1!
1%
#414360000000
0!
0%
#414365000000
1!
1%
#414370000000
0!
0%
#414375000000
1!
1%
#414380000000
0!
0%
#414385000000
1!
1%
#414390000000
0!
0%
#414395000000
1!
1%
#414400000000
0!
0%
#414405000000
1!
1%
#414410000000
0!
0%
#414415000000
1!
1%
#414420000000
0!
0%
#414425000000
1!
1%
#414430000000
0!
0%
#414435000000
1!
1%
#414440000000
0!
0%
#414445000000
1!
1%
#414450000000
0!
0%
#414455000000
1!
1%
#414460000000
0!
0%
#414465000000
1!
1%
#414470000000
0!
0%
#414475000000
1!
1%
#414480000000
0!
0%
#414485000000
1!
1%
#414490000000
0!
0%
#414495000000
1!
1%
#414500000000
0!
0%
#414505000000
1!
1%
#414510000000
0!
0%
#414515000000
1!
1%
#414520000000
0!
0%
#414525000000
1!
1%
#414530000000
0!
0%
#414535000000
1!
1%
#414540000000
0!
0%
#414545000000
1!
1%
#414550000000
0!
0%
#414555000000
1!
1%
#414560000000
0!
0%
#414565000000
1!
1%
#414570000000
0!
0%
#414575000000
1!
1%
#414580000000
0!
0%
#414585000000
1!
1%
#414590000000
0!
0%
#414595000000
1!
1%
#414600000000
0!
0%
#414605000000
1!
1%
#414610000000
0!
0%
#414615000000
1!
1%
#414620000000
0!
0%
#414625000000
1!
1%
#414630000000
0!
0%
#414635000000
1!
1%
#414640000000
0!
0%
#414645000000
1!
1%
#414650000000
0!
0%
#414655000000
1!
1%
#414660000000
0!
0%
#414665000000
1!
1%
#414670000000
0!
0%
#414675000000
1!
1%
#414680000000
0!
0%
#414685000000
1!
1%
#414690000000
0!
0%
#414695000000
1!
1%
#414700000000
0!
0%
#414705000000
1!
1%
#414710000000
0!
0%
#414715000000
1!
1%
#414720000000
0!
0%
#414725000000
1!
1%
#414730000000
0!
0%
#414735000000
1!
1%
#414740000000
0!
0%
#414745000000
1!
1%
#414750000000
0!
0%
#414755000000
1!
1%
#414760000000
0!
0%
#414765000000
1!
1%
#414770000000
0!
0%
#414775000000
1!
1%
#414780000000
0!
0%
#414785000000
1!
1%
#414790000000
0!
0%
#414795000000
1!
1%
#414800000000
0!
0%
#414805000000
1!
1%
#414810000000
0!
0%
#414815000000
1!
1%
#414820000000
0!
0%
#414825000000
1!
1%
#414830000000
0!
0%
#414835000000
1!
1%
#414840000000
0!
0%
#414845000000
1!
1%
#414850000000
0!
0%
#414855000000
1!
1%
#414860000000
0!
0%
#414865000000
1!
1%
#414870000000
0!
0%
#414875000000
1!
1%
#414880000000
0!
0%
#414885000000
1!
1%
#414890000000
0!
0%
#414895000000
1!
1%
#414900000000
0!
0%
#414905000000
1!
1%
#414910000000
0!
0%
#414915000000
1!
1%
#414920000000
0!
0%
#414925000000
1!
1%
#414930000000
0!
0%
#414935000000
1!
1%
#414940000000
0!
0%
#414945000000
1!
1%
#414950000000
0!
0%
#414955000000
1!
1%
#414960000000
0!
0%
#414965000000
1!
1%
#414970000000
0!
0%
#414975000000
1!
1%
#414980000000
0!
0%
#414985000000
1!
1%
#414990000000
0!
0%
#414995000000
1!
1%
#415000000000
0!
0%
#415005000000
1!
1%
#415010000000
0!
0%
#415015000000
1!
1%
#415020000000
0!
0%
#415025000000
1!
1%
#415030000000
0!
0%
#415035000000
1!
1%
#415040000000
0!
0%
#415045000000
1!
1%
#415050000000
0!
0%
#415055000000
1!
1%
#415060000000
0!
0%
#415065000000
1!
1%
#415070000000
0!
0%
#415075000000
1!
1%
#415080000000
0!
0%
#415085000000
1!
1%
#415090000000
0!
0%
#415095000000
1!
1%
#415100000000
0!
0%
#415105000000
1!
1%
#415110000000
0!
0%
#415115000000
1!
1%
#415120000000
0!
0%
#415125000000
1!
1%
#415130000000
0!
0%
#415135000000
1!
1%
#415140000000
0!
0%
#415145000000
1!
1%
#415150000000
0!
0%
#415155000000
1!
1%
#415160000000
0!
0%
#415165000000
1!
1%
#415170000000
0!
0%
#415175000000
1!
1%
#415180000000
0!
0%
#415185000000
1!
1%
#415190000000
0!
0%
#415195000000
1!
1%
#415200000000
0!
0%
#415205000000
1!
1%
#415210000000
0!
0%
#415215000000
1!
1%
#415220000000
0!
0%
#415225000000
1!
1%
#415230000000
0!
0%
#415235000000
1!
1%
#415240000000
0!
0%
#415245000000
1!
1%
#415250000000
0!
0%
#415255000000
1!
1%
#415260000000
0!
0%
#415265000000
1!
1%
#415270000000
0!
0%
#415275000000
1!
1%
#415280000000
0!
0%
#415285000000
1!
1%
#415290000000
0!
0%
#415295000000
1!
1%
#415300000000
0!
0%
#415305000000
1!
1%
#415310000000
0!
0%
#415315000000
1!
1%
#415320000000
0!
0%
#415325000000
1!
1%
#415330000000
0!
0%
#415335000000
1!
1%
#415340000000
0!
0%
#415345000000
1!
1%
#415350000000
0!
0%
#415355000000
1!
1%
#415360000000
0!
0%
#415365000000
1!
1%
#415370000000
0!
0%
#415375000000
1!
1%
#415380000000
0!
0%
#415385000000
1!
1%
#415390000000
0!
0%
#415395000000
1!
1%
#415400000000
0!
0%
#415405000000
1!
1%
#415410000000
0!
0%
#415415000000
1!
1%
#415420000000
0!
0%
#415425000000
1!
1%
#415430000000
0!
0%
#415435000000
1!
1%
#415440000000
0!
0%
#415445000000
1!
1%
#415450000000
0!
0%
#415455000000
1!
1%
#415460000000
0!
0%
#415465000000
1!
1%
#415470000000
0!
0%
#415475000000
1!
1%
#415480000000
0!
0%
#415485000000
1!
1%
#415490000000
0!
0%
#415495000000
1!
1%
#415500000000
0!
0%
#415505000000
1!
1%
#415510000000
0!
0%
#415515000000
1!
1%
#415520000000
0!
0%
#415525000000
1!
1%
#415530000000
0!
0%
#415535000000
1!
1%
#415540000000
0!
0%
#415545000000
1!
1%
#415550000000
0!
0%
#415555000000
1!
1%
#415560000000
0!
0%
#415565000000
1!
1%
#415570000000
0!
0%
#415575000000
1!
1%
#415580000000
0!
0%
#415585000000
1!
1%
#415590000000
0!
0%
#415595000000
1!
1%
#415600000000
0!
0%
#415605000000
1!
1%
#415610000000
0!
0%
#415615000000
1!
1%
#415620000000
0!
0%
#415625000000
1!
1%
#415630000000
0!
0%
#415635000000
1!
1%
#415640000000
0!
0%
#415645000000
1!
1%
#415650000000
0!
0%
#415655000000
1!
1%
#415660000000
0!
0%
#415665000000
1!
1%
#415670000000
0!
0%
#415675000000
1!
1%
#415680000000
0!
0%
#415685000000
1!
1%
#415690000000
0!
0%
#415695000000
1!
1%
#415700000000
0!
0%
#415705000000
1!
1%
#415710000000
0!
0%
#415715000000
1!
1%
#415720000000
0!
0%
#415725000000
1!
1%
#415730000000
0!
0%
#415735000000
1!
1%
#415740000000
0!
0%
#415745000000
1!
1%
#415750000000
0!
0%
#415755000000
1!
1%
#415760000000
0!
0%
#415765000000
1!
1%
#415770000000
0!
0%
#415775000000
1!
1%
#415780000000
0!
0%
#415785000000
1!
1%
#415790000000
0!
0%
#415795000000
1!
1%
#415800000000
0!
0%
#415805000000
1!
1%
#415810000000
0!
0%
#415815000000
1!
1%
#415820000000
0!
0%
#415825000000
1!
1%
#415830000000
0!
0%
#415835000000
1!
1%
#415840000000
0!
0%
#415845000000
1!
1%
#415850000000
0!
0%
#415855000000
1!
1%
#415860000000
0!
0%
#415865000000
1!
1%
#415870000000
0!
0%
#415875000000
1!
1%
#415880000000
0!
0%
#415885000000
1!
1%
#415890000000
0!
0%
#415895000000
1!
1%
#415900000000
0!
0%
#415905000000
1!
1%
#415910000000
0!
0%
#415915000000
1!
1%
#415920000000
0!
0%
#415925000000
1!
1%
#415930000000
0!
0%
#415935000000
1!
1%
#415940000000
0!
0%
#415945000000
1!
1%
#415950000000
0!
0%
#415955000000
1!
1%
#415960000000
0!
0%
#415965000000
1!
1%
#415970000000
0!
0%
#415975000000
1!
1%
#415980000000
0!
0%
#415985000000
1!
1%
#415990000000
0!
0%
#415995000000
1!
1%
#416000000000
0!
0%
#416005000000
1!
1%
#416010000000
0!
0%
#416015000000
1!
1%
#416020000000
0!
0%
#416025000000
1!
1%
#416030000000
0!
0%
#416035000000
1!
1%
#416040000000
0!
0%
#416045000000
1!
1%
#416050000000
0!
0%
#416055000000
1!
1%
#416060000000
0!
0%
#416065000000
1!
1%
#416070000000
0!
0%
#416075000000
1!
1%
#416080000000
0!
0%
#416085000000
1!
1%
#416090000000
0!
0%
#416095000000
1!
1%
#416100000000
0!
0%
#416105000000
1!
1%
#416110000000
0!
0%
#416115000000
1!
1%
#416120000000
0!
0%
#416125000000
1!
1%
#416130000000
0!
0%
#416135000000
1!
1%
#416140000000
0!
0%
#416145000000
1!
1%
#416150000000
0!
0%
#416155000000
1!
1%
#416160000000
0!
0%
#416165000000
1!
1%
#416170000000
0!
0%
#416175000000
1!
1%
#416180000000
0!
0%
#416185000000
1!
1%
#416190000000
0!
0%
#416195000000
1!
1%
#416200000000
0!
0%
#416205000000
1!
1%
#416210000000
0!
0%
#416215000000
1!
1%
#416220000000
0!
0%
#416225000000
1!
1%
#416230000000
0!
0%
#416235000000
1!
1%
#416240000000
0!
0%
#416245000000
1!
1%
#416250000000
0!
0%
#416255000000
1!
1%
#416260000000
0!
0%
#416265000000
1!
1%
#416270000000
0!
0%
#416275000000
1!
1%
#416280000000
0!
0%
#416285000000
1!
1%
#416290000000
0!
0%
#416295000000
1!
1%
#416300000000
0!
0%
#416305000000
1!
1%
#416310000000
0!
0%
#416315000000
1!
1%
#416320000000
0!
0%
#416325000000
1!
1%
#416330000000
0!
0%
#416335000000
1!
1%
#416340000000
0!
0%
#416345000000
1!
1%
#416350000000
0!
0%
#416355000000
1!
1%
#416360000000
0!
0%
#416365000000
1!
1%
#416370000000
0!
0%
#416375000000
1!
1%
#416380000000
0!
0%
#416385000000
1!
1%
#416390000000
0!
0%
#416395000000
1!
1%
#416400000000
0!
0%
#416405000000
1!
1%
#416410000000
0!
0%
#416415000000
1!
1%
#416420000000
0!
0%
#416425000000
1!
1%
#416430000000
0!
0%
#416435000000
1!
1%
#416440000000
0!
0%
#416445000000
1!
1%
#416450000000
0!
0%
#416455000000
1!
1%
#416460000000
0!
0%
#416465000000
1!
1%
#416470000000
0!
0%
#416475000000
1!
1%
#416480000000
0!
0%
#416485000000
1!
1%
#416490000000
0!
0%
#416495000000
1!
1%
#416500000000
0!
0%
#416505000000
1!
1%
#416510000000
0!
0%
#416515000000
1!
1%
#416520000000
0!
0%
#416525000000
1!
1%
#416530000000
0!
0%
#416535000000
1!
1%
#416540000000
0!
0%
#416545000000
1!
1%
#416550000000
0!
0%
#416555000000
1!
1%
#416560000000
0!
0%
#416565000000
1!
1%
#416570000000
0!
0%
#416575000000
1!
1%
#416580000000
0!
0%
#416585000000
1!
1%
#416590000000
0!
0%
#416595000000
1!
1%
#416600000000
0!
0%
#416605000000
1!
1%
#416610000000
0!
0%
#416615000000
1!
1%
#416620000000
0!
0%
#416625000000
1!
1%
#416630000000
0!
0%
#416635000000
1!
1%
#416640000000
0!
0%
#416645000000
1!
1%
#416650000000
0!
0%
#416655000000
1!
1%
#416660000000
0!
0%
#416665000000
1!
1%
#416670000000
0!
0%
#416675000000
1!
1%
#416680000000
0!
0%
#416685000000
1!
1%
#416690000000
0!
0%
#416695000000
1!
1%
#416700000000
0!
0%
#416705000000
1!
1%
#416710000000
0!
0%
#416715000000
1!
1%
#416720000000
0!
0%
#416725000000
1!
1%
#416730000000
0!
0%
#416735000000
1!
1%
#416740000000
0!
0%
#416745000000
1!
1%
#416750000000
0!
0%
#416755000000
1!
1%
#416760000000
0!
0%
#416765000000
1!
1%
#416770000000
0!
0%
#416775000000
1!
1%
#416780000000
0!
0%
#416785000000
1!
1%
#416790000000
0!
0%
#416795000000
1!
1%
#416800000000
0!
0%
#416805000000
1!
1%
#416810000000
0!
0%
#416815000000
1!
1%
#416820000000
0!
0%
#416825000000
1!
1%
#416830000000
0!
0%
#416835000000
1!
1%
#416840000000
0!
0%
#416845000000
1!
1%
#416850000000
0!
0%
#416855000000
1!
1%
#416860000000
0!
0%
#416865000000
1!
1%
#416870000000
0!
0%
#416875000000
1!
1%
#416880000000
0!
0%
#416885000000
1!
1%
#416890000000
0!
0%
#416895000000
1!
1%
#416900000000
0!
0%
#416905000000
1!
1%
#416910000000
0!
0%
#416915000000
1!
1%
#416920000000
0!
0%
#416925000000
1!
1%
#416930000000
0!
0%
#416935000000
1!
1%
#416940000000
0!
0%
#416945000000
1!
1%
#416950000000
0!
0%
#416955000000
1!
1%
#416960000000
0!
0%
#416965000000
1!
1%
#416970000000
0!
0%
#416975000000
1!
1%
#416980000000
0!
0%
#416985000000
1!
1%
#416990000000
0!
0%
#416995000000
1!
1%
#417000000000
0!
0%
#417005000000
1!
1%
#417010000000
0!
0%
#417015000000
1!
1%
#417020000000
0!
0%
#417025000000
1!
1%
#417030000000
0!
0%
#417035000000
1!
1%
#417040000000
0!
0%
#417045000000
1!
1%
#417050000000
0!
0%
#417055000000
1!
1%
#417060000000
0!
0%
#417065000000
1!
1%
#417070000000
0!
0%
#417075000000
1!
1%
#417080000000
0!
0%
#417085000000
1!
1%
#417090000000
0!
0%
#417095000000
1!
1%
#417100000000
0!
0%
#417105000000
1!
1%
#417110000000
0!
0%
#417115000000
1!
1%
#417120000000
0!
0%
#417125000000
1!
1%
#417130000000
0!
0%
#417135000000
1!
1%
#417140000000
0!
0%
#417145000000
1!
1%
#417150000000
0!
0%
#417155000000
1!
1%
#417160000000
0!
0%
#417165000000
1!
1%
#417170000000
0!
0%
#417175000000
1!
1%
#417180000000
0!
0%
#417185000000
1!
1%
#417190000000
0!
0%
#417195000000
1!
1%
#417200000000
0!
0%
#417205000000
1!
1%
#417210000000
0!
0%
#417215000000
1!
1%
#417220000000
0!
0%
#417225000000
1!
1%
#417230000000
0!
0%
#417235000000
1!
1%
#417240000000
0!
0%
#417245000000
1!
1%
#417250000000
0!
0%
#417255000000
1!
1%
#417260000000
0!
0%
#417265000000
1!
1%
#417270000000
0!
0%
#417275000000
1!
1%
#417280000000
0!
0%
#417285000000
1!
1%
#417290000000
0!
0%
#417295000000
1!
1%
#417300000000
0!
0%
#417305000000
1!
1%
#417310000000
0!
0%
#417315000000
1!
1%
#417320000000
0!
0%
#417325000000
1!
1%
#417330000000
0!
0%
#417335000000
1!
1%
#417340000000
0!
0%
#417345000000
1!
1%
#417350000000
0!
0%
#417355000000
1!
1%
#417360000000
0!
0%
#417365000000
1!
1%
#417370000000
0!
0%
#417375000000
1!
1%
#417380000000
0!
0%
#417385000000
1!
1%
#417390000000
0!
0%
#417395000000
1!
1%
#417400000000
0!
0%
#417405000000
1!
1%
#417410000000
0!
0%
#417415000000
1!
1%
#417420000000
0!
0%
#417425000000
1!
1%
#417430000000
0!
0%
#417435000000
1!
1%
#417440000000
0!
0%
#417445000000
1!
1%
#417450000000
0!
0%
#417455000000
1!
1%
#417460000000
0!
0%
#417465000000
1!
1%
#417470000000
0!
0%
#417475000000
1!
1%
#417480000000
0!
0%
#417485000000
1!
1%
#417490000000
0!
0%
#417495000000
1!
1%
#417500000000
0!
0%
#417505000000
1!
1%
#417510000000
0!
0%
#417515000000
1!
1%
#417520000000
0!
0%
#417525000000
1!
1%
#417530000000
0!
0%
#417535000000
1!
1%
#417540000000
0!
0%
#417545000000
1!
1%
#417550000000
0!
0%
#417555000000
1!
1%
#417560000000
0!
0%
#417565000000
1!
1%
#417570000000
0!
0%
#417575000000
1!
1%
#417580000000
0!
0%
#417585000000
1!
1%
#417590000000
0!
0%
#417595000000
1!
1%
#417600000000
0!
0%
#417605000000
1!
1%
#417610000000
0!
0%
#417615000000
1!
1%
#417620000000
0!
0%
#417625000000
1!
1%
#417630000000
0!
0%
#417635000000
1!
1%
#417640000000
0!
0%
#417645000000
1!
1%
#417650000000
0!
0%
#417655000000
1!
1%
#417660000000
0!
0%
#417665000000
1!
1%
#417670000000
0!
0%
#417675000000
1!
1%
#417680000000
0!
0%
#417685000000
1!
1%
#417690000000
0!
0%
#417695000000
1!
1%
#417700000000
0!
0%
#417705000000
1!
1%
#417710000000
0!
0%
#417715000000
1!
1%
#417720000000
0!
0%
#417725000000
1!
1%
#417730000000
0!
0%
#417735000000
1!
1%
#417740000000
0!
0%
#417745000000
1!
1%
#417750000000
0!
0%
#417755000000
1!
1%
#417760000000
0!
0%
#417765000000
1!
1%
#417770000000
0!
0%
#417775000000
1!
1%
#417780000000
0!
0%
#417785000000
1!
1%
#417790000000
0!
0%
#417795000000
1!
1%
#417800000000
0!
0%
#417805000000
1!
1%
#417810000000
0!
0%
#417815000000
1!
1%
#417820000000
0!
0%
#417825000000
1!
1%
#417830000000
0!
0%
#417835000000
1!
1%
#417840000000
0!
0%
#417845000000
1!
1%
#417850000000
0!
0%
#417855000000
1!
1%
#417860000000
0!
0%
#417865000000
1!
1%
#417870000000
0!
0%
#417875000000
1!
1%
#417880000000
0!
0%
#417885000000
1!
1%
#417890000000
0!
0%
#417895000000
1!
1%
#417900000000
0!
0%
#417905000000
1!
1%
#417910000000
0!
0%
#417915000000
1!
1%
#417920000000
0!
0%
#417925000000
1!
1%
#417930000000
0!
0%
#417935000000
1!
1%
#417940000000
0!
0%
#417945000000
1!
1%
#417950000000
0!
0%
#417955000000
1!
1%
#417960000000
0!
0%
#417965000000
1!
1%
#417970000000
0!
0%
#417975000000
1!
1%
#417980000000
0!
0%
#417985000000
1!
1%
#417990000000
0!
0%
#417995000000
1!
1%
#418000000000
0!
0%
#418005000000
1!
1%
#418010000000
0!
0%
#418015000000
1!
1%
#418020000000
0!
0%
#418025000000
1!
1%
#418030000000
0!
0%
#418035000000
1!
1%
#418040000000
0!
0%
#418045000000
1!
1%
#418050000000
0!
0%
#418055000000
1!
1%
#418060000000
0!
0%
#418065000000
1!
1%
#418070000000
0!
0%
#418075000000
1!
1%
#418080000000
0!
0%
#418085000000
1!
1%
#418090000000
0!
0%
#418095000000
1!
1%
#418100000000
0!
0%
#418105000000
1!
1%
#418110000000
0!
0%
#418115000000
1!
1%
#418120000000
0!
0%
#418125000000
1!
1%
#418130000000
0!
0%
#418135000000
1!
1%
#418140000000
0!
0%
#418145000000
1!
1%
#418150000000
0!
0%
#418155000000
1!
1%
#418160000000
0!
0%
#418165000000
1!
1%
#418170000000
0!
0%
#418175000000
1!
1%
#418180000000
0!
0%
#418185000000
1!
1%
#418190000000
0!
0%
#418195000000
1!
1%
#418200000000
0!
0%
#418205000000
1!
1%
#418210000000
0!
0%
#418215000000
1!
1%
#418220000000
0!
0%
#418225000000
1!
1%
#418230000000
0!
0%
#418235000000
1!
1%
#418240000000
0!
0%
#418245000000
1!
1%
#418250000000
0!
0%
#418255000000
1!
1%
#418260000000
0!
0%
#418265000000
1!
1%
#418270000000
0!
0%
#418275000000
1!
1%
#418280000000
0!
0%
#418285000000
1!
1%
#418290000000
0!
0%
#418295000000
1!
1%
#418300000000
0!
0%
#418305000000
1!
1%
#418310000000
0!
0%
#418315000000
1!
1%
#418320000000
0!
0%
#418325000000
1!
1%
#418330000000
0!
0%
#418335000000
1!
1%
#418340000000
0!
0%
#418345000000
1!
1%
#418350000000
0!
0%
#418355000000
1!
1%
#418360000000
0!
0%
#418365000000
1!
1%
#418370000000
0!
0%
#418375000000
1!
1%
#418380000000
0!
0%
#418385000000
1!
1%
#418390000000
0!
0%
#418395000000
1!
1%
#418400000000
0!
0%
#418405000000
1!
1%
#418410000000
0!
0%
#418415000000
1!
1%
#418420000000
0!
0%
#418425000000
1!
1%
#418430000000
0!
0%
#418435000000
1!
1%
#418440000000
0!
0%
#418445000000
1!
1%
#418450000000
0!
0%
#418455000000
1!
1%
#418460000000
0!
0%
#418465000000
1!
1%
#418470000000
0!
0%
#418475000000
1!
1%
#418480000000
0!
0%
#418485000000
1!
1%
#418490000000
0!
0%
#418495000000
1!
1%
#418500000000
0!
0%
#418505000000
1!
1%
#418510000000
0!
0%
#418515000000
1!
1%
#418520000000
0!
0%
#418525000000
1!
1%
#418530000000
0!
0%
#418535000000
1!
1%
#418540000000
0!
0%
#418545000000
1!
1%
#418550000000
0!
0%
#418555000000
1!
1%
#418560000000
0!
0%
#418565000000
1!
1%
#418570000000
0!
0%
#418575000000
1!
1%
#418580000000
0!
0%
#418585000000
1!
1%
#418590000000
0!
0%
#418595000000
1!
1%
#418600000000
0!
0%
#418605000000
1!
1%
#418610000000
0!
0%
#418615000000
1!
1%
#418620000000
0!
0%
#418625000000
1!
1%
#418630000000
0!
0%
#418635000000
1!
1%
#418640000000
0!
0%
#418645000000
1!
1%
#418650000000
0!
0%
#418655000000
1!
1%
#418660000000
0!
0%
#418665000000
1!
1%
#418670000000
0!
0%
#418675000000
1!
1%
#418680000000
0!
0%
#418685000000
1!
1%
#418690000000
0!
0%
#418695000000
1!
1%
#418700000000
0!
0%
#418705000000
1!
1%
#418710000000
0!
0%
#418715000000
1!
1%
#418720000000
0!
0%
#418725000000
1!
1%
#418730000000
0!
0%
#418735000000
1!
1%
#418740000000
0!
0%
#418745000000
1!
1%
#418750000000
0!
0%
#418755000000
1!
1%
#418760000000
0!
0%
#418765000000
1!
1%
#418770000000
0!
0%
#418775000000
1!
1%
#418780000000
0!
0%
#418785000000
1!
1%
#418790000000
0!
0%
#418795000000
1!
1%
#418800000000
0!
0%
#418805000000
1!
1%
#418810000000
0!
0%
#418815000000
1!
1%
#418820000000
0!
0%
#418825000000
1!
1%
#418830000000
0!
0%
#418835000000
1!
1%
#418840000000
0!
0%
#418845000000
1!
1%
#418850000000
0!
0%
#418855000000
1!
1%
#418860000000
0!
0%
#418865000000
1!
1%
#418870000000
0!
0%
#418875000000
1!
1%
#418880000000
0!
0%
#418885000000
1!
1%
#418890000000
0!
0%
#418895000000
1!
1%
#418900000000
0!
0%
#418905000000
1!
1%
#418910000000
0!
0%
#418915000000
1!
1%
#418920000000
0!
0%
#418925000000
1!
1%
#418930000000
0!
0%
#418935000000
1!
1%
#418940000000
0!
0%
#418945000000
1!
1%
#418950000000
0!
0%
#418955000000
1!
1%
#418960000000
0!
0%
#418965000000
1!
1%
#418970000000
0!
0%
#418975000000
1!
1%
#418980000000
0!
0%
#418985000000
1!
1%
#418990000000
0!
0%
#418995000000
1!
1%
#419000000000
0!
0%
#419005000000
1!
1%
#419010000000
0!
0%
#419015000000
1!
1%
#419020000000
0!
0%
#419025000000
1!
1%
#419030000000
0!
0%
#419035000000
1!
1%
#419040000000
0!
0%
#419045000000
1!
1%
#419050000000
0!
0%
#419055000000
1!
1%
#419060000000
0!
0%
#419065000000
1!
1%
#419070000000
0!
0%
#419075000000
1!
1%
#419080000000
0!
0%
#419085000000
1!
1%
#419090000000
0!
0%
#419095000000
1!
1%
#419100000000
0!
0%
#419105000000
1!
1%
#419110000000
0!
0%
#419115000000
1!
1%
#419120000000
0!
0%
#419125000000
1!
1%
#419130000000
0!
0%
#419135000000
1!
1%
#419140000000
0!
0%
#419145000000
1!
1%
#419150000000
0!
0%
#419155000000
1!
1%
#419160000000
0!
0%
#419165000000
1!
1%
#419170000000
0!
0%
#419175000000
1!
1%
#419180000000
0!
0%
#419185000000
1!
1%
#419190000000
0!
0%
#419195000000
1!
1%
#419200000000
0!
0%
#419205000000
1!
1%
#419210000000
0!
0%
#419215000000
1!
1%
#419220000000
0!
0%
#419225000000
1!
1%
#419230000000
0!
0%
#419235000000
1!
1%
#419240000000
0!
0%
#419245000000
1!
1%
#419250000000
0!
0%
#419255000000
1!
1%
#419260000000
0!
0%
#419265000000
1!
1%
#419270000000
0!
0%
#419275000000
1!
1%
#419280000000
0!
0%
#419285000000
1!
1%
#419290000000
0!
0%
#419295000000
1!
1%
#419300000000
0!
0%
#419305000000
1!
1%
#419310000000
0!
0%
#419315000000
1!
1%
#419320000000
0!
0%
#419325000000
1!
1%
#419330000000
0!
0%
#419335000000
1!
1%
#419340000000
0!
0%
#419345000000
1!
1%
#419350000000
0!
0%
#419355000000
1!
1%
#419360000000
0!
0%
#419365000000
1!
1%
#419370000000
0!
0%
#419375000000
1!
1%
#419380000000
0!
0%
#419385000000
1!
1%
#419390000000
0!
0%
#419395000000
1!
1%
#419400000000
0!
0%
#419405000000
1!
1%
#419410000000
0!
0%
#419415000000
1!
1%
#419420000000
0!
0%
#419425000000
1!
1%
#419430000000
0!
0%
#419435000000
1!
1%
#419440000000
0!
0%
#419445000000
1!
1%
#419450000000
0!
0%
#419455000000
1!
1%
#419460000000
0!
0%
#419465000000
1!
1%
#419470000000
0!
0%
#419475000000
1!
1%
#419480000000
0!
0%
#419485000000
1!
1%
#419490000000
0!
0%
#419495000000
1!
1%
#419500000000
0!
0%
#419505000000
1!
1%
#419510000000
0!
0%
#419515000000
1!
1%
#419520000000
0!
0%
#419525000000
1!
1%
#419530000000
0!
0%
#419535000000
1!
1%
#419540000000
0!
0%
#419545000000
1!
1%
#419550000000
0!
0%
#419555000000
1!
1%
#419560000000
0!
0%
#419565000000
1!
1%
#419570000000
0!
0%
#419575000000
1!
1%
#419580000000
0!
0%
#419585000000
1!
1%
#419590000000
0!
0%
#419595000000
1!
1%
#419600000000
0!
0%
#419605000000
1!
1%
#419610000000
0!
0%
#419615000000
1!
1%
#419620000000
0!
0%
#419625000000
1!
1%
#419630000000
0!
0%
#419635000000
1!
1%
#419640000000
0!
0%
#419645000000
1!
1%
#419650000000
0!
0%
#419655000000
1!
1%
#419660000000
0!
0%
#419665000000
1!
1%
#419670000000
0!
0%
#419675000000
1!
1%
#419680000000
0!
0%
#419685000000
1!
1%
#419690000000
0!
0%
#419695000000
1!
1%
#419700000000
0!
0%
#419705000000
1!
1%
#419710000000
0!
0%
#419715000000
1!
1%
#419720000000
0!
0%
#419725000000
1!
1%
#419730000000
0!
0%
#419735000000
1!
1%
#419740000000
0!
0%
#419745000000
1!
1%
#419750000000
0!
0%
#419755000000
1!
1%
#419760000000
0!
0%
#419765000000
1!
1%
#419770000000
0!
0%
#419775000000
1!
1%
#419780000000
0!
0%
#419785000000
1!
1%
#419790000000
0!
0%
#419795000000
1!
1%
#419800000000
0!
0%
#419805000000
1!
1%
#419810000000
0!
0%
#419815000000
1!
1%
#419820000000
0!
0%
#419825000000
1!
1%
#419830000000
0!
0%
#419835000000
1!
1%
#419840000000
0!
0%
#419845000000
1!
1%
#419850000000
0!
0%
#419855000000
1!
1%
#419860000000
0!
0%
#419865000000
1!
1%
#419870000000
0!
0%
#419875000000
1!
1%
#419880000000
0!
0%
#419885000000
1!
1%
#419890000000
0!
0%
#419895000000
1!
1%
#419900000000
0!
0%
#419905000000
1!
1%
#419910000000
0!
0%
#419915000000
1!
1%
#419920000000
0!
0%
#419925000000
1!
1%
#419930000000
0!
0%
#419935000000
1!
1%
#419940000000
0!
0%
#419945000000
1!
1%
#419950000000
0!
0%
#419955000000
1!
1%
#419960000000
0!
0%
#419965000000
1!
1%
#419970000000
0!
0%
#419975000000
1!
1%
#419980000000
0!
0%
#419985000000
1!
1%
#419990000000
0!
0%
#419995000000
1!
1%
#420000000000
0!
0%
#420005000000
1!
1%
#420010000000
0!
0%
#420015000000
1!
1%
#420020000000
0!
0%
#420025000000
1!
1%
#420030000000
0!
0%
#420035000000
1!
1%
#420040000000
0!
0%
#420045000000
1!
1%
#420050000000
0!
0%
#420055000000
1!
1%
#420060000000
0!
0%
#420065000000
1!
1%
#420070000000
0!
0%
#420075000000
1!
1%
#420080000000
0!
0%
#420085000000
1!
1%
#420090000000
0!
0%
#420095000000
1!
1%
#420100000000
0!
0%
#420105000000
1!
1%
#420110000000
0!
0%
#420115000000
1!
1%
#420120000000
0!
0%
#420125000000
1!
1%
#420130000000
0!
0%
#420135000000
1!
1%
#420140000000
0!
0%
#420145000000
1!
1%
#420150000000
0!
0%
#420155000000
1!
1%
#420160000000
0!
0%
#420165000000
1!
1%
#420170000000
0!
0%
#420175000000
1!
1%
#420180000000
0!
0%
#420185000000
1!
1%
#420190000000
0!
0%
#420195000000
1!
1%
#420200000000
0!
0%
#420205000000
1!
1%
#420210000000
0!
0%
#420215000000
1!
1%
#420220000000
0!
0%
#420225000000
1!
1%
#420230000000
0!
0%
#420235000000
1!
1%
#420240000000
0!
0%
#420245000000
1!
1%
#420250000000
0!
0%
#420255000000
1!
1%
#420260000000
0!
0%
#420265000000
1!
1%
#420270000000
0!
0%
#420275000000
1!
1%
#420280000000
0!
0%
#420285000000
1!
1%
#420290000000
0!
0%
#420295000000
1!
1%
#420300000000
0!
0%
#420305000000
1!
1%
#420310000000
0!
0%
#420315000000
1!
1%
#420320000000
0!
0%
#420325000000
1!
1%
#420330000000
0!
0%
#420335000000
1!
1%
#420340000000
0!
0%
#420345000000
1!
1%
#420350000000
0!
0%
#420355000000
1!
1%
#420360000000
0!
0%
#420365000000
1!
1%
#420370000000
0!
0%
#420375000000
1!
1%
#420380000000
0!
0%
#420385000000
1!
1%
#420390000000
0!
0%
#420395000000
1!
1%
#420400000000
0!
0%
#420405000000
1!
1%
#420410000000
0!
0%
#420415000000
1!
1%
#420420000000
0!
0%
#420425000000
1!
1%
#420430000000
0!
0%
#420435000000
1!
1%
#420440000000
0!
0%
#420445000000
1!
1%
#420450000000
0!
0%
#420455000000
1!
1%
#420460000000
0!
0%
#420465000000
1!
1%
#420470000000
0!
0%
#420475000000
1!
1%
#420480000000
0!
0%
#420485000000
1!
1%
#420490000000
0!
0%
#420495000000
1!
1%
#420500000000
0!
0%
#420505000000
1!
1%
#420510000000
0!
0%
#420515000000
1!
1%
#420520000000
0!
0%
#420525000000
1!
1%
#420530000000
0!
0%
#420535000000
1!
1%
#420540000000
0!
0%
#420545000000
1!
1%
#420550000000
0!
0%
#420555000000
1!
1%
#420560000000
0!
0%
#420565000000
1!
1%
#420570000000
0!
0%
#420575000000
1!
1%
#420580000000
0!
0%
#420585000000
1!
1%
#420590000000
0!
0%
#420595000000
1!
1%
#420600000000
0!
0%
#420605000000
1!
1%
#420610000000
0!
0%
#420615000000
1!
1%
#420620000000
0!
0%
#420625000000
1!
1%
#420630000000
0!
0%
#420635000000
1!
1%
#420640000000
0!
0%
#420645000000
1!
1%
#420650000000
0!
0%
#420655000000
1!
1%
#420660000000
0!
0%
#420665000000
1!
1%
#420670000000
0!
0%
#420675000000
1!
1%
#420680000000
0!
0%
#420685000000
1!
1%
#420690000000
0!
0%
#420695000000
1!
1%
#420700000000
0!
0%
#420705000000
1!
1%
#420710000000
0!
0%
#420715000000
1!
1%
#420720000000
0!
0%
#420725000000
1!
1%
#420730000000
0!
0%
#420735000000
1!
1%
#420740000000
0!
0%
#420745000000
1!
1%
#420750000000
0!
0%
#420755000000
1!
1%
#420760000000
0!
0%
#420765000000
1!
1%
#420770000000
0!
0%
#420775000000
1!
1%
#420780000000
0!
0%
#420785000000
1!
1%
#420790000000
0!
0%
#420795000000
1!
1%
#420800000000
0!
0%
#420805000000
1!
1%
#420810000000
0!
0%
#420815000000
1!
1%
#420820000000
0!
0%
#420825000000
1!
1%
#420830000000
0!
0%
#420835000000
1!
1%
#420840000000
0!
0%
#420845000000
1!
1%
#420850000000
0!
0%
#420855000000
1!
1%
#420860000000
0!
0%
#420865000000
1!
1%
#420870000000
0!
0%
#420875000000
1!
1%
#420880000000
0!
0%
#420885000000
1!
1%
#420890000000
0!
0%
#420895000000
1!
1%
#420900000000
0!
0%
#420905000000
1!
1%
#420910000000
0!
0%
#420915000000
1!
1%
#420920000000
0!
0%
#420925000000
1!
1%
#420930000000
0!
0%
#420935000000
1!
1%
#420940000000
0!
0%
#420945000000
1!
1%
#420950000000
0!
0%
#420955000000
1!
1%
#420960000000
0!
0%
#420965000000
1!
1%
#420970000000
0!
0%
#420975000000
1!
1%
#420980000000
0!
0%
#420985000000
1!
1%
#420990000000
0!
0%
#420995000000
1!
1%
#421000000000
0!
0%
#421005000000
1!
1%
#421010000000
0!
0%
#421015000000
1!
1%
#421020000000
0!
0%
#421025000000
1!
1%
#421030000000
0!
0%
#421035000000
1!
1%
#421040000000
0!
0%
#421045000000
1!
1%
#421050000000
0!
0%
#421055000000
1!
1%
#421060000000
0!
0%
#421065000000
1!
1%
#421070000000
0!
0%
#421075000000
1!
1%
#421080000000
0!
0%
#421085000000
1!
1%
#421090000000
0!
0%
#421095000000
1!
1%
#421100000000
0!
0%
#421105000000
1!
1%
#421110000000
0!
0%
#421115000000
1!
1%
#421120000000
0!
0%
#421125000000
1!
1%
#421130000000
0!
0%
#421135000000
1!
1%
#421140000000
0!
0%
#421145000000
1!
1%
#421150000000
0!
0%
#421155000000
1!
1%
#421160000000
0!
0%
#421165000000
1!
1%
#421170000000
0!
0%
#421175000000
1!
1%
#421180000000
0!
0%
#421185000000
1!
1%
#421190000000
0!
0%
#421195000000
1!
1%
#421200000000
0!
0%
#421205000000
1!
1%
#421210000000
0!
0%
#421215000000
1!
1%
#421220000000
0!
0%
#421225000000
1!
1%
#421230000000
0!
0%
#421235000000
1!
1%
#421240000000
0!
0%
#421245000000
1!
1%
#421250000000
0!
0%
#421255000000
1!
1%
#421260000000
0!
0%
#421265000000
1!
1%
#421270000000
0!
0%
#421275000000
1!
1%
#421280000000
0!
0%
#421285000000
1!
1%
#421290000000
0!
0%
#421295000000
1!
1%
#421300000000
0!
0%
#421305000000
1!
1%
#421310000000
0!
0%
#421315000000
1!
1%
#421320000000
0!
0%
#421325000000
1!
1%
#421330000000
0!
0%
#421335000000
1!
1%
#421340000000
0!
0%
#421345000000
1!
1%
#421350000000
0!
0%
#421355000000
1!
1%
#421360000000
0!
0%
#421365000000
1!
1%
#421370000000
0!
0%
#421375000000
1!
1%
#421380000000
0!
0%
#421385000000
1!
1%
#421390000000
0!
0%
#421395000000
1!
1%
#421400000000
0!
0%
#421405000000
1!
1%
#421410000000
0!
0%
#421415000000
1!
1%
#421420000000
0!
0%
#421425000000
1!
1%
#421430000000
0!
0%
#421435000000
1!
1%
#421440000000
0!
0%
#421445000000
1!
1%
#421450000000
0!
0%
#421455000000
1!
1%
#421460000000
0!
0%
#421465000000
1!
1%
#421470000000
0!
0%
#421475000000
1!
1%
#421480000000
0!
0%
#421485000000
1!
1%
#421490000000
0!
0%
#421495000000
1!
1%
#421500000000
0!
0%
#421505000000
1!
1%
#421510000000
0!
0%
#421515000000
1!
1%
#421520000000
0!
0%
#421525000000
1!
1%
#421530000000
0!
0%
#421535000000
1!
1%
#421540000000
0!
0%
#421545000000
1!
1%
#421550000000
0!
0%
#421555000000
1!
1%
#421560000000
0!
0%
#421565000000
1!
1%
#421570000000
0!
0%
#421575000000
1!
1%
#421580000000
0!
0%
#421585000000
1!
1%
#421590000000
0!
0%
#421595000000
1!
1%
#421600000000
0!
0%
#421605000000
1!
1%
#421610000000
0!
0%
#421615000000
1!
1%
#421620000000
0!
0%
#421625000000
1!
1%
#421630000000
0!
0%
#421635000000
1!
1%
#421640000000
0!
0%
#421645000000
1!
1%
#421650000000
0!
0%
#421655000000
1!
1%
#421660000000
0!
0%
#421665000000
1!
1%
#421670000000
0!
0%
#421675000000
1!
1%
#421680000000
0!
0%
#421685000000
1!
1%
#421690000000
0!
0%
#421695000000
1!
1%
#421700000000
0!
0%
#421705000000
1!
1%
#421710000000
0!
0%
#421715000000
1!
1%
#421720000000
0!
0%
#421725000000
1!
1%
#421730000000
0!
0%
#421735000000
1!
1%
#421740000000
0!
0%
#421745000000
1!
1%
#421750000000
0!
0%
#421755000000
1!
1%
#421760000000
0!
0%
#421765000000
1!
1%
#421770000000
0!
0%
#421775000000
1!
1%
#421780000000
0!
0%
#421785000000
1!
1%
#421790000000
0!
0%
#421795000000
1!
1%
#421800000000
0!
0%
#421805000000
1!
1%
#421810000000
0!
0%
#421815000000
1!
1%
#421820000000
0!
0%
#421825000000
1!
1%
#421830000000
0!
0%
#421835000000
1!
1%
#421840000000
0!
0%
#421845000000
1!
1%
#421850000000
0!
0%
#421855000000
1!
1%
#421860000000
0!
0%
#421865000000
1!
1%
#421870000000
0!
0%
#421875000000
1!
1%
#421880000000
0!
0%
#421885000000
1!
1%
#421890000000
0!
0%
#421895000000
1!
1%
#421900000000
0!
0%
#421905000000
1!
1%
#421910000000
0!
0%
#421915000000
1!
1%
#421920000000
0!
0%
#421925000000
1!
1%
#421930000000
0!
0%
#421935000000
1!
1%
#421940000000
0!
0%
#421945000000
1!
1%
#421950000000
0!
0%
#421955000000
1!
1%
#421960000000
0!
0%
#421965000000
1!
1%
#421970000000
0!
0%
#421975000000
1!
1%
#421980000000
0!
0%
#421985000000
1!
1%
#421990000000
0!
0%
#421995000000
1!
1%
#422000000000
0!
0%
#422005000000
1!
1%
#422010000000
0!
0%
#422015000000
1!
1%
#422020000000
0!
0%
#422025000000
1!
1%
#422030000000
0!
0%
#422035000000
1!
1%
#422040000000
0!
0%
#422045000000
1!
1%
#422050000000
0!
0%
#422055000000
1!
1%
#422060000000
0!
0%
#422065000000
1!
1%
#422070000000
0!
0%
#422075000000
1!
1%
#422080000000
0!
0%
#422085000000
1!
1%
#422090000000
0!
0%
#422095000000
1!
1%
#422100000000
0!
0%
#422105000000
1!
1%
#422110000000
0!
0%
#422115000000
1!
1%
#422120000000
0!
0%
#422125000000
1!
1%
#422130000000
0!
0%
#422135000000
1!
1%
#422140000000
0!
0%
#422145000000
1!
1%
#422150000000
0!
0%
#422155000000
1!
1%
#422160000000
0!
0%
#422165000000
1!
1%
#422170000000
0!
0%
#422175000000
1!
1%
#422180000000
0!
0%
#422185000000
1!
1%
#422190000000
0!
0%
#422195000000
1!
1%
#422200000000
0!
0%
#422205000000
1!
1%
#422210000000
0!
0%
#422215000000
1!
1%
#422220000000
0!
0%
#422225000000
1!
1%
#422230000000
0!
0%
#422235000000
1!
1%
#422240000000
0!
0%
#422245000000
1!
1%
#422250000000
0!
0%
#422255000000
1!
1%
#422260000000
0!
0%
#422265000000
1!
1%
#422270000000
0!
0%
#422275000000
1!
1%
#422280000000
0!
0%
#422285000000
1!
1%
#422290000000
0!
0%
#422295000000
1!
1%
#422300000000
0!
0%
#422305000000
1!
1%
#422310000000
0!
0%
#422315000000
1!
1%
#422320000000
0!
0%
#422325000000
1!
1%
#422330000000
0!
0%
#422335000000
1!
1%
#422340000000
0!
0%
#422345000000
1!
1%
#422350000000
0!
0%
#422355000000
1!
1%
#422360000000
0!
0%
#422365000000
1!
1%
#422370000000
0!
0%
#422375000000
1!
1%
#422380000000
0!
0%
#422385000000
1!
1%
#422390000000
0!
0%
#422395000000
1!
1%
#422400000000
0!
0%
#422405000000
1!
1%
#422410000000
0!
0%
#422415000000
1!
1%
#422420000000
0!
0%
#422425000000
1!
1%
#422430000000
0!
0%
#422435000000
1!
1%
#422440000000
0!
0%
#422445000000
1!
1%
#422450000000
0!
0%
#422455000000
1!
1%
#422460000000
0!
0%
#422465000000
1!
1%
#422470000000
0!
0%
#422475000000
1!
1%
#422480000000
0!
0%
#422485000000
1!
1%
#422490000000
0!
0%
#422495000000
1!
1%
#422500000000
0!
0%
#422505000000
1!
1%
#422510000000
0!
0%
#422515000000
1!
1%
#422520000000
0!
0%
#422525000000
1!
1%
#422530000000
0!
0%
#422535000000
1!
1%
#422540000000
0!
0%
#422545000000
1!
1%
#422550000000
0!
0%
#422555000000
1!
1%
#422560000000
0!
0%
#422565000000
1!
1%
#422570000000
0!
0%
#422575000000
1!
1%
#422580000000
0!
0%
#422585000000
1!
1%
#422590000000
0!
0%
#422595000000
1!
1%
#422600000000
0!
0%
#422605000000
1!
1%
#422610000000
0!
0%
#422615000000
1!
1%
#422620000000
0!
0%
#422625000000
1!
1%
#422630000000
0!
0%
#422635000000
1!
1%
#422640000000
0!
0%
#422645000000
1!
1%
#422650000000
0!
0%
#422655000000
1!
1%
#422660000000
0!
0%
#422665000000
1!
1%
#422670000000
0!
0%
#422675000000
1!
1%
#422680000000
0!
0%
#422685000000
1!
1%
#422690000000
0!
0%
#422695000000
1!
1%
#422700000000
0!
0%
#422705000000
1!
1%
#422710000000
0!
0%
#422715000000
1!
1%
#422720000000
0!
0%
#422725000000
1!
1%
#422730000000
0!
0%
#422735000000
1!
1%
#422740000000
0!
0%
#422745000000
1!
1%
#422750000000
0!
0%
#422755000000
1!
1%
#422760000000
0!
0%
#422765000000
1!
1%
#422770000000
0!
0%
#422775000000
1!
1%
#422780000000
0!
0%
#422785000000
1!
1%
#422790000000
0!
0%
#422795000000
1!
1%
#422800000000
0!
0%
#422805000000
1!
1%
#422810000000
0!
0%
#422815000000
1!
1%
#422820000000
0!
0%
#422825000000
1!
1%
#422830000000
0!
0%
#422835000000
1!
1%
#422840000000
0!
0%
#422845000000
1!
1%
#422850000000
0!
0%
#422855000000
1!
1%
#422860000000
0!
0%
#422865000000
1!
1%
#422870000000
0!
0%
#422875000000
1!
1%
#422880000000
0!
0%
#422885000000
1!
1%
#422890000000
0!
0%
#422895000000
1!
1%
#422900000000
0!
0%
#422905000000
1!
1%
#422910000000
0!
0%
#422915000000
1!
1%
#422920000000
0!
0%
#422925000000
1!
1%
#422930000000
0!
0%
#422935000000
1!
1%
#422940000000
0!
0%
#422945000000
1!
1%
#422950000000
0!
0%
#422955000000
1!
1%
#422960000000
0!
0%
#422965000000
1!
1%
#422970000000
0!
0%
#422975000000
1!
1%
#422980000000
0!
0%
#422985000000
1!
1%
#422990000000
0!
0%
#422995000000
1!
1%
#423000000000
0!
0%
#423005000000
1!
1%
#423010000000
0!
0%
#423015000000
1!
1%
#423020000000
0!
0%
#423025000000
1!
1%
#423030000000
0!
0%
#423035000000
1!
1%
#423040000000
0!
0%
#423045000000
1!
1%
#423050000000
0!
0%
#423055000000
1!
1%
#423060000000
0!
0%
#423065000000
1!
1%
#423070000000
0!
0%
#423075000000
1!
1%
#423080000000
0!
0%
#423085000000
1!
1%
#423090000000
0!
0%
#423095000000
1!
1%
#423100000000
0!
0%
#423105000000
1!
1%
#423110000000
0!
0%
#423115000000
1!
1%
#423120000000
0!
0%
#423125000000
1!
1%
#423130000000
0!
0%
#423135000000
1!
1%
#423140000000
0!
0%
#423145000000
1!
1%
#423150000000
0!
0%
#423155000000
1!
1%
#423160000000
0!
0%
#423165000000
1!
1%
#423170000000
0!
0%
#423175000000
1!
1%
#423180000000
0!
0%
#423185000000
1!
1%
#423190000000
0!
0%
#423195000000
1!
1%
#423200000000
0!
0%
#423205000000
1!
1%
#423210000000
0!
0%
#423215000000
1!
1%
#423220000000
0!
0%
#423225000000
1!
1%
#423230000000
0!
0%
#423235000000
1!
1%
#423240000000
0!
0%
#423245000000
1!
1%
#423250000000
0!
0%
#423255000000
1!
1%
#423260000000
0!
0%
#423265000000
1!
1%
#423270000000
0!
0%
#423275000000
1!
1%
#423280000000
0!
0%
#423285000000
1!
1%
#423290000000
0!
0%
#423295000000
1!
1%
#423300000000
0!
0%
#423305000000
1!
1%
#423310000000
0!
0%
#423315000000
1!
1%
#423320000000
0!
0%
#423325000000
1!
1%
#423330000000
0!
0%
#423335000000
1!
1%
#423340000000
0!
0%
#423345000000
1!
1%
#423350000000
0!
0%
#423355000000
1!
1%
#423360000000
0!
0%
#423365000000
1!
1%
#423370000000
0!
0%
#423375000000
1!
1%
#423380000000
0!
0%
#423385000000
1!
1%
#423390000000
0!
0%
#423395000000
1!
1%
#423400000000
0!
0%
#423405000000
1!
1%
#423410000000
0!
0%
#423415000000
1!
1%
#423420000000
0!
0%
#423425000000
1!
1%
#423430000000
0!
0%
#423435000000
1!
1%
#423440000000
0!
0%
#423445000000
1!
1%
#423450000000
0!
0%
#423455000000
1!
1%
#423460000000
0!
0%
#423465000000
1!
1%
#423470000000
0!
0%
#423475000000
1!
1%
#423480000000
0!
0%
#423485000000
1!
1%
#423490000000
0!
0%
#423495000000
1!
1%
#423500000000
0!
0%
#423505000000
1!
1%
#423510000000
0!
0%
#423515000000
1!
1%
#423520000000
0!
0%
#423525000000
1!
1%
#423530000000
0!
0%
#423535000000
1!
1%
#423540000000
0!
0%
#423545000000
1!
1%
#423550000000
0!
0%
#423555000000
1!
1%
#423560000000
0!
0%
#423565000000
1!
1%
#423570000000
0!
0%
#423575000000
1!
1%
#423580000000
0!
0%
#423585000000
1!
1%
#423590000000
0!
0%
#423595000000
1!
1%
#423600000000
0!
0%
#423605000000
1!
1%
#423610000000
0!
0%
#423615000000
1!
1%
#423620000000
0!
0%
#423625000000
1!
1%
#423630000000
0!
0%
#423635000000
1!
1%
#423640000000
0!
0%
#423645000000
1!
1%
#423650000000
0!
0%
#423655000000
1!
1%
#423660000000
0!
0%
#423665000000
1!
1%
#423670000000
0!
0%
#423675000000
1!
1%
#423680000000
0!
0%
#423685000000
1!
1%
#423690000000
0!
0%
#423695000000
1!
1%
#423700000000
0!
0%
#423705000000
1!
1%
#423710000000
0!
0%
#423715000000
1!
1%
#423720000000
0!
0%
#423725000000
1!
1%
#423730000000
0!
0%
#423735000000
1!
1%
#423740000000
0!
0%
#423745000000
1!
1%
#423750000000
0!
0%
#423755000000
1!
1%
#423760000000
0!
0%
#423765000000
1!
1%
#423770000000
0!
0%
#423775000000
1!
1%
#423780000000
0!
0%
#423785000000
1!
1%
#423790000000
0!
0%
#423795000000
1!
1%
#423800000000
0!
0%
#423805000000
1!
1%
#423810000000
0!
0%
#423815000000
1!
1%
#423820000000
0!
0%
#423825000000
1!
1%
#423830000000
0!
0%
#423835000000
1!
1%
#423840000000
0!
0%
#423845000000
1!
1%
#423850000000
0!
0%
#423855000000
1!
1%
#423860000000
0!
0%
#423865000000
1!
1%
#423870000000
0!
0%
#423875000000
1!
1%
#423880000000
0!
0%
#423885000000
1!
1%
#423890000000
0!
0%
#423895000000
1!
1%
#423900000000
0!
0%
#423905000000
1!
1%
#423910000000
0!
0%
#423915000000
1!
1%
#423920000000
0!
0%
#423925000000
1!
1%
#423930000000
0!
0%
#423935000000
1!
1%
#423940000000
0!
0%
#423945000000
1!
1%
#423950000000
0!
0%
#423955000000
1!
1%
#423960000000
0!
0%
#423965000000
1!
1%
#423970000000
0!
0%
#423975000000
1!
1%
#423980000000
0!
0%
#423985000000
1!
1%
#423990000000
0!
0%
#423995000000
1!
1%
#424000000000
0!
0%
#424005000000
1!
1%
#424010000000
0!
0%
#424015000000
1!
1%
#424020000000
0!
0%
#424025000000
1!
1%
#424030000000
0!
0%
#424035000000
1!
1%
#424040000000
0!
0%
#424045000000
1!
1%
#424050000000
0!
0%
#424055000000
1!
1%
#424060000000
0!
0%
#424065000000
1!
1%
#424070000000
0!
0%
#424075000000
1!
1%
#424080000000
0!
0%
#424085000000
1!
1%
#424090000000
0!
0%
#424095000000
1!
1%
#424100000000
0!
0%
#424105000000
1!
1%
#424110000000
0!
0%
#424115000000
1!
1%
#424120000000
0!
0%
#424125000000
1!
1%
#424130000000
0!
0%
#424135000000
1!
1%
#424140000000
0!
0%
#424145000000
1!
1%
#424150000000
0!
0%
#424155000000
1!
1%
#424160000000
0!
0%
#424165000000
1!
1%
#424170000000
0!
0%
#424175000000
1!
1%
#424180000000
0!
0%
#424185000000
1!
1%
#424190000000
0!
0%
#424195000000
1!
1%
#424200000000
0!
0%
#424205000000
1!
1%
#424210000000
0!
0%
#424215000000
1!
1%
#424220000000
0!
0%
#424225000000
1!
1%
#424230000000
0!
0%
#424235000000
1!
1%
#424240000000
0!
0%
#424245000000
1!
1%
#424250000000
0!
0%
#424255000000
1!
1%
#424260000000
0!
0%
#424265000000
1!
1%
#424270000000
0!
0%
#424275000000
1!
1%
#424280000000
0!
0%
#424285000000
1!
1%
#424290000000
0!
0%
#424295000000
1!
1%
#424300000000
0!
0%
#424305000000
1!
1%
#424310000000
0!
0%
#424315000000
1!
1%
#424320000000
0!
0%
#424325000000
1!
1%
#424330000000
0!
0%
#424335000000
1!
1%
#424340000000
0!
0%
#424345000000
1!
1%
#424350000000
0!
0%
#424355000000
1!
1%
#424360000000
0!
0%
#424365000000
1!
1%
#424370000000
0!
0%
#424375000000
1!
1%
#424380000000
0!
0%
#424385000000
1!
1%
#424390000000
0!
0%
#424395000000
1!
1%
#424400000000
0!
0%
#424405000000
1!
1%
#424410000000
0!
0%
#424415000000
1!
1%
#424420000000
0!
0%
#424425000000
1!
1%
#424430000000
0!
0%
#424435000000
1!
1%
#424440000000
0!
0%
#424445000000
1!
1%
#424450000000
0!
0%
#424455000000
1!
1%
#424460000000
0!
0%
#424465000000
1!
1%
#424470000000
0!
0%
#424475000000
1!
1%
#424480000000
0!
0%
#424485000000
1!
1%
#424490000000
0!
0%
#424495000000
1!
1%
#424500000000
0!
0%
#424505000000
1!
1%
#424510000000
0!
0%
#424515000000
1!
1%
#424520000000
0!
0%
#424525000000
1!
1%
#424530000000
0!
0%
#424535000000
1!
1%
#424540000000
0!
0%
#424545000000
1!
1%
#424550000000
0!
0%
#424555000000
1!
1%
#424560000000
0!
0%
#424565000000
1!
1%
#424570000000
0!
0%
#424575000000
1!
1%
#424580000000
0!
0%
#424585000000
1!
1%
#424590000000
0!
0%
#424595000000
1!
1%
#424600000000
0!
0%
#424605000000
1!
1%
#424610000000
0!
0%
#424615000000
1!
1%
#424620000000
0!
0%
#424625000000
1!
1%
#424630000000
0!
0%
#424635000000
1!
1%
#424640000000
0!
0%
#424645000000
1!
1%
#424650000000
0!
0%
#424655000000
1!
1%
#424660000000
0!
0%
#424665000000
1!
1%
#424670000000
0!
0%
#424675000000
1!
1%
#424680000000
0!
0%
#424685000000
1!
1%
#424690000000
0!
0%
#424695000000
1!
1%
#424700000000
0!
0%
#424705000000
1!
1%
#424710000000
0!
0%
#424715000000
1!
1%
#424720000000
0!
0%
#424725000000
1!
1%
#424730000000
0!
0%
#424735000000
1!
1%
#424740000000
0!
0%
#424745000000
1!
1%
#424750000000
0!
0%
#424755000000
1!
1%
#424760000000
0!
0%
#424765000000
1!
1%
#424770000000
0!
0%
#424775000000
1!
1%
#424780000000
0!
0%
#424785000000
1!
1%
#424790000000
0!
0%
#424795000000
1!
1%
#424800000000
0!
0%
#424805000000
1!
1%
#424810000000
0!
0%
#424815000000
1!
1%
#424820000000
0!
0%
#424825000000
1!
1%
#424830000000
0!
0%
#424835000000
1!
1%
#424840000000
0!
0%
#424845000000
1!
1%
#424850000000
0!
0%
#424855000000
1!
1%
#424860000000
0!
0%
#424865000000
1!
1%
#424870000000
0!
0%
#424875000000
1!
1%
#424880000000
0!
0%
#424885000000
1!
1%
#424890000000
0!
0%
#424895000000
1!
1%
#424900000000
0!
0%
#424905000000
1!
1%
#424910000000
0!
0%
#424915000000
1!
1%
#424920000000
0!
0%
#424925000000
1!
1%
#424930000000
0!
0%
#424935000000
1!
1%
#424940000000
0!
0%
#424945000000
1!
1%
#424950000000
0!
0%
#424955000000
1!
1%
#424960000000
0!
0%
#424965000000
1!
1%
#424970000000
0!
0%
#424975000000
1!
1%
#424980000000
0!
0%
#424985000000
1!
1%
#424990000000
0!
0%
#424995000000
1!
1%
#425000000000
0!
0%
#425005000000
1!
1%
#425010000000
0!
0%
#425015000000
1!
1%
#425020000000
0!
0%
#425025000000
1!
1%
#425030000000
0!
0%
#425035000000
1!
1%
#425040000000
0!
0%
#425045000000
1!
1%
#425050000000
0!
0%
#425055000000
1!
1%
#425060000000
0!
0%
#425065000000
1!
1%
#425070000000
0!
0%
#425075000000
1!
1%
#425080000000
0!
0%
#425085000000
1!
1%
#425090000000
0!
0%
#425095000000
1!
1%
#425100000000
0!
0%
#425105000000
1!
1%
#425110000000
0!
0%
#425115000000
1!
1%
#425120000000
0!
0%
#425125000000
1!
1%
#425130000000
0!
0%
#425135000000
1!
1%
#425140000000
0!
0%
#425145000000
1!
1%
#425150000000
0!
0%
#425155000000
1!
1%
#425160000000
0!
0%
#425165000000
1!
1%
#425170000000
0!
0%
#425175000000
1!
1%
#425180000000
0!
0%
#425185000000
1!
1%
#425190000000
0!
0%
#425195000000
1!
1%
#425200000000
0!
0%
#425205000000
1!
1%
#425210000000
0!
0%
#425215000000
1!
1%
#425220000000
0!
0%
#425225000000
1!
1%
#425230000000
0!
0%
#425235000000
1!
1%
#425240000000
0!
0%
#425245000000
1!
1%
#425250000000
0!
0%
#425255000000
1!
1%
#425260000000
0!
0%
#425265000000
1!
1%
#425270000000
0!
0%
#425275000000
1!
1%
#425280000000
0!
0%
#425285000000
1!
1%
#425290000000
0!
0%
#425295000000
1!
1%
#425300000000
0!
0%
#425305000000
1!
1%
#425310000000
0!
0%
#425315000000
1!
1%
#425320000000
0!
0%
#425325000000
1!
1%
#425330000000
0!
0%
#425335000000
1!
1%
#425340000000
0!
0%
#425345000000
1!
1%
#425350000000
0!
0%
#425355000000
1!
1%
#425360000000
0!
0%
#425365000000
1!
1%
#425370000000
0!
0%
#425375000000
1!
1%
#425380000000
0!
0%
#425385000000
1!
1%
#425390000000
0!
0%
#425395000000
1!
1%
#425400000000
0!
0%
#425405000000
1!
1%
#425410000000
0!
0%
#425415000000
1!
1%
#425420000000
0!
0%
#425425000000
1!
1%
#425430000000
0!
0%
#425435000000
1!
1%
#425440000000
0!
0%
#425445000000
1!
1%
#425450000000
0!
0%
#425455000000
1!
1%
#425460000000
0!
0%
#425465000000
1!
1%
#425470000000
0!
0%
#425475000000
1!
1%
#425480000000
0!
0%
#425485000000
1!
1%
#425490000000
0!
0%
#425495000000
1!
1%
#425500000000
0!
0%
#425505000000
1!
1%
#425510000000
0!
0%
#425515000000
1!
1%
#425520000000
0!
0%
#425525000000
1!
1%
#425530000000
0!
0%
#425535000000
1!
1%
#425540000000
0!
0%
#425545000000
1!
1%
#425550000000
0!
0%
#425555000000
1!
1%
#425560000000
0!
0%
#425565000000
1!
1%
#425570000000
0!
0%
#425575000000
1!
1%
#425580000000
0!
0%
#425585000000
1!
1%
#425590000000
0!
0%
#425595000000
1!
1%
#425600000000
0!
0%
#425605000000
1!
1%
#425610000000
0!
0%
#425615000000
1!
1%
#425620000000
0!
0%
#425625000000
1!
1%
#425630000000
0!
0%
#425635000000
1!
1%
#425640000000
0!
0%
#425645000000
1!
1%
#425650000000
0!
0%
#425655000000
1!
1%
#425660000000
0!
0%
#425665000000
1!
1%
#425670000000
0!
0%
#425675000000
1!
1%
#425680000000
0!
0%
#425685000000
1!
1%
#425690000000
0!
0%
#425695000000
1!
1%
#425700000000
0!
0%
#425705000000
1!
1%
#425710000000
0!
0%
#425715000000
1!
1%
#425720000000
0!
0%
#425725000000
1!
1%
#425730000000
0!
0%
#425735000000
1!
1%
#425740000000
0!
0%
#425745000000
1!
1%
#425750000000
0!
0%
#425755000000
1!
1%
#425760000000
0!
0%
#425765000000
1!
1%
#425770000000
0!
0%
#425775000000
1!
1%
#425780000000
0!
0%
#425785000000
1!
1%
#425790000000
0!
0%
#425795000000
1!
1%
#425800000000
0!
0%
#425805000000
1!
1%
#425810000000
0!
0%
#425815000000
1!
1%
#425820000000
0!
0%
#425825000000
1!
1%
#425830000000
0!
0%
#425835000000
1!
1%
#425840000000
0!
0%
#425845000000
1!
1%
#425850000000
0!
0%
#425855000000
1!
1%
#425860000000
0!
0%
#425865000000
1!
1%
#425870000000
0!
0%
#425875000000
1!
1%
#425880000000
0!
0%
#425885000000
1!
1%
#425890000000
0!
0%
#425895000000
1!
1%
#425900000000
0!
0%
#425905000000
1!
1%
#425910000000
0!
0%
#425915000000
1!
1%
#425920000000
0!
0%
#425925000000
1!
1%
#425930000000
0!
0%
#425935000000
1!
1%
#425940000000
0!
0%
#425945000000
1!
1%
#425950000000
0!
0%
#425955000000
1!
1%
#425960000000
0!
0%
#425965000000
1!
1%
#425970000000
0!
0%
#425975000000
1!
1%
#425980000000
0!
0%
#425985000000
1!
1%
#425990000000
0!
0%
#425995000000
1!
1%
#426000000000
0!
0%
#426005000000
1!
1%
#426010000000
0!
0%
#426015000000
1!
1%
#426020000000
0!
0%
#426025000000
1!
1%
#426030000000
0!
0%
#426035000000
1!
1%
#426040000000
0!
0%
#426045000000
1!
1%
#426050000000
0!
0%
#426055000000
1!
1%
#426060000000
0!
0%
#426065000000
1!
1%
#426070000000
0!
0%
#426075000000
1!
1%
#426080000000
0!
0%
#426085000000
1!
1%
#426090000000
0!
0%
#426095000000
1!
1%
#426100000000
0!
0%
#426105000000
1!
1%
#426110000000
0!
0%
#426115000000
1!
1%
#426120000000
0!
0%
#426125000000
1!
1%
#426130000000
0!
0%
#426135000000
1!
1%
#426140000000
0!
0%
#426145000000
1!
1%
#426150000000
0!
0%
#426155000000
1!
1%
#426160000000
0!
0%
#426165000000
1!
1%
#426170000000
0!
0%
#426175000000
1!
1%
#426180000000
0!
0%
#426185000000
1!
1%
#426190000000
0!
0%
#426195000000
1!
1%
#426200000000
0!
0%
#426205000000
1!
1%
#426210000000
0!
0%
#426215000000
1!
1%
#426220000000
0!
0%
#426225000000
1!
1%
#426230000000
0!
0%
#426235000000
1!
1%
#426240000000
0!
0%
#426245000000
1!
1%
#426250000000
0!
0%
#426255000000
1!
1%
#426260000000
0!
0%
#426265000000
1!
1%
#426270000000
0!
0%
#426275000000
1!
1%
#426280000000
0!
0%
#426285000000
1!
1%
#426290000000
0!
0%
#426295000000
1!
1%
#426300000000
0!
0%
#426305000000
1!
1%
#426310000000
0!
0%
#426315000000
1!
1%
#426320000000
0!
0%
#426325000000
1!
1%
#426330000000
0!
0%
#426335000000
1!
1%
#426340000000
0!
0%
#426345000000
1!
1%
#426350000000
0!
0%
#426355000000
1!
1%
#426360000000
0!
0%
#426365000000
1!
1%
#426370000000
0!
0%
#426375000000
1!
1%
#426380000000
0!
0%
#426385000000
1!
1%
#426390000000
0!
0%
#426395000000
1!
1%
#426400000000
0!
0%
#426405000000
1!
1%
#426410000000
0!
0%
#426415000000
1!
1%
#426420000000
0!
0%
#426425000000
1!
1%
#426430000000
0!
0%
#426435000000
1!
1%
#426440000000
0!
0%
#426445000000
1!
1%
#426450000000
0!
0%
#426455000000
1!
1%
#426460000000
0!
0%
#426465000000
1!
1%
#426470000000
0!
0%
#426475000000
1!
1%
#426480000000
0!
0%
#426485000000
1!
1%
#426490000000
0!
0%
#426495000000
1!
1%
#426500000000
0!
0%
#426505000000
1!
1%
#426510000000
0!
0%
#426515000000
1!
1%
#426520000000
0!
0%
#426525000000
1!
1%
#426530000000
0!
0%
#426535000000
1!
1%
#426540000000
0!
0%
#426545000000
1!
1%
#426550000000
0!
0%
#426555000000
1!
1%
#426560000000
0!
0%
#426565000000
1!
1%
#426570000000
0!
0%
#426575000000
1!
1%
#426580000000
0!
0%
#426585000000
1!
1%
#426590000000
0!
0%
#426595000000
1!
1%
#426600000000
0!
0%
#426605000000
1!
1%
#426610000000
0!
0%
#426615000000
1!
1%
#426620000000
0!
0%
#426625000000
1!
1%
#426630000000
0!
0%
#426635000000
1!
1%
#426640000000
0!
0%
#426645000000
1!
1%
#426650000000
0!
0%
#426655000000
1!
1%
#426660000000
0!
0%
#426665000000
1!
1%
#426670000000
0!
0%
#426675000000
1!
1%
#426680000000
0!
0%
#426685000000
1!
1%
#426690000000
0!
0%
#426695000000
1!
1%
#426700000000
0!
0%
#426705000000
1!
1%
#426710000000
0!
0%
#426715000000
1!
1%
#426720000000
0!
0%
#426725000000
1!
1%
#426730000000
0!
0%
#426735000000
1!
1%
#426740000000
0!
0%
#426745000000
1!
1%
#426750000000
0!
0%
#426755000000
1!
1%
#426760000000
0!
0%
#426765000000
1!
1%
#426770000000
0!
0%
#426775000000
1!
1%
#426780000000
0!
0%
#426785000000
1!
1%
#426790000000
0!
0%
#426795000000
1!
1%
#426800000000
0!
0%
#426805000000
1!
1%
#426810000000
0!
0%
#426815000000
1!
1%
#426820000000
0!
0%
#426825000000
1!
1%
#426830000000
0!
0%
#426835000000
1!
1%
#426840000000
0!
0%
#426845000000
1!
1%
#426850000000
0!
0%
#426855000000
1!
1%
#426860000000
0!
0%
#426865000000
1!
1%
#426870000000
0!
0%
#426875000000
1!
1%
#426880000000
0!
0%
#426885000000
1!
1%
#426890000000
0!
0%
#426895000000
1!
1%
#426900000000
0!
0%
#426905000000
1!
1%
#426910000000
0!
0%
#426915000000
1!
1%
#426920000000
0!
0%
#426925000000
1!
1%
#426930000000
0!
0%
#426935000000
1!
1%
#426940000000
0!
0%
#426945000000
1!
1%
#426950000000
0!
0%
#426955000000
1!
1%
#426960000000
0!
0%
#426965000000
1!
1%
#426970000000
0!
0%
#426975000000
1!
1%
#426980000000
0!
0%
#426985000000
1!
1%
#426990000000
0!
0%
#426995000000
1!
1%
#427000000000
0!
0%
#427005000000
1!
1%
#427010000000
0!
0%
#427015000000
1!
1%
#427020000000
0!
0%
#427025000000
1!
1%
#427030000000
0!
0%
#427035000000
1!
1%
#427040000000
0!
0%
#427045000000
1!
1%
#427050000000
0!
0%
#427055000000
1!
1%
#427060000000
0!
0%
#427065000000
1!
1%
#427070000000
0!
0%
#427075000000
1!
1%
#427080000000
0!
0%
#427085000000
1!
1%
#427090000000
0!
0%
#427095000000
1!
1%
#427100000000
0!
0%
#427105000000
1!
1%
#427110000000
0!
0%
#427115000000
1!
1%
#427120000000
0!
0%
#427125000000
1!
1%
#427130000000
0!
0%
#427135000000
1!
1%
#427140000000
0!
0%
#427145000000
1!
1%
#427150000000
0!
0%
#427155000000
1!
1%
#427160000000
0!
0%
#427165000000
1!
1%
#427170000000
0!
0%
#427175000000
1!
1%
#427180000000
0!
0%
#427185000000
1!
1%
#427190000000
0!
0%
#427195000000
1!
1%
#427200000000
0!
0%
#427205000000
1!
1%
#427210000000
0!
0%
#427215000000
1!
1%
#427220000000
0!
0%
#427225000000
1!
1%
#427230000000
0!
0%
#427235000000
1!
1%
#427240000000
0!
0%
#427245000000
1!
1%
#427250000000
0!
0%
#427255000000
1!
1%
#427260000000
0!
0%
#427265000000
1!
1%
#427270000000
0!
0%
#427275000000
1!
1%
#427280000000
0!
0%
#427285000000
1!
1%
#427290000000
0!
0%
#427295000000
1!
1%
#427300000000
0!
0%
#427305000000
1!
1%
#427310000000
0!
0%
#427315000000
1!
1%
#427320000000
0!
0%
#427325000000
1!
1%
#427330000000
0!
0%
#427335000000
1!
1%
#427340000000
0!
0%
#427345000000
1!
1%
#427350000000
0!
0%
#427355000000
1!
1%
#427360000000
0!
0%
#427365000000
1!
1%
#427370000000
0!
0%
#427375000000
1!
1%
#427380000000
0!
0%
#427385000000
1!
1%
#427390000000
0!
0%
#427395000000
1!
1%
#427400000000
0!
0%
#427405000000
1!
1%
#427410000000
0!
0%
#427415000000
1!
1%
#427420000000
0!
0%
#427425000000
1!
1%
#427430000000
0!
0%
#427435000000
1!
1%
#427440000000
0!
0%
#427445000000
1!
1%
#427450000000
0!
0%
#427455000000
1!
1%
#427460000000
0!
0%
#427465000000
1!
1%
#427470000000
0!
0%
#427475000000
1!
1%
#427480000000
0!
0%
#427485000000
1!
1%
#427490000000
0!
0%
#427495000000
1!
1%
#427500000000
0!
0%
#427505000000
1!
1%
#427510000000
0!
0%
#427515000000
1!
1%
#427520000000
0!
0%
#427525000000
1!
1%
#427530000000
0!
0%
#427535000000
1!
1%
#427540000000
0!
0%
#427545000000
1!
1%
#427550000000
0!
0%
#427555000000
1!
1%
#427560000000
0!
0%
#427565000000
1!
1%
#427570000000
0!
0%
#427575000000
1!
1%
#427580000000
0!
0%
#427585000000
1!
1%
#427590000000
0!
0%
#427595000000
1!
1%
#427600000000
0!
0%
#427605000000
1!
1%
#427610000000
0!
0%
#427615000000
1!
1%
#427620000000
0!
0%
#427625000000
1!
1%
#427630000000
0!
0%
#427635000000
1!
1%
#427640000000
0!
0%
#427645000000
1!
1%
#427650000000
0!
0%
#427655000000
1!
1%
#427660000000
0!
0%
#427665000000
1!
1%
#427670000000
0!
0%
#427675000000
1!
1%
#427680000000
0!
0%
#427685000000
1!
1%
#427690000000
0!
0%
#427695000000
1!
1%
#427700000000
0!
0%
#427705000000
1!
1%
#427710000000
0!
0%
#427715000000
1!
1%
#427720000000
0!
0%
#427725000000
1!
1%
#427730000000
0!
0%
#427735000000
1!
1%
#427740000000
0!
0%
#427745000000
1!
1%
#427750000000
0!
0%
#427755000000
1!
1%
#427760000000
0!
0%
#427765000000
1!
1%
#427770000000
0!
0%
#427775000000
1!
1%
#427780000000
0!
0%
#427785000000
1!
1%
#427790000000
0!
0%
#427795000000
1!
1%
#427800000000
0!
0%
#427805000000
1!
1%
#427810000000
0!
0%
#427815000000
1!
1%
#427820000000
0!
0%
#427825000000
1!
1%
#427830000000
0!
0%
#427835000000
1!
1%
#427840000000
0!
0%
#427845000000
1!
1%
#427850000000
0!
0%
#427855000000
1!
1%
#427860000000
0!
0%
#427865000000
1!
1%
#427870000000
0!
0%
#427875000000
1!
1%
#427880000000
0!
0%
#427885000000
1!
1%
#427890000000
0!
0%
#427895000000
1!
1%
#427900000000
0!
0%
#427905000000
1!
1%
#427910000000
0!
0%
#427915000000
1!
1%
#427920000000
0!
0%
#427925000000
1!
1%
#427930000000
0!
0%
#427935000000
1!
1%
#427940000000
0!
0%
#427945000000
1!
1%
#427950000000
0!
0%
#427955000000
1!
1%
#427960000000
0!
0%
#427965000000
1!
1%
#427970000000
0!
0%
#427975000000
1!
1%
#427980000000
0!
0%
#427985000000
1!
1%
#427990000000
0!
0%
#427995000000
1!
1%
#428000000000
0!
0%
#428005000000
1!
1%
#428010000000
0!
0%
#428015000000
1!
1%
#428020000000
0!
0%
#428025000000
1!
1%
#428030000000
0!
0%
#428035000000
1!
1%
#428040000000
0!
0%
#428045000000
1!
1%
#428050000000
0!
0%
#428055000000
1!
1%
#428060000000
0!
0%
#428065000000
1!
1%
#428070000000
0!
0%
#428075000000
1!
1%
#428080000000
0!
0%
#428085000000
1!
1%
#428090000000
0!
0%
#428095000000
1!
1%
#428100000000
0!
0%
#428105000000
1!
1%
#428110000000
0!
0%
#428115000000
1!
1%
#428120000000
0!
0%
#428125000000
1!
1%
#428130000000
0!
0%
#428135000000
1!
1%
#428140000000
0!
0%
#428145000000
1!
1%
#428150000000
0!
0%
#428155000000
1!
1%
#428160000000
0!
0%
#428165000000
1!
1%
#428170000000
0!
0%
#428175000000
1!
1%
#428180000000
0!
0%
#428185000000
1!
1%
#428190000000
0!
0%
#428195000000
1!
1%
#428200000000
0!
0%
#428205000000
1!
1%
#428210000000
0!
0%
#428215000000
1!
1%
#428220000000
0!
0%
#428225000000
1!
1%
#428230000000
0!
0%
#428235000000
1!
1%
#428240000000
0!
0%
#428245000000
1!
1%
#428250000000
0!
0%
#428255000000
1!
1%
#428260000000
0!
0%
#428265000000
1!
1%
#428270000000
0!
0%
#428275000000
1!
1%
#428280000000
0!
0%
#428285000000
1!
1%
#428290000000
0!
0%
#428295000000
1!
1%
#428300000000
0!
0%
#428305000000
1!
1%
#428310000000
0!
0%
#428315000000
1!
1%
#428320000000
0!
0%
#428325000000
1!
1%
#428330000000
0!
0%
#428335000000
1!
1%
#428340000000
0!
0%
#428345000000
1!
1%
#428350000000
0!
0%
#428355000000
1!
1%
#428360000000
0!
0%
#428365000000
1!
1%
#428370000000
0!
0%
#428375000000
1!
1%
#428380000000
0!
0%
#428385000000
1!
1%
#428390000000
0!
0%
#428395000000
1!
1%
#428400000000
0!
0%
#428405000000
1!
1%
#428410000000
0!
0%
#428415000000
1!
1%
#428420000000
0!
0%
#428425000000
1!
1%
#428430000000
0!
0%
#428435000000
1!
1%
#428440000000
0!
0%
#428445000000
1!
1%
#428450000000
0!
0%
#428455000000
1!
1%
#428460000000
0!
0%
#428465000000
1!
1%
#428470000000
0!
0%
#428475000000
1!
1%
#428480000000
0!
0%
#428485000000
1!
1%
#428490000000
0!
0%
#428495000000
1!
1%
#428500000000
0!
0%
#428505000000
1!
1%
#428510000000
0!
0%
#428515000000
1!
1%
#428520000000
0!
0%
#428525000000
1!
1%
#428530000000
0!
0%
#428535000000
1!
1%
#428540000000
0!
0%
#428545000000
1!
1%
#428550000000
0!
0%
#428555000000
1!
1%
#428560000000
0!
0%
#428565000000
1!
1%
#428570000000
0!
0%
#428575000000
1!
1%
#428580000000
0!
0%
#428585000000
1!
1%
#428590000000
0!
0%
#428595000000
1!
1%
#428600000000
0!
0%
#428605000000
1!
1%
#428610000000
0!
0%
#428615000000
1!
1%
#428620000000
0!
0%
#428625000000
1!
1%
#428630000000
0!
0%
#428635000000
1!
1%
#428640000000
0!
0%
#428645000000
1!
1%
#428650000000
0!
0%
#428655000000
1!
1%
#428660000000
0!
0%
#428665000000
1!
1%
#428670000000
0!
0%
#428675000000
1!
1%
#428680000000
0!
0%
#428685000000
1!
1%
#428690000000
0!
0%
#428695000000
1!
1%
#428700000000
0!
0%
#428705000000
1!
1%
#428710000000
0!
0%
#428715000000
1!
1%
#428720000000
0!
0%
#428725000000
1!
1%
#428730000000
0!
0%
#428735000000
1!
1%
#428740000000
0!
0%
#428745000000
1!
1%
#428750000000
0!
0%
#428755000000
1!
1%
#428760000000
0!
0%
#428765000000
1!
1%
#428770000000
0!
0%
#428775000000
1!
1%
#428780000000
0!
0%
#428785000000
1!
1%
#428790000000
0!
0%
#428795000000
1!
1%
#428800000000
0!
0%
#428805000000
1!
1%
#428810000000
0!
0%
#428815000000
1!
1%
#428820000000
0!
0%
#428825000000
1!
1%
#428830000000
0!
0%
#428835000000
1!
1%
#428840000000
0!
0%
#428845000000
1!
1%
#428850000000
0!
0%
#428855000000
1!
1%
#428860000000
0!
0%
#428865000000
1!
1%
#428870000000
0!
0%
#428875000000
1!
1%
#428880000000
0!
0%
#428885000000
1!
1%
#428890000000
0!
0%
#428895000000
1!
1%
#428900000000
0!
0%
#428905000000
1!
1%
#428910000000
0!
0%
#428915000000
1!
1%
#428920000000
0!
0%
#428925000000
1!
1%
#428930000000
0!
0%
#428935000000
1!
1%
#428940000000
0!
0%
#428945000000
1!
1%
#428950000000
0!
0%
#428955000000
1!
1%
#428960000000
0!
0%
#428965000000
1!
1%
#428970000000
0!
0%
#428975000000
1!
1%
#428980000000
0!
0%
#428985000000
1!
1%
#428990000000
0!
0%
#428995000000
1!
1%
#429000000000
0!
0%
#429005000000
1!
1%
#429010000000
0!
0%
#429015000000
1!
1%
#429020000000
0!
0%
#429025000000
1!
1%
#429030000000
0!
0%
#429035000000
1!
1%
#429040000000
0!
0%
#429045000000
1!
1%
#429050000000
0!
0%
#429055000000
1!
1%
#429060000000
0!
0%
#429065000000
1!
1%
#429070000000
0!
0%
#429075000000
1!
1%
#429080000000
0!
0%
#429085000000
1!
1%
#429090000000
0!
0%
#429095000000
1!
1%
#429100000000
0!
0%
#429105000000
1!
1%
#429110000000
0!
0%
#429115000000
1!
1%
#429120000000
0!
0%
#429125000000
1!
1%
#429130000000
0!
0%
#429135000000
1!
1%
#429140000000
0!
0%
#429145000000
1!
1%
#429150000000
0!
0%
#429155000000
1!
1%
#429160000000
0!
0%
#429165000000
1!
1%
#429170000000
0!
0%
#429175000000
1!
1%
#429180000000
0!
0%
#429185000000
1!
1%
#429190000000
0!
0%
#429195000000
1!
1%
#429200000000
0!
0%
#429205000000
1!
1%
#429210000000
0!
0%
#429215000000
1!
1%
#429220000000
0!
0%
#429225000000
1!
1%
#429230000000
0!
0%
#429235000000
1!
1%
#429240000000
0!
0%
#429245000000
1!
1%
#429250000000
0!
0%
#429255000000
1!
1%
#429260000000
0!
0%
#429265000000
1!
1%
#429270000000
0!
0%
#429275000000
1!
1%
#429280000000
0!
0%
#429285000000
1!
1%
#429290000000
0!
0%
#429295000000
1!
1%
#429300000000
0!
0%
#429305000000
1!
1%
#429310000000
0!
0%
#429315000000
1!
1%
#429320000000
0!
0%
#429325000000
1!
1%
#429330000000
0!
0%
#429335000000
1!
1%
#429340000000
0!
0%
#429345000000
1!
1%
#429350000000
0!
0%
#429355000000
1!
1%
#429360000000
0!
0%
#429365000000
1!
1%
#429370000000
0!
0%
#429375000000
1!
1%
#429380000000
0!
0%
#429385000000
1!
1%
#429390000000
0!
0%
#429395000000
1!
1%
#429400000000
0!
0%
#429405000000
1!
1%
#429410000000
0!
0%
#429415000000
1!
1%
#429420000000
0!
0%
#429425000000
1!
1%
#429430000000
0!
0%
#429435000000
1!
1%
#429440000000
0!
0%
#429445000000
1!
1%
#429450000000
0!
0%
#429455000000
1!
1%
#429460000000
0!
0%
#429465000000
1!
1%
#429470000000
0!
0%
#429475000000
1!
1%
#429480000000
0!
0%
#429485000000
1!
1%
#429490000000
0!
0%
#429495000000
1!
1%
#429500000000
0!
0%
#429505000000
1!
1%
#429510000000
0!
0%
#429515000000
1!
1%
#429520000000
0!
0%
#429525000000
1!
1%
#429530000000
0!
0%
#429535000000
1!
1%
#429540000000
0!
0%
#429545000000
1!
1%
#429550000000
0!
0%
#429555000000
1!
1%
#429560000000
0!
0%
#429565000000
1!
1%
#429570000000
0!
0%
#429575000000
1!
1%
#429580000000
0!
0%
#429585000000
1!
1%
#429590000000
0!
0%
#429595000000
1!
1%
#429600000000
0!
0%
#429605000000
1!
1%
#429610000000
0!
0%
#429615000000
1!
1%
#429620000000
0!
0%
#429625000000
1!
1%
#429630000000
0!
0%
#429635000000
1!
1%
#429640000000
0!
0%
#429645000000
1!
1%
#429650000000
0!
0%
#429655000000
1!
1%
#429660000000
0!
0%
#429665000000
1!
1%
#429670000000
0!
0%
#429675000000
1!
1%
#429680000000
0!
0%
#429685000000
1!
1%
#429690000000
0!
0%
#429695000000
1!
1%
#429700000000
0!
0%
#429705000000
1!
1%
#429710000000
0!
0%
#429715000000
1!
1%
#429720000000
0!
0%
#429725000000
1!
1%
#429730000000
0!
0%
#429735000000
1!
1%
#429740000000
0!
0%
#429745000000
1!
1%
#429750000000
0!
0%
#429755000000
1!
1%
#429760000000
0!
0%
#429765000000
1!
1%
#429770000000
0!
0%
#429775000000
1!
1%
#429780000000
0!
0%
#429785000000
1!
1%
#429790000000
0!
0%
#429795000000
1!
1%
#429800000000
0!
0%
#429805000000
1!
1%
#429810000000
0!
0%
#429815000000
1!
1%
#429820000000
0!
0%
#429825000000
1!
1%
#429830000000
0!
0%
#429835000000
1!
1%
#429840000000
0!
0%
#429845000000
1!
1%
#429850000000
0!
0%
#429855000000
1!
1%
#429860000000
0!
0%
#429865000000
1!
1%
#429870000000
0!
0%
#429875000000
1!
1%
#429880000000
0!
0%
#429885000000
1!
1%
#429890000000
0!
0%
#429895000000
1!
1%
#429900000000
0!
0%
#429905000000
1!
1%
#429910000000
0!
0%
#429915000000
1!
1%
#429920000000
0!
0%
#429925000000
1!
1%
#429930000000
0!
0%
#429935000000
1!
1%
#429940000000
0!
0%
#429945000000
1!
1%
#429950000000
0!
0%
#429955000000
1!
1%
#429960000000
0!
0%
#429965000000
1!
1%
#429970000000
0!
0%
#429975000000
1!
1%
#429980000000
0!
0%
#429985000000
1!
1%
#429990000000
0!
0%
#429995000000
1!
1%
#430000000000
0!
0%
#430005000000
1!
1%
#430010000000
0!
0%
#430015000000
1!
1%
#430020000000
0!
0%
#430025000000
1!
1%
#430030000000
0!
0%
#430035000000
1!
1%
#430040000000
0!
0%
#430045000000
1!
1%
#430050000000
0!
0%
#430055000000
1!
1%
#430060000000
0!
0%
#430065000000
1!
1%
#430070000000
0!
0%
#430075000000
1!
1%
#430080000000
0!
0%
#430085000000
1!
1%
#430090000000
0!
0%
#430095000000
1!
1%
#430100000000
0!
0%
#430105000000
1!
1%
#430110000000
0!
0%
#430115000000
1!
1%
#430120000000
0!
0%
#430125000000
1!
1%
#430130000000
0!
0%
#430135000000
1!
1%
#430140000000
0!
0%
#430145000000
1!
1%
#430150000000
0!
0%
#430155000000
1!
1%
#430160000000
0!
0%
#430165000000
1!
1%
#430170000000
0!
0%
#430175000000
1!
1%
#430180000000
0!
0%
#430185000000
1!
1%
#430190000000
0!
0%
#430195000000
1!
1%
#430200000000
0!
0%
#430205000000
1!
1%
#430210000000
0!
0%
#430215000000
1!
1%
#430220000000
0!
0%
#430225000000
1!
1%
#430230000000
0!
0%
#430235000000
1!
1%
#430240000000
0!
0%
#430245000000
1!
1%
#430250000000
0!
0%
#430255000000
1!
1%
#430260000000
0!
0%
#430265000000
1!
1%
#430270000000
0!
0%
#430275000000
1!
1%
#430280000000
0!
0%
#430285000000
1!
1%
#430290000000
0!
0%
#430295000000
1!
1%
#430300000000
0!
0%
#430305000000
1!
1%
#430310000000
0!
0%
#430315000000
1!
1%
#430320000000
0!
0%
#430325000000
1!
1%
#430330000000
0!
0%
#430335000000
1!
1%
#430340000000
0!
0%
#430345000000
1!
1%
#430350000000
0!
0%
#430355000000
1!
1%
#430360000000
0!
0%
#430365000000
1!
1%
#430370000000
0!
0%
#430375000000
1!
1%
#430380000000
0!
0%
#430385000000
1!
1%
#430390000000
0!
0%
#430395000000
1!
1%
#430400000000
0!
0%
#430405000000
1!
1%
#430410000000
0!
0%
#430415000000
1!
1%
#430420000000
0!
0%
#430425000000
1!
1%
#430430000000
0!
0%
#430435000000
1!
1%
#430440000000
0!
0%
#430445000000
1!
1%
#430450000000
0!
0%
#430455000000
1!
1%
#430460000000
0!
0%
#430465000000
1!
1%
#430470000000
0!
0%
#430475000000
1!
1%
#430480000000
0!
0%
#430485000000
1!
1%
#430490000000
0!
0%
#430495000000
1!
1%
#430500000000
0!
0%
#430505000000
1!
1%
#430510000000
0!
0%
#430515000000
1!
1%
#430520000000
0!
0%
#430525000000
1!
1%
#430530000000
0!
0%
#430535000000
1!
1%
#430540000000
0!
0%
#430545000000
1!
1%
#430550000000
0!
0%
#430555000000
1!
1%
#430560000000
0!
0%
#430565000000
1!
1%
#430570000000
0!
0%
#430575000000
1!
1%
#430580000000
0!
0%
#430585000000
1!
1%
#430590000000
0!
0%
#430595000000
1!
1%
#430600000000
0!
0%
#430605000000
1!
1%
#430610000000
0!
0%
#430615000000
1!
1%
#430620000000
0!
0%
#430625000000
1!
1%
#430630000000
0!
0%
#430635000000
1!
1%
#430640000000
0!
0%
#430645000000
1!
1%
#430650000000
0!
0%
#430655000000
1!
1%
#430660000000
0!
0%
#430665000000
1!
1%
#430670000000
0!
0%
#430675000000
1!
1%
#430680000000
0!
0%
#430685000000
1!
1%
#430690000000
0!
0%
#430695000000
1!
1%
#430700000000
0!
0%
#430705000000
1!
1%
#430710000000
0!
0%
#430715000000
1!
1%
#430720000000
0!
0%
#430725000000
1!
1%
#430730000000
0!
0%
#430735000000
1!
1%
#430740000000
0!
0%
#430745000000
1!
1%
#430750000000
0!
0%
#430755000000
1!
1%
#430760000000
0!
0%
#430765000000
1!
1%
#430770000000
0!
0%
#430775000000
1!
1%
#430780000000
0!
0%
#430785000000
1!
1%
#430790000000
0!
0%
#430795000000
1!
1%
#430800000000
0!
0%
#430805000000
1!
1%
#430810000000
0!
0%
#430815000000
1!
1%
#430820000000
0!
0%
#430825000000
1!
1%
#430830000000
0!
0%
#430835000000
1!
1%
#430840000000
0!
0%
#430845000000
1!
1%
#430850000000
0!
0%
#430855000000
1!
1%
#430860000000
0!
0%
#430865000000
1!
1%
#430870000000
0!
0%
#430875000000
1!
1%
#430880000000
0!
0%
#430885000000
1!
1%
#430890000000
0!
0%
#430895000000
1!
1%
#430900000000
0!
0%
#430905000000
1!
1%
#430910000000
0!
0%
#430915000000
1!
1%
#430920000000
0!
0%
#430925000000
1!
1%
#430930000000
0!
0%
#430935000000
1!
1%
#430940000000
0!
0%
#430945000000
1!
1%
#430950000000
0!
0%
#430955000000
1!
1%
#430960000000
0!
0%
#430965000000
1!
1%
#430970000000
0!
0%
#430975000000
1!
1%
#430980000000
0!
0%
#430985000000
1!
1%
#430990000000
0!
0%
#430995000000
1!
1%
#431000000000
0!
0%
#431005000000
1!
1%
#431010000000
0!
0%
#431015000000
1!
1%
#431020000000
0!
0%
#431025000000
1!
1%
#431030000000
0!
0%
#431035000000
1!
1%
#431040000000
0!
0%
#431045000000
1!
1%
#431050000000
0!
0%
#431055000000
1!
1%
#431060000000
0!
0%
#431065000000
1!
1%
#431070000000
0!
0%
#431075000000
1!
1%
#431080000000
0!
0%
#431085000000
1!
1%
#431090000000
0!
0%
#431095000000
1!
1%
#431100000000
0!
0%
#431105000000
1!
1%
#431110000000
0!
0%
#431115000000
1!
1%
#431120000000
0!
0%
#431125000000
1!
1%
#431130000000
0!
0%
#431135000000
1!
1%
#431140000000
0!
0%
#431145000000
1!
1%
#431150000000
0!
0%
#431155000000
1!
1%
#431160000000
0!
0%
#431165000000
1!
1%
#431170000000
0!
0%
#431175000000
1!
1%
#431180000000
0!
0%
#431185000000
1!
1%
#431190000000
0!
0%
#431195000000
1!
1%
#431200000000
0!
0%
#431205000000
1!
1%
#431210000000
0!
0%
#431215000000
1!
1%
#431220000000
0!
0%
#431225000000
1!
1%
#431230000000
0!
0%
#431235000000
1!
1%
#431240000000
0!
0%
#431245000000
1!
1%
#431250000000
0!
0%
#431255000000
1!
1%
#431260000000
0!
0%
#431265000000
1!
1%
#431270000000
0!
0%
#431275000000
1!
1%
#431280000000
0!
0%
#431285000000
1!
1%
#431290000000
0!
0%
#431295000000
1!
1%
#431300000000
0!
0%
#431305000000
1!
1%
#431310000000
0!
0%
#431315000000
1!
1%
#431320000000
0!
0%
#431325000000
1!
1%
#431330000000
0!
0%
#431335000000
1!
1%
#431340000000
0!
0%
#431345000000
1!
1%
#431350000000
0!
0%
#431355000000
1!
1%
#431360000000
0!
0%
#431365000000
1!
1%
#431370000000
0!
0%
#431375000000
1!
1%
#431380000000
0!
0%
#431385000000
1!
1%
#431390000000
0!
0%
#431395000000
1!
1%
#431400000000
0!
0%
#431405000000
1!
1%
#431410000000
0!
0%
#431415000000
1!
1%
#431420000000
0!
0%
#431425000000
1!
1%
#431430000000
0!
0%
#431435000000
1!
1%
#431440000000
0!
0%
#431445000000
1!
1%
#431450000000
0!
0%
#431455000000
1!
1%
#431460000000
0!
0%
#431465000000
1!
1%
#431470000000
0!
0%
#431475000000
1!
1%
#431480000000
0!
0%
#431485000000
1!
1%
#431490000000
0!
0%
#431495000000
1!
1%
#431500000000
0!
0%
#431505000000
1!
1%
#431510000000
0!
0%
#431515000000
1!
1%
#431520000000
0!
0%
#431525000000
1!
1%
#431530000000
0!
0%
#431535000000
1!
1%
#431540000000
0!
0%
#431545000000
1!
1%
#431550000000
0!
0%
#431555000000
1!
1%
#431560000000
0!
0%
#431565000000
1!
1%
#431570000000
0!
0%
#431575000000
1!
1%
#431580000000
0!
0%
#431585000000
1!
1%
#431590000000
0!
0%
#431595000000
1!
1%
#431600000000
0!
0%
#431605000000
1!
1%
#431610000000
0!
0%
#431615000000
1!
1%
#431620000000
0!
0%
#431625000000
1!
1%
#431630000000
0!
0%
#431635000000
1!
1%
#431640000000
0!
0%
#431645000000
1!
1%
#431650000000
0!
0%
#431655000000
1!
1%
#431660000000
0!
0%
#431665000000
1!
1%
#431670000000
0!
0%
#431675000000
1!
1%
#431680000000
0!
0%
#431685000000
1!
1%
#431690000000
0!
0%
#431695000000
1!
1%
#431700000000
0!
0%
#431705000000
1!
1%
#431710000000
0!
0%
#431715000000
1!
1%
#431720000000
0!
0%
#431725000000
1!
1%
#431730000000
0!
0%
#431735000000
1!
1%
#431740000000
0!
0%
#431745000000
1!
1%
#431750000000
0!
0%
#431755000000
1!
1%
#431760000000
0!
0%
#431765000000
1!
1%
#431770000000
0!
0%
#431775000000
1!
1%
#431780000000
0!
0%
#431785000000
1!
1%
#431790000000
0!
0%
#431795000000
1!
1%
#431800000000
0!
0%
#431805000000
1!
1%
#431810000000
0!
0%
#431815000000
1!
1%
#431820000000
0!
0%
#431825000000
1!
1%
#431830000000
0!
0%
#431835000000
1!
1%
#431840000000
0!
0%
#431845000000
1!
1%
#431850000000
0!
0%
#431855000000
1!
1%
#431860000000
0!
0%
#431865000000
1!
1%
#431870000000
0!
0%
#431875000000
1!
1%
#431880000000
0!
0%
#431885000000
1!
1%
#431890000000
0!
0%
#431895000000
1!
1%
#431900000000
0!
0%
#431905000000
1!
1%
#431910000000
0!
0%
#431915000000
1!
1%
#431920000000
0!
0%
#431925000000
1!
1%
#431930000000
0!
0%
#431935000000
1!
1%
#431940000000
0!
0%
#431945000000
1!
1%
#431950000000
0!
0%
#431955000000
1!
1%
#431960000000
0!
0%
#431965000000
1!
1%
#431970000000
0!
0%
#431975000000
1!
1%
#431980000000
0!
0%
#431985000000
1!
1%
#431990000000
0!
0%
#431995000000
1!
1%
#432000000000
0!
0%
#432005000000
1!
1%
#432010000000
0!
0%
#432015000000
1!
1%
#432020000000
0!
0%
#432025000000
1!
1%
#432030000000
0!
0%
#432035000000
1!
1%
#432040000000
0!
0%
#432045000000
1!
1%
#432050000000
0!
0%
#432055000000
1!
1%
#432060000000
0!
0%
#432065000000
1!
1%
#432070000000
0!
0%
#432075000000
1!
1%
#432080000000
0!
0%
#432085000000
1!
1%
#432090000000
0!
0%
#432095000000
1!
1%
#432100000000
0!
0%
#432105000000
1!
1%
#432110000000
0!
0%
#432115000000
1!
1%
#432120000000
0!
0%
#432125000000
1!
1%
#432130000000
0!
0%
#432135000000
1!
1%
#432140000000
0!
0%
#432145000000
1!
1%
#432150000000
0!
0%
#432155000000
1!
1%
#432160000000
0!
0%
#432165000000
1!
1%
#432170000000
0!
0%
#432175000000
1!
1%
#432180000000
0!
0%
#432185000000
1!
1%
#432190000000
0!
0%
#432195000000
1!
1%
#432200000000
0!
0%
#432205000000
1!
1%
#432210000000
0!
0%
#432215000000
1!
1%
#432220000000
0!
0%
#432225000000
1!
1%
#432230000000
0!
0%
#432235000000
1!
1%
#432240000000
0!
0%
#432245000000
1!
1%
#432250000000
0!
0%
#432255000000
1!
1%
#432260000000
0!
0%
#432265000000
1!
1%
#432270000000
0!
0%
#432275000000
1!
1%
#432280000000
0!
0%
#432285000000
1!
1%
#432290000000
0!
0%
#432295000000
1!
1%
#432300000000
0!
0%
#432305000000
1!
1%
#432310000000
0!
0%
#432315000000
1!
1%
#432320000000
0!
0%
#432325000000
1!
1%
#432330000000
0!
0%
#432335000000
1!
1%
#432340000000
0!
0%
#432345000000
1!
1%
#432350000000
0!
0%
#432355000000
1!
1%
#432360000000
0!
0%
#432365000000
1!
1%
#432370000000
0!
0%
#432375000000
1!
1%
#432380000000
0!
0%
#432385000000
1!
1%
#432390000000
0!
0%
#432395000000
1!
1%
#432400000000
0!
0%
#432405000000
1!
1%
#432410000000
0!
0%
#432415000000
1!
1%
#432420000000
0!
0%
#432425000000
1!
1%
#432430000000
0!
0%
#432435000000
1!
1%
#432440000000
0!
0%
#432445000000
1!
1%
#432450000000
0!
0%
#432455000000
1!
1%
#432460000000
0!
0%
#432465000000
1!
1%
#432470000000
0!
0%
#432475000000
1!
1%
#432480000000
0!
0%
#432485000000
1!
1%
#432490000000
0!
0%
#432495000000
1!
1%
#432500000000
0!
0%
#432505000000
1!
1%
#432510000000
0!
0%
#432515000000
1!
1%
#432520000000
0!
0%
#432525000000
1!
1%
#432530000000
0!
0%
#432535000000
1!
1%
#432540000000
0!
0%
#432545000000
1!
1%
#432550000000
0!
0%
#432555000000
1!
1%
#432560000000
0!
0%
#432565000000
1!
1%
#432570000000
0!
0%
#432575000000
1!
1%
#432580000000
0!
0%
#432585000000
1!
1%
#432590000000
0!
0%
#432595000000
1!
1%
#432600000000
0!
0%
#432605000000
1!
1%
#432610000000
0!
0%
#432615000000
1!
1%
#432620000000
0!
0%
#432625000000
1!
1%
#432630000000
0!
0%
#432635000000
1!
1%
#432640000000
0!
0%
#432645000000
1!
1%
#432650000000
0!
0%
#432655000000
1!
1%
#432660000000
0!
0%
#432665000000
1!
1%
#432670000000
0!
0%
#432675000000
1!
1%
#432680000000
0!
0%
#432685000000
1!
1%
#432690000000
0!
0%
#432695000000
1!
1%
#432700000000
0!
0%
#432705000000
1!
1%
#432710000000
0!
0%
#432715000000
1!
1%
#432720000000
0!
0%
#432725000000
1!
1%
#432730000000
0!
0%
#432735000000
1!
1%
#432740000000
0!
0%
#432745000000
1!
1%
#432750000000
0!
0%
#432755000000
1!
1%
#432760000000
0!
0%
#432765000000
1!
1%
#432770000000
0!
0%
#432775000000
1!
1%
#432780000000
0!
0%
#432785000000
1!
1%
#432790000000
0!
0%
#432795000000
1!
1%
#432800000000
0!
0%
#432805000000
1!
1%
#432810000000
0!
0%
#432815000000
1!
1%
#432820000000
0!
0%
#432825000000
1!
1%
#432830000000
0!
0%
#432835000000
1!
1%
#432840000000
0!
0%
#432845000000
1!
1%
#432850000000
0!
0%
#432855000000
1!
1%
#432860000000
0!
0%
#432865000000
1!
1%
#432870000000
0!
0%
#432875000000
1!
1%
#432880000000
0!
0%
#432885000000
1!
1%
#432890000000
0!
0%
#432895000000
1!
1%
#432900000000
0!
0%
#432905000000
1!
1%
#432910000000
0!
0%
#432915000000
1!
1%
#432920000000
0!
0%
#432925000000
1!
1%
#432930000000
0!
0%
#432935000000
1!
1%
#432940000000
0!
0%
#432945000000
1!
1%
#432950000000
0!
0%
#432955000000
1!
1%
#432960000000
0!
0%
#432965000000
1!
1%
#432970000000
0!
0%
#432975000000
1!
1%
#432980000000
0!
0%
#432985000000
1!
1%
#432990000000
0!
0%
#432995000000
1!
1%
#433000000000
0!
0%
#433005000000
1!
1%
#433010000000
0!
0%
#433015000000
1!
1%
#433020000000
0!
0%
#433025000000
1!
1%
#433030000000
0!
0%
#433035000000
1!
1%
#433040000000
0!
0%
#433045000000
1!
1%
#433050000000
0!
0%
#433055000000
1!
1%
#433060000000
0!
0%
#433065000000
1!
1%
#433070000000
0!
0%
#433075000000
1!
1%
#433080000000
0!
0%
#433085000000
1!
1%
#433090000000
0!
0%
#433095000000
1!
1%
#433100000000
0!
0%
#433105000000
1!
1%
#433110000000
0!
0%
#433115000000
1!
1%
#433120000000
0!
0%
#433125000000
1!
1%
#433130000000
0!
0%
#433135000000
1!
1%
#433140000000
0!
0%
#433145000000
1!
1%
#433150000000
0!
0%
#433155000000
1!
1%
#433160000000
0!
0%
#433165000000
1!
1%
#433170000000
0!
0%
#433175000000
1!
1%
#433180000000
0!
0%
#433185000000
1!
1%
#433190000000
0!
0%
#433195000000
1!
1%
#433200000000
0!
0%
#433205000000
1!
1%
#433210000000
0!
0%
#433215000000
1!
1%
#433220000000
0!
0%
#433225000000
1!
1%
#433230000000
0!
0%
#433235000000
1!
1%
#433240000000
0!
0%
#433245000000
1!
1%
#433250000000
0!
0%
#433255000000
1!
1%
#433260000000
0!
0%
#433265000000
1!
1%
#433270000000
0!
0%
#433275000000
1!
1%
#433280000000
0!
0%
#433285000000
1!
1%
#433290000000
0!
0%
#433295000000
1!
1%
#433300000000
0!
0%
#433305000000
1!
1%
#433310000000
0!
0%
#433315000000
1!
1%
#433320000000
0!
0%
#433325000000
1!
1%
#433330000000
0!
0%
#433335000000
1!
1%
#433340000000
0!
0%
#433345000000
1!
1%
#433350000000
0!
0%
#433355000000
1!
1%
#433360000000
0!
0%
#433365000000
1!
1%
#433370000000
0!
0%
#433375000000
1!
1%
#433380000000
0!
0%
#433385000000
1!
1%
#433390000000
0!
0%
#433395000000
1!
1%
#433400000000
0!
0%
#433405000000
1!
1%
#433410000000
0!
0%
#433415000000
1!
1%
#433420000000
0!
0%
#433425000000
1!
1%
#433430000000
0!
0%
#433435000000
1!
1%
#433440000000
0!
0%
#433445000000
1!
1%
#433450000000
0!
0%
#433455000000
1!
1%
#433460000000
0!
0%
#433465000000
1!
1%
#433470000000
0!
0%
#433475000000
1!
1%
#433480000000
0!
0%
#433485000000
1!
1%
#433490000000
0!
0%
#433495000000
1!
1%
#433500000000
0!
0%
#433505000000
1!
1%
#433510000000
0!
0%
#433515000000
1!
1%
#433520000000
0!
0%
#433525000000
1!
1%
#433530000000
0!
0%
#433535000000
1!
1%
#433540000000
0!
0%
#433545000000
1!
1%
#433550000000
0!
0%
#433555000000
1!
1%
#433560000000
0!
0%
#433565000000
1!
1%
#433570000000
0!
0%
#433575000000
1!
1%
#433580000000
0!
0%
#433585000000
1!
1%
#433590000000
0!
0%
#433595000000
1!
1%
#433600000000
0!
0%
#433605000000
1!
1%
#433610000000
0!
0%
#433615000000
1!
1%
#433620000000
0!
0%
#433625000000
1!
1%
#433630000000
0!
0%
#433635000000
1!
1%
#433640000000
0!
0%
#433645000000
1!
1%
#433650000000
0!
0%
#433655000000
1!
1%
#433660000000
0!
0%
#433665000000
1!
1%
#433670000000
0!
0%
#433675000000
1!
1%
#433680000000
0!
0%
#433685000000
1!
1%
#433690000000
0!
0%
#433695000000
1!
1%
#433700000000
0!
0%
#433705000000
1!
1%
#433710000000
0!
0%
#433715000000
1!
1%
#433720000000
0!
0%
#433725000000
1!
1%
#433730000000
0!
0%
#433735000000
1!
1%
#433740000000
0!
0%
#433745000000
1!
1%
#433750000000
0!
0%
#433755000000
1!
1%
#433760000000
0!
0%
#433765000000
1!
1%
#433770000000
0!
0%
#433775000000
1!
1%
#433780000000
0!
0%
#433785000000
1!
1%
#433790000000
0!
0%
#433795000000
1!
1%
#433800000000
0!
0%
#433805000000
1!
1%
#433810000000
0!
0%
#433815000000
1!
1%
#433820000000
0!
0%
#433825000000
1!
1%
#433830000000
0!
0%
#433835000000
1!
1%
#433840000000
0!
0%
#433845000000
1!
1%
#433850000000
0!
0%
#433855000000
1!
1%
#433860000000
0!
0%
#433865000000
1!
1%
#433870000000
0!
0%
#433875000000
1!
1%
#433880000000
0!
0%
#433885000000
1!
1%
#433890000000
0!
0%
#433895000000
1!
1%
#433900000000
0!
0%
#433905000000
1!
1%
#433910000000
0!
0%
#433915000000
1!
1%
#433920000000
0!
0%
#433925000000
1!
1%
#433930000000
0!
0%
#433935000000
1!
1%
#433940000000
0!
0%
#433945000000
1!
1%
#433950000000
0!
0%
#433955000000
1!
1%
#433960000000
0!
0%
#433965000000
1!
1%
#433970000000
0!
0%
#433975000000
1!
1%
#433980000000
0!
0%
#433985000000
1!
1%
#433990000000
0!
0%
#433995000000
1!
1%
#434000000000
0!
0%
#434005000000
1!
1%
#434010000000
0!
0%
#434015000000
1!
1%
#434020000000
0!
0%
#434025000000
1!
1%
#434030000000
0!
0%
#434035000000
1!
1%
#434040000000
0!
0%
#434045000000
1!
1%
#434050000000
0!
0%
#434055000000
1!
1%
#434060000000
0!
0%
#434065000000
1!
1%
#434070000000
0!
0%
#434075000000
1!
1%
#434080000000
0!
0%
#434085000000
1!
1%
#434090000000
0!
0%
#434095000000
1!
1%
#434100000000
0!
0%
#434105000000
1!
1%
#434110000000
0!
0%
#434115000000
1!
1%
#434120000000
0!
0%
#434125000000
1!
1%
#434130000000
0!
0%
#434135000000
1!
1%
#434140000000
0!
0%
#434145000000
1!
1%
#434150000000
0!
0%
#434155000000
1!
1%
#434160000000
0!
0%
#434165000000
1!
1%
#434170000000
0!
0%
#434175000000
1!
1%
#434180000000
0!
0%
#434185000000
1!
1%
#434190000000
0!
0%
#434195000000
1!
1%
#434200000000
0!
0%
#434205000000
1!
1%
#434210000000
0!
0%
#434215000000
1!
1%
#434220000000
0!
0%
#434225000000
1!
1%
#434230000000
0!
0%
#434235000000
1!
1%
#434240000000
0!
0%
#434245000000
1!
1%
#434250000000
0!
0%
#434255000000
1!
1%
#434260000000
0!
0%
#434265000000
1!
1%
#434270000000
0!
0%
#434275000000
1!
1%
#434280000000
0!
0%
#434285000000
1!
1%
#434290000000
0!
0%
#434295000000
1!
1%
#434300000000
0!
0%
#434305000000
1!
1%
#434310000000
0!
0%
#434315000000
1!
1%
#434320000000
0!
0%
#434325000000
1!
1%
#434330000000
0!
0%
#434335000000
1!
1%
#434340000000
0!
0%
#434345000000
1!
1%
#434350000000
0!
0%
#434355000000
1!
1%
#434360000000
0!
0%
#434365000000
1!
1%
#434370000000
0!
0%
#434375000000
1!
1%
#434380000000
0!
0%
#434385000000
1!
1%
#434390000000
0!
0%
#434395000000
1!
1%
#434400000000
0!
0%
#434405000000
1!
1%
#434410000000
0!
0%
#434415000000
1!
1%
#434420000000
0!
0%
#434425000000
1!
1%
#434430000000
0!
0%
#434435000000
1!
1%
#434440000000
0!
0%
#434445000000
1!
1%
#434450000000
0!
0%
#434455000000
1!
1%
#434460000000
0!
0%
#434465000000
1!
1%
#434470000000
0!
0%
#434475000000
1!
1%
#434480000000
0!
0%
#434485000000
1!
1%
#434490000000
0!
0%
#434495000000
1!
1%
#434500000000
0!
0%
#434505000000
1!
1%
#434510000000
0!
0%
#434515000000
1!
1%
#434520000000
0!
0%
#434525000000
1!
1%
#434530000000
0!
0%
#434535000000
1!
1%
#434540000000
0!
0%
#434545000000
1!
1%
#434550000000
0!
0%
#434555000000
1!
1%
#434560000000
0!
0%
#434565000000
1!
1%
#434570000000
0!
0%
#434575000000
1!
1%
#434580000000
0!
0%
#434585000000
1!
1%
#434590000000
0!
0%
#434595000000
1!
1%
#434600000000
0!
0%
#434605000000
1!
1%
#434610000000
0!
0%
#434615000000
1!
1%
#434620000000
0!
0%
#434625000000
1!
1%
#434630000000
0!
0%
#434635000000
1!
1%
#434640000000
0!
0%
#434645000000
1!
1%
#434650000000
0!
0%
#434655000000
1!
1%
#434660000000
0!
0%
#434665000000
1!
1%
#434670000000
0!
0%
#434675000000
1!
1%
#434680000000
0!
0%
#434685000000
1!
1%
#434690000000
0!
0%
#434695000000
1!
1%
#434700000000
0!
0%
#434705000000
1!
1%
#434710000000
0!
0%
#434715000000
1!
1%
#434720000000
0!
0%
#434725000000
1!
1%
#434730000000
0!
0%
#434735000000
1!
1%
#434740000000
0!
0%
#434745000000
1!
1%
#434750000000
0!
0%
#434755000000
1!
1%
#434760000000
0!
0%
#434765000000
1!
1%
#434770000000
0!
0%
#434775000000
1!
1%
#434780000000
0!
0%
#434785000000
1!
1%
#434790000000
0!
0%
#434795000000
1!
1%
#434800000000
0!
0%
#434805000000
1!
1%
#434810000000
0!
0%
#434815000000
1!
1%
#434820000000
0!
0%
#434825000000
1!
1%
#434830000000
0!
0%
#434835000000
1!
1%
#434840000000
0!
0%
#434845000000
1!
1%
#434850000000
0!
0%
#434855000000
1!
1%
#434860000000
0!
0%
#434865000000
1!
1%
#434870000000
0!
0%
#434875000000
1!
1%
#434880000000
0!
0%
#434885000000
1!
1%
#434890000000
0!
0%
#434895000000
1!
1%
#434900000000
0!
0%
#434905000000
1!
1%
#434910000000
0!
0%
#434915000000
1!
1%
#434920000000
0!
0%
#434925000000
1!
1%
#434930000000
0!
0%
#434935000000
1!
1%
#434940000000
0!
0%
#434945000000
1!
1%
#434950000000
0!
0%
#434955000000
1!
1%
#434960000000
0!
0%
#434965000000
1!
1%
#434970000000
0!
0%
#434975000000
1!
1%
#434980000000
0!
0%
#434985000000
1!
1%
#434990000000
0!
0%
#434995000000
1!
1%
#435000000000
0!
0%
#435005000000
1!
1%
#435010000000
0!
0%
#435015000000
1!
1%
#435020000000
0!
0%
#435025000000
1!
1%
#435030000000
0!
0%
#435035000000
1!
1%
#435040000000
0!
0%
#435045000000
1!
1%
#435050000000
0!
0%
#435055000000
1!
1%
#435060000000
0!
0%
#435065000000
1!
1%
#435070000000
0!
0%
#435075000000
1!
1%
#435080000000
0!
0%
#435085000000
1!
1%
#435090000000
0!
0%
#435095000000
1!
1%
#435100000000
0!
0%
#435105000000
1!
1%
#435110000000
0!
0%
#435115000000
1!
1%
#435120000000
0!
0%
#435125000000
1!
1%
#435130000000
0!
0%
#435135000000
1!
1%
#435140000000
0!
0%
#435145000000
1!
1%
#435150000000
0!
0%
#435155000000
1!
1%
#435160000000
0!
0%
#435165000000
1!
1%
#435170000000
0!
0%
#435175000000
1!
1%
#435180000000
0!
0%
#435185000000
1!
1%
#435190000000
0!
0%
#435195000000
1!
1%
#435200000000
0!
0%
#435205000000
1!
1%
#435210000000
0!
0%
#435215000000
1!
1%
#435220000000
0!
0%
#435225000000
1!
1%
#435230000000
0!
0%
#435235000000
1!
1%
#435240000000
0!
0%
#435245000000
1!
1%
#435250000000
0!
0%
#435255000000
1!
1%
#435260000000
0!
0%
#435265000000
1!
1%
#435270000000
0!
0%
#435275000000
1!
1%
#435280000000
0!
0%
#435285000000
1!
1%
#435290000000
0!
0%
#435295000000
1!
1%
#435300000000
0!
0%
#435305000000
1!
1%
#435310000000
0!
0%
#435315000000
1!
1%
#435320000000
0!
0%
#435325000000
1!
1%
#435330000000
0!
0%
#435335000000
1!
1%
#435340000000
0!
0%
#435345000000
1!
1%
#435350000000
0!
0%
#435355000000
1!
1%
#435360000000
0!
0%
#435365000000
1!
1%
#435370000000
0!
0%
#435375000000
1!
1%
#435380000000
0!
0%
#435385000000
1!
1%
#435390000000
0!
0%
#435395000000
1!
1%
#435400000000
0!
0%
#435405000000
1!
1%
#435410000000
0!
0%
#435415000000
1!
1%
#435420000000
0!
0%
#435425000000
1!
1%
#435430000000
0!
0%
#435435000000
1!
1%
#435440000000
0!
0%
#435445000000
1!
1%
#435450000000
0!
0%
#435455000000
1!
1%
#435460000000
0!
0%
#435465000000
1!
1%
#435470000000
0!
0%
#435475000000
1!
1%
#435480000000
0!
0%
#435485000000
1!
1%
#435490000000
0!
0%
#435495000000
1!
1%
#435500000000
0!
0%
#435505000000
1!
1%
#435510000000
0!
0%
#435515000000
1!
1%
#435520000000
0!
0%
#435525000000
1!
1%
#435530000000
0!
0%
#435535000000
1!
1%
#435540000000
0!
0%
#435545000000
1!
1%
#435550000000
0!
0%
#435555000000
1!
1%
#435560000000
0!
0%
#435565000000
1!
1%
#435570000000
0!
0%
#435575000000
1!
1%
#435580000000
0!
0%
#435585000000
1!
1%
#435590000000
0!
0%
#435595000000
1!
1%
#435600000000
0!
0%
#435605000000
1!
1%
#435610000000
0!
0%
#435615000000
1!
1%
#435620000000
0!
0%
#435625000000
1!
1%
#435630000000
0!
0%
#435635000000
1!
1%
#435640000000
0!
0%
#435645000000
1!
1%
#435650000000
0!
0%
#435655000000
1!
1%
#435660000000
0!
0%
#435665000000
1!
1%
#435670000000
0!
0%
#435675000000
1!
1%
#435680000000
0!
0%
#435685000000
1!
1%
#435690000000
0!
0%
#435695000000
1!
1%
#435700000000
0!
0%
#435705000000
1!
1%
#435710000000
0!
0%
#435715000000
1!
1%
#435720000000
0!
0%
#435725000000
1!
1%
#435730000000
0!
0%
#435735000000
1!
1%
#435740000000
0!
0%
#435745000000
1!
1%
#435750000000
0!
0%
#435755000000
1!
1%
#435760000000
0!
0%
#435765000000
1!
1%
#435770000000
0!
0%
#435775000000
1!
1%
#435780000000
0!
0%
#435785000000
1!
1%
#435790000000
0!
0%
#435795000000
1!
1%
#435800000000
0!
0%
#435805000000
1!
1%
#435810000000
0!
0%
#435815000000
1!
1%
#435820000000
0!
0%
#435825000000
1!
1%
#435830000000
0!
0%
#435835000000
1!
1%
#435840000000
0!
0%
#435845000000
1!
1%
#435850000000
0!
0%
#435855000000
1!
1%
#435860000000
0!
0%
#435865000000
1!
1%
#435870000000
0!
0%
#435875000000
1!
1%
#435880000000
0!
0%
#435885000000
1!
1%
#435890000000
0!
0%
#435895000000
1!
1%
#435900000000
0!
0%
#435905000000
1!
1%
#435910000000
0!
0%
#435915000000
1!
1%
#435920000000
0!
0%
#435925000000
1!
1%
#435930000000
0!
0%
#435935000000
1!
1%
#435940000000
0!
0%
#435945000000
1!
1%
#435950000000
0!
0%
#435955000000
1!
1%
#435960000000
0!
0%
#435965000000
1!
1%
#435970000000
0!
0%
#435975000000
1!
1%
#435980000000
0!
0%
#435985000000
1!
1%
#435990000000
0!
0%
#435995000000
1!
1%
#436000000000
0!
0%
#436005000000
1!
1%
#436010000000
0!
0%
#436015000000
1!
1%
#436020000000
0!
0%
#436025000000
1!
1%
#436030000000
0!
0%
#436035000000
1!
1%
#436040000000
0!
0%
#436045000000
1!
1%
#436050000000
0!
0%
#436055000000
1!
1%
#436060000000
0!
0%
#436065000000
1!
1%
#436070000000
0!
0%
#436075000000
1!
1%
#436080000000
0!
0%
#436085000000
1!
1%
#436090000000
0!
0%
#436095000000
1!
1%
#436100000000
0!
0%
#436105000000
1!
1%
#436110000000
0!
0%
#436115000000
1!
1%
#436120000000
0!
0%
#436125000000
1!
1%
#436130000000
0!
0%
#436135000000
1!
1%
#436140000000
0!
0%
#436145000000
1!
1%
#436150000000
0!
0%
#436155000000
1!
1%
#436160000000
0!
0%
#436165000000
1!
1%
#436170000000
0!
0%
#436175000000
1!
1%
#436180000000
0!
0%
#436185000000
1!
1%
#436190000000
0!
0%
#436195000000
1!
1%
#436200000000
0!
0%
#436205000000
1!
1%
#436210000000
0!
0%
#436215000000
1!
1%
#436220000000
0!
0%
#436225000000
1!
1%
#436230000000
0!
0%
#436235000000
1!
1%
#436240000000
0!
0%
#436245000000
1!
1%
#436250000000
0!
0%
#436255000000
1!
1%
#436260000000
0!
0%
#436265000000
1!
1%
#436270000000
0!
0%
#436275000000
1!
1%
#436280000000
0!
0%
#436285000000
1!
1%
#436290000000
0!
0%
#436295000000
1!
1%
#436300000000
0!
0%
#436305000000
1!
1%
#436310000000
0!
0%
#436315000000
1!
1%
#436320000000
0!
0%
#436325000000
1!
1%
#436330000000
0!
0%
#436335000000
1!
1%
#436340000000
0!
0%
#436345000000
1!
1%
#436350000000
0!
0%
#436355000000
1!
1%
#436360000000
0!
0%
#436365000000
1!
1%
#436370000000
0!
0%
#436375000000
1!
1%
#436380000000
0!
0%
#436385000000
1!
1%
#436390000000
0!
0%
#436395000000
1!
1%
#436400000000
0!
0%
#436405000000
1!
1%
#436410000000
0!
0%
#436415000000
1!
1%
#436420000000
0!
0%
#436425000000
1!
1%
#436430000000
0!
0%
#436435000000
1!
1%
#436440000000
0!
0%
#436445000000
1!
1%
#436450000000
0!
0%
#436455000000
1!
1%
#436460000000
0!
0%
#436465000000
1!
1%
#436470000000
0!
0%
#436475000000
1!
1%
#436480000000
0!
0%
#436485000000
1!
1%
#436490000000
0!
0%
#436495000000
1!
1%
#436500000000
0!
0%
#436505000000
1!
1%
#436510000000
0!
0%
#436515000000
1!
1%
#436520000000
0!
0%
#436525000000
1!
1%
#436530000000
0!
0%
#436535000000
1!
1%
#436540000000
0!
0%
#436545000000
1!
1%
#436550000000
0!
0%
#436555000000
1!
1%
#436560000000
0!
0%
#436565000000
1!
1%
#436570000000
0!
0%
#436575000000
1!
1%
#436580000000
0!
0%
#436585000000
1!
1%
#436590000000
0!
0%
#436595000000
1!
1%
#436600000000
0!
0%
#436605000000
1!
1%
#436610000000
0!
0%
#436615000000
1!
1%
#436620000000
0!
0%
#436625000000
1!
1%
#436630000000
0!
0%
#436635000000
1!
1%
#436640000000
0!
0%
#436645000000
1!
1%
#436650000000
0!
0%
#436655000000
1!
1%
#436660000000
0!
0%
#436665000000
1!
1%
#436670000000
0!
0%
#436675000000
1!
1%
#436680000000
0!
0%
#436685000000
1!
1%
#436690000000
0!
0%
#436695000000
1!
1%
#436700000000
0!
0%
#436705000000
1!
1%
#436710000000
0!
0%
#436715000000
1!
1%
#436720000000
0!
0%
#436725000000
1!
1%
#436730000000
0!
0%
#436735000000
1!
1%
#436740000000
0!
0%
#436745000000
1!
1%
#436750000000
0!
0%
#436755000000
1!
1%
#436760000000
0!
0%
#436765000000
1!
1%
#436770000000
0!
0%
#436775000000
1!
1%
#436780000000
0!
0%
#436785000000
1!
1%
#436790000000
0!
0%
#436795000000
1!
1%
#436800000000
0!
0%
#436805000000
1!
1%
#436810000000
0!
0%
#436815000000
1!
1%
#436820000000
0!
0%
#436825000000
1!
1%
#436830000000
0!
0%
#436835000000
1!
1%
#436840000000
0!
0%
#436845000000
1!
1%
#436850000000
0!
0%
#436855000000
1!
1%
#436860000000
0!
0%
#436865000000
1!
1%
#436870000000
0!
0%
#436875000000
1!
1%
#436880000000
0!
0%
#436885000000
1!
1%
#436890000000
0!
0%
#436895000000
1!
1%
#436900000000
0!
0%
#436905000000
1!
1%
#436910000000
0!
0%
#436915000000
1!
1%
#436920000000
0!
0%
#436925000000
1!
1%
#436930000000
0!
0%
#436935000000
1!
1%
#436940000000
0!
0%
#436945000000
1!
1%
#436950000000
0!
0%
#436955000000
1!
1%
#436960000000
0!
0%
#436965000000
1!
1%
#436970000000
0!
0%
#436975000000
1!
1%
#436980000000
0!
0%
#436985000000
1!
1%
#436990000000
0!
0%
#436995000000
1!
1%
#437000000000
0!
0%
#437005000000
1!
1%
#437010000000
0!
0%
#437015000000
1!
1%
#437020000000
0!
0%
#437025000000
1!
1%
#437030000000
0!
0%
#437035000000
1!
1%
#437040000000
0!
0%
#437045000000
1!
1%
#437050000000
0!
0%
#437055000000
1!
1%
#437060000000
0!
0%
#437065000000
1!
1%
#437070000000
0!
0%
#437075000000
1!
1%
#437080000000
0!
0%
#437085000000
1!
1%
#437090000000
0!
0%
#437095000000
1!
1%
#437100000000
0!
0%
#437105000000
1!
1%
#437110000000
0!
0%
#437115000000
1!
1%
#437120000000
0!
0%
#437125000000
1!
1%
#437130000000
0!
0%
#437135000000
1!
1%
#437140000000
0!
0%
#437145000000
1!
1%
#437150000000
0!
0%
#437155000000
1!
1%
#437160000000
0!
0%
#437165000000
1!
1%
#437170000000
0!
0%
#437175000000
1!
1%
#437180000000
0!
0%
#437185000000
1!
1%
#437190000000
0!
0%
#437195000000
1!
1%
#437200000000
0!
0%
#437205000000
1!
1%
#437210000000
0!
0%
#437215000000
1!
1%
#437220000000
0!
0%
#437225000000
1!
1%
#437230000000
0!
0%
#437235000000
1!
1%
#437240000000
0!
0%
#437245000000
1!
1%
#437250000000
0!
0%
#437255000000
1!
1%
#437260000000
0!
0%
#437265000000
1!
1%
#437270000000
0!
0%
#437275000000
1!
1%
#437280000000
0!
0%
#437285000000
1!
1%
#437290000000
0!
0%
#437295000000
1!
1%
#437300000000
0!
0%
#437305000000
1!
1%
#437310000000
0!
0%
#437315000000
1!
1%
#437320000000
0!
0%
#437325000000
1!
1%
#437330000000
0!
0%
#437335000000
1!
1%
#437340000000
0!
0%
#437345000000
1!
1%
#437350000000
0!
0%
#437355000000
1!
1%
#437360000000
0!
0%
#437365000000
1!
1%
#437370000000
0!
0%
#437375000000
1!
1%
#437380000000
0!
0%
#437385000000
1!
1%
#437390000000
0!
0%
#437395000000
1!
1%
#437400000000
0!
0%
#437405000000
1!
1%
#437410000000
0!
0%
#437415000000
1!
1%
#437420000000
0!
0%
#437425000000
1!
1%
#437430000000
0!
0%
#437435000000
1!
1%
#437440000000
0!
0%
#437445000000
1!
1%
#437450000000
0!
0%
#437455000000
1!
1%
#437460000000
0!
0%
#437465000000
1!
1%
#437470000000
0!
0%
#437475000000
1!
1%
#437480000000
0!
0%
#437485000000
1!
1%
#437490000000
0!
0%
#437495000000
1!
1%
#437500000000
0!
0%
#437505000000
1!
1%
#437510000000
0!
0%
#437515000000
1!
1%
#437520000000
0!
0%
#437525000000
1!
1%
#437530000000
0!
0%
#437535000000
1!
1%
#437540000000
0!
0%
#437545000000
1!
1%
#437550000000
0!
0%
#437555000000
1!
1%
#437560000000
0!
0%
#437565000000
1!
1%
#437570000000
0!
0%
#437575000000
1!
1%
#437580000000
0!
0%
#437585000000
1!
1%
#437590000000
0!
0%
#437595000000
1!
1%
#437600000000
0!
0%
#437605000000
1!
1%
#437610000000
0!
0%
#437615000000
1!
1%
#437620000000
0!
0%
#437625000000
1!
1%
#437630000000
0!
0%
#437635000000
1!
1%
#437640000000
0!
0%
#437645000000
1!
1%
#437650000000
0!
0%
#437655000000
1!
1%
#437660000000
0!
0%
#437665000000
1!
1%
#437670000000
0!
0%
#437675000000
1!
1%
#437680000000
0!
0%
#437685000000
1!
1%
#437690000000
0!
0%
#437695000000
1!
1%
#437700000000
0!
0%
#437705000000
1!
1%
#437710000000
0!
0%
#437715000000
1!
1%
#437720000000
0!
0%
#437725000000
1!
1%
#437730000000
0!
0%
#437735000000
1!
1%
#437740000000
0!
0%
#437745000000
1!
1%
#437750000000
0!
0%
#437755000000
1!
1%
#437760000000
0!
0%
#437765000000
1!
1%
#437770000000
0!
0%
#437775000000
1!
1%
#437780000000
0!
0%
#437785000000
1!
1%
#437790000000
0!
0%
#437795000000
1!
1%
#437800000000
0!
0%
#437805000000
1!
1%
#437810000000
0!
0%
#437815000000
1!
1%
#437820000000
0!
0%
#437825000000
1!
1%
#437830000000
0!
0%
#437835000000
1!
1%
#437840000000
0!
0%
#437845000000
1!
1%
#437850000000
0!
0%
#437855000000
1!
1%
#437860000000
0!
0%
#437865000000
1!
1%
#437870000000
0!
0%
#437875000000
1!
1%
#437880000000
0!
0%
#437885000000
1!
1%
#437890000000
0!
0%
#437895000000
1!
1%
#437900000000
0!
0%
#437905000000
1!
1%
#437910000000
0!
0%
#437915000000
1!
1%
#437920000000
0!
0%
#437925000000
1!
1%
#437930000000
0!
0%
#437935000000
1!
1%
#437940000000
0!
0%
#437945000000
1!
1%
#437950000000
0!
0%
#437955000000
1!
1%
#437960000000
0!
0%
#437965000000
1!
1%
#437970000000
0!
0%
#437975000000
1!
1%
#437980000000
0!
0%
#437985000000
1!
1%
#437990000000
0!
0%
#437995000000
1!
1%
#438000000000
0!
0%
#438005000000
1!
1%
#438010000000
0!
0%
#438015000000
1!
1%
#438020000000
0!
0%
#438025000000
1!
1%
#438030000000
0!
0%
#438035000000
1!
1%
#438040000000
0!
0%
#438045000000
1!
1%
#438050000000
0!
0%
#438055000000
1!
1%
#438060000000
0!
0%
#438065000000
1!
1%
#438070000000
0!
0%
#438075000000
1!
1%
#438080000000
0!
0%
#438085000000
1!
1%
#438090000000
0!
0%
#438095000000
1!
1%
#438100000000
0!
0%
#438105000000
1!
1%
#438110000000
0!
0%
#438115000000
1!
1%
#438120000000
0!
0%
#438125000000
1!
1%
#438130000000
0!
0%
#438135000000
1!
1%
#438140000000
0!
0%
#438145000000
1!
1%
#438150000000
0!
0%
#438155000000
1!
1%
#438160000000
0!
0%
#438165000000
1!
1%
#438170000000
0!
0%
#438175000000
1!
1%
#438180000000
0!
0%
#438185000000
1!
1%
#438190000000
0!
0%
#438195000000
1!
1%
#438200000000
0!
0%
#438205000000
1!
1%
#438210000000
0!
0%
#438215000000
1!
1%
#438220000000
0!
0%
#438225000000
1!
1%
#438230000000
0!
0%
#438235000000
1!
1%
#438240000000
0!
0%
#438245000000
1!
1%
#438250000000
0!
0%
#438255000000
1!
1%
#438260000000
0!
0%
#438265000000
1!
1%
#438270000000
0!
0%
#438275000000
1!
1%
#438280000000
0!
0%
#438285000000
1!
1%
#438290000000
0!
0%
#438295000000
1!
1%
#438300000000
0!
0%
#438305000000
1!
1%
#438310000000
0!
0%
#438315000000
1!
1%
#438320000000
0!
0%
#438325000000
1!
1%
#438330000000
0!
0%
#438335000000
1!
1%
#438340000000
0!
0%
#438345000000
1!
1%
#438350000000
0!
0%
#438355000000
1!
1%
#438360000000
0!
0%
#438365000000
1!
1%
#438370000000
0!
0%
#438375000000
1!
1%
#438380000000
0!
0%
#438385000000
1!
1%
#438390000000
0!
0%
#438395000000
1!
1%
#438400000000
0!
0%
#438405000000
1!
1%
#438410000000
0!
0%
#438415000000
1!
1%
#438420000000
0!
0%
#438425000000
1!
1%
#438430000000
0!
0%
#438435000000
1!
1%
#438440000000
0!
0%
#438445000000
1!
1%
#438450000000
0!
0%
#438455000000
1!
1%
#438460000000
0!
0%
#438465000000
1!
1%
#438470000000
0!
0%
#438475000000
1!
1%
#438480000000
0!
0%
#438485000000
1!
1%
#438490000000
0!
0%
#438495000000
1!
1%
#438500000000
0!
0%
#438505000000
1!
1%
#438510000000
0!
0%
#438515000000
1!
1%
#438520000000
0!
0%
#438525000000
1!
1%
#438530000000
0!
0%
#438535000000
1!
1%
#438540000000
0!
0%
#438545000000
1!
1%
#438550000000
0!
0%
#438555000000
1!
1%
#438560000000
0!
0%
#438565000000
1!
1%
#438570000000
0!
0%
#438575000000
1!
1%
#438580000000
0!
0%
#438585000000
1!
1%
#438590000000
0!
0%
#438595000000
1!
1%
#438600000000
0!
0%
#438605000000
1!
1%
#438610000000
0!
0%
#438615000000
1!
1%
#438620000000
0!
0%
#438625000000
1!
1%
#438630000000
0!
0%
#438635000000
1!
1%
#438640000000
0!
0%
#438645000000
1!
1%
#438650000000
0!
0%
#438655000000
1!
1%
#438660000000
0!
0%
#438665000000
1!
1%
#438670000000
0!
0%
#438675000000
1!
1%
#438680000000
0!
0%
#438685000000
1!
1%
#438690000000
0!
0%
#438695000000
1!
1%
#438700000000
0!
0%
#438705000000
1!
1%
#438710000000
0!
0%
#438715000000
1!
1%
#438720000000
0!
0%
#438725000000
1!
1%
#438730000000
0!
0%
#438735000000
1!
1%
#438740000000
0!
0%
#438745000000
1!
1%
#438750000000
0!
0%
#438755000000
1!
1%
#438760000000
0!
0%
#438765000000
1!
1%
#438770000000
0!
0%
#438775000000
1!
1%
#438780000000
0!
0%
#438785000000
1!
1%
#438790000000
0!
0%
#438795000000
1!
1%
#438800000000
0!
0%
#438805000000
1!
1%
#438810000000
0!
0%
#438815000000
1!
1%
#438820000000
0!
0%
#438825000000
1!
1%
#438830000000
0!
0%
#438835000000
1!
1%
#438840000000
0!
0%
#438845000000
1!
1%
#438850000000
0!
0%
#438855000000
1!
1%
#438860000000
0!
0%
#438865000000
1!
1%
#438870000000
0!
0%
#438875000000
1!
1%
#438880000000
0!
0%
#438885000000
1!
1%
#438890000000
0!
0%
#438895000000
1!
1%
#438900000000
0!
0%
#438905000000
1!
1%
#438910000000
0!
0%
#438915000000
1!
1%
#438920000000
0!
0%
#438925000000
1!
1%
#438930000000
0!
0%
#438935000000
1!
1%
#438940000000
0!
0%
#438945000000
1!
1%
#438950000000
0!
0%
#438955000000
1!
1%
#438960000000
0!
0%
#438965000000
1!
1%
#438970000000
0!
0%
#438975000000
1!
1%
#438980000000
0!
0%
#438985000000
1!
1%
#438990000000
0!
0%
#438995000000
1!
1%
#439000000000
0!
0%
#439005000000
1!
1%
#439010000000
0!
0%
#439015000000
1!
1%
#439020000000
0!
0%
#439025000000
1!
1%
#439030000000
0!
0%
#439035000000
1!
1%
#439040000000
0!
0%
#439045000000
1!
1%
#439050000000
0!
0%
#439055000000
1!
1%
#439060000000
0!
0%
#439065000000
1!
1%
#439070000000
0!
0%
#439075000000
1!
1%
#439080000000
0!
0%
#439085000000
1!
1%
#439090000000
0!
0%
#439095000000
1!
1%
#439100000000
0!
0%
#439105000000
1!
1%
#439110000000
0!
0%
#439115000000
1!
1%
#439120000000
0!
0%
#439125000000
1!
1%
#439130000000
0!
0%
#439135000000
1!
1%
#439140000000
0!
0%
#439145000000
1!
1%
#439150000000
0!
0%
#439155000000
1!
1%
#439160000000
0!
0%
#439165000000
1!
1%
#439170000000
0!
0%
#439175000000
1!
1%
#439180000000
0!
0%
#439185000000
1!
1%
#439190000000
0!
0%
#439195000000
1!
1%
#439200000000
0!
0%
#439205000000
1!
1%
#439210000000
0!
0%
#439215000000
1!
1%
#439220000000
0!
0%
#439225000000
1!
1%
#439230000000
0!
0%
#439235000000
1!
1%
#439240000000
0!
0%
#439245000000
1!
1%
#439250000000
0!
0%
#439255000000
1!
1%
#439260000000
0!
0%
#439265000000
1!
1%
#439270000000
0!
0%
#439275000000
1!
1%
#439280000000
0!
0%
#439285000000
1!
1%
#439290000000
0!
0%
#439295000000
1!
1%
#439300000000
0!
0%
#439305000000
1!
1%
#439310000000
0!
0%
#439315000000
1!
1%
#439320000000
0!
0%
#439325000000
1!
1%
#439330000000
0!
0%
#439335000000
1!
1%
#439340000000
0!
0%
#439345000000
1!
1%
#439350000000
0!
0%
#439355000000
1!
1%
#439360000000
0!
0%
#439365000000
1!
1%
#439370000000
0!
0%
#439375000000
1!
1%
#439380000000
0!
0%
#439385000000
1!
1%
#439390000000
0!
0%
#439395000000
1!
1%
#439400000000
0!
0%
#439405000000
1!
1%
#439410000000
0!
0%
#439415000000
1!
1%
#439420000000
0!
0%
#439425000000
1!
1%
#439430000000
0!
0%
#439435000000
1!
1%
#439440000000
0!
0%
#439445000000
1!
1%
#439450000000
0!
0%
#439455000000
1!
1%
#439460000000
0!
0%
#439465000000
1!
1%
#439470000000
0!
0%
#439475000000
1!
1%
#439480000000
0!
0%
#439485000000
1!
1%
#439490000000
0!
0%
#439495000000
1!
1%
#439500000000
0!
0%
#439505000000
1!
1%
#439510000000
0!
0%
#439515000000
1!
1%
#439520000000
0!
0%
#439525000000
1!
1%
#439530000000
0!
0%
#439535000000
1!
1%
#439540000000
0!
0%
#439545000000
1!
1%
#439550000000
0!
0%
#439555000000
1!
1%
#439560000000
0!
0%
#439565000000
1!
1%
#439570000000
0!
0%
#439575000000
1!
1%
#439580000000
0!
0%
#439585000000
1!
1%
#439590000000
0!
0%
#439595000000
1!
1%
#439600000000
0!
0%
#439605000000
1!
1%
#439610000000
0!
0%
#439615000000
1!
1%
#439620000000
0!
0%
#439625000000
1!
1%
#439630000000
0!
0%
#439635000000
1!
1%
#439640000000
0!
0%
#439645000000
1!
1%
#439650000000
0!
0%
#439655000000
1!
1%
#439660000000
0!
0%
#439665000000
1!
1%
#439670000000
0!
0%
#439675000000
1!
1%
#439680000000
0!
0%
#439685000000
1!
1%
#439690000000
0!
0%
#439695000000
1!
1%
#439700000000
0!
0%
#439705000000
1!
1%
#439710000000
0!
0%
#439715000000
1!
1%
#439720000000
0!
0%
#439725000000
1!
1%
#439730000000
0!
0%
#439735000000
1!
1%
#439740000000
0!
0%
#439745000000
1!
1%
#439750000000
0!
0%
#439755000000
1!
1%
#439760000000
0!
0%
#439765000000
1!
1%
#439770000000
0!
0%
#439775000000
1!
1%
#439780000000
0!
0%
#439785000000
1!
1%
#439790000000
0!
0%
#439795000000
1!
1%
#439800000000
0!
0%
#439805000000
1!
1%
#439810000000
0!
0%
#439815000000
1!
1%
#439820000000
0!
0%
#439825000000
1!
1%
#439830000000
0!
0%
#439835000000
1!
1%
#439840000000
0!
0%
#439845000000
1!
1%
#439850000000
0!
0%
#439855000000
1!
1%
#439860000000
0!
0%
#439865000000
1!
1%
#439870000000
0!
0%
#439875000000
1!
1%
#439880000000
0!
0%
#439885000000
1!
1%
#439890000000
0!
0%
#439895000000
1!
1%
#439900000000
0!
0%
#439905000000
1!
1%
#439910000000
0!
0%
#439915000000
1!
1%
#439920000000
0!
0%
#439925000000
1!
1%
#439930000000
0!
0%
#439935000000
1!
1%
#439940000000
0!
0%
#439945000000
1!
1%
#439950000000
0!
0%
#439955000000
1!
1%
#439960000000
0!
0%
#439965000000
1!
1%
#439970000000
0!
0%
#439975000000
1!
1%
#439980000000
0!
0%
#439985000000
1!
1%
#439990000000
0!
0%
#439995000000
1!
1%
#440000000000
0!
0%
#440005000000
1!
1%
#440010000000
0!
0%
#440015000000
1!
1%
#440020000000
0!
0%
#440025000000
1!
1%
#440030000000
0!
0%
#440035000000
1!
1%
#440040000000
0!
0%
#440045000000
1!
1%
#440050000000
0!
0%
#440055000000
1!
1%
#440060000000
0!
0%
#440065000000
1!
1%
#440070000000
0!
0%
#440075000000
1!
1%
#440080000000
0!
0%
#440085000000
1!
1%
#440090000000
0!
0%
#440095000000
1!
1%
#440100000000
0!
0%
#440105000000
1!
1%
#440110000000
0!
0%
#440115000000
1!
1%
#440120000000
0!
0%
#440125000000
1!
1%
#440130000000
0!
0%
#440135000000
1!
1%
#440140000000
0!
0%
#440145000000
1!
1%
#440150000000
0!
0%
#440155000000
1!
1%
#440160000000
0!
0%
#440165000000
1!
1%
#440170000000
0!
0%
#440175000000
1!
1%
#440180000000
0!
0%
#440185000000
1!
1%
#440190000000
0!
0%
#440195000000
1!
1%
#440200000000
0!
0%
#440205000000
1!
1%
#440210000000
0!
0%
#440215000000
1!
1%
#440220000000
0!
0%
#440225000000
1!
1%
#440230000000
0!
0%
#440235000000
1!
1%
#440240000000
0!
0%
#440245000000
1!
1%
#440250000000
0!
0%
#440255000000
1!
1%
#440260000000
0!
0%
#440265000000
1!
1%
#440270000000
0!
0%
#440275000000
1!
1%
#440280000000
0!
0%
#440285000000
1!
1%
#440290000000
0!
0%
#440295000000
1!
1%
#440300000000
0!
0%
#440305000000
1!
1%
#440310000000
0!
0%
#440315000000
1!
1%
#440320000000
0!
0%
#440325000000
1!
1%
#440330000000
0!
0%
#440335000000
1!
1%
#440340000000
0!
0%
#440345000000
1!
1%
#440350000000
0!
0%
#440355000000
1!
1%
#440360000000
0!
0%
#440365000000
1!
1%
#440370000000
0!
0%
#440375000000
1!
1%
#440380000000
0!
0%
#440385000000
1!
1%
#440390000000
0!
0%
#440395000000
1!
1%
#440400000000
0!
0%
#440405000000
1!
1%
#440410000000
0!
0%
#440415000000
1!
1%
#440420000000
0!
0%
#440425000000
1!
1%
#440430000000
0!
0%
#440435000000
1!
1%
#440440000000
0!
0%
#440445000000
1!
1%
#440450000000
0!
0%
#440455000000
1!
1%
#440460000000
0!
0%
#440465000000
1!
1%
#440470000000
0!
0%
#440475000000
1!
1%
#440480000000
0!
0%
#440485000000
1!
1%
#440490000000
0!
0%
#440495000000
1!
1%
#440500000000
0!
0%
#440505000000
1!
1%
#440510000000
0!
0%
#440515000000
1!
1%
#440520000000
0!
0%
#440525000000
1!
1%
#440530000000
0!
0%
#440535000000
1!
1%
#440540000000
0!
0%
#440545000000
1!
1%
#440550000000
0!
0%
#440555000000
1!
1%
#440560000000
0!
0%
#440565000000
1!
1%
#440570000000
0!
0%
#440575000000
1!
1%
#440580000000
0!
0%
#440585000000
1!
1%
#440590000000
0!
0%
#440595000000
1!
1%
#440600000000
0!
0%
#440605000000
1!
1%
#440610000000
0!
0%
#440615000000
1!
1%
#440620000000
0!
0%
#440625000000
1!
1%
#440630000000
0!
0%
#440635000000
1!
1%
#440640000000
0!
0%
#440645000000
1!
1%
#440650000000
0!
0%
#440655000000
1!
1%
#440660000000
0!
0%
#440665000000
1!
1%
#440670000000
0!
0%
#440675000000
1!
1%
#440680000000
0!
0%
#440685000000
1!
1%
#440690000000
0!
0%
#440695000000
1!
1%
#440700000000
0!
0%
#440705000000
1!
1%
#440710000000
0!
0%
#440715000000
1!
1%
#440720000000
0!
0%
#440725000000
1!
1%
#440730000000
0!
0%
#440735000000
1!
1%
#440740000000
0!
0%
#440745000000
1!
1%
#440750000000
0!
0%
#440755000000
1!
1%
#440760000000
0!
0%
#440765000000
1!
1%
#440770000000
0!
0%
#440775000000
1!
1%
#440780000000
0!
0%
#440785000000
1!
1%
#440790000000
0!
0%
#440795000000
1!
1%
#440800000000
0!
0%
#440805000000
1!
1%
#440810000000
0!
0%
#440815000000
1!
1%
#440820000000
0!
0%
#440825000000
1!
1%
#440830000000
0!
0%
#440835000000
1!
1%
#440840000000
0!
0%
#440845000000
1!
1%
#440850000000
0!
0%
#440855000000
1!
1%
#440860000000
0!
0%
#440865000000
1!
1%
#440870000000
0!
0%
#440875000000
1!
1%
#440880000000
0!
0%
#440885000000
1!
1%
#440890000000
0!
0%
#440895000000
1!
1%
#440900000000
0!
0%
#440905000000
1!
1%
#440910000000
0!
0%
#440915000000
1!
1%
#440920000000
0!
0%
#440925000000
1!
1%
#440930000000
0!
0%
#440935000000
1!
1%
#440940000000
0!
0%
#440945000000
1!
1%
#440950000000
0!
0%
#440955000000
1!
1%
#440960000000
0!
0%
#440965000000
1!
1%
#440970000000
0!
0%
#440975000000
1!
1%
#440980000000
0!
0%
#440985000000
1!
1%
#440990000000
0!
0%
#440995000000
1!
1%
#441000000000
0!
0%
#441005000000
1!
1%
#441010000000
0!
0%
#441015000000
1!
1%
#441020000000
0!
0%
#441025000000
1!
1%
#441030000000
0!
0%
#441035000000
1!
1%
#441040000000
0!
0%
#441045000000
1!
1%
#441050000000
0!
0%
#441055000000
1!
1%
#441060000000
0!
0%
#441065000000
1!
1%
#441070000000
0!
0%
#441075000000
1!
1%
#441080000000
0!
0%
#441085000000
1!
1%
#441090000000
0!
0%
#441095000000
1!
1%
#441100000000
0!
0%
#441105000000
1!
1%
#441110000000
0!
0%
#441115000000
1!
1%
#441120000000
0!
0%
#441125000000
1!
1%
#441130000000
0!
0%
#441135000000
1!
1%
#441140000000
0!
0%
#441145000000
1!
1%
#441150000000
0!
0%
#441155000000
1!
1%
#441160000000
0!
0%
#441165000000
1!
1%
#441170000000
0!
0%
#441175000000
1!
1%
#441180000000
0!
0%
#441185000000
1!
1%
#441190000000
0!
0%
#441195000000
1!
1%
#441200000000
0!
0%
#441205000000
1!
1%
#441210000000
0!
0%
#441215000000
1!
1%
#441220000000
0!
0%
#441225000000
1!
1%
#441230000000
0!
0%
#441235000000
1!
1%
#441240000000
0!
0%
#441245000000
1!
1%
#441250000000
0!
0%
#441255000000
1!
1%
#441260000000
0!
0%
#441265000000
1!
1%
#441270000000
0!
0%
#441275000000
1!
1%
#441280000000
0!
0%
#441285000000
1!
1%
#441290000000
0!
0%
#441295000000
1!
1%
#441300000000
0!
0%
#441305000000
1!
1%
#441310000000
0!
0%
#441315000000
1!
1%
#441320000000
0!
0%
#441325000000
1!
1%
#441330000000
0!
0%
#441335000000
1!
1%
#441340000000
0!
0%
#441345000000
1!
1%
#441350000000
0!
0%
#441355000000
1!
1%
#441360000000
0!
0%
#441365000000
1!
1%
#441370000000
0!
0%
#441375000000
1!
1%
#441380000000
0!
0%
#441385000000
1!
1%
#441390000000
0!
0%
#441395000000
1!
1%
#441400000000
0!
0%
#441405000000
1!
1%
#441410000000
0!
0%
#441415000000
1!
1%
#441420000000
0!
0%
#441425000000
1!
1%
#441430000000
0!
0%
#441435000000
1!
1%
#441440000000
0!
0%
#441445000000
1!
1%
#441450000000
0!
0%
#441455000000
1!
1%
#441460000000
0!
0%
#441465000000
1!
1%
#441470000000
0!
0%
#441475000000
1!
1%
#441480000000
0!
0%
#441485000000
1!
1%
#441490000000
0!
0%
#441495000000
1!
1%
#441500000000
0!
0%
#441505000000
1!
1%
#441510000000
0!
0%
#441515000000
1!
1%
#441520000000
0!
0%
#441525000000
1!
1%
#441530000000
0!
0%
#441535000000
1!
1%
#441540000000
0!
0%
#441545000000
1!
1%
#441550000000
0!
0%
#441555000000
1!
1%
#441560000000
0!
0%
#441565000000
1!
1%
#441570000000
0!
0%
#441575000000
1!
1%
#441580000000
0!
0%
#441585000000
1!
1%
#441590000000
0!
0%
#441595000000
1!
1%
#441600000000
0!
0%
#441605000000
1!
1%
#441610000000
0!
0%
#441615000000
1!
1%
#441620000000
0!
0%
#441625000000
1!
1%
#441630000000
0!
0%
#441635000000
1!
1%
#441640000000
0!
0%
#441645000000
1!
1%
#441650000000
0!
0%
#441655000000
1!
1%
#441660000000
0!
0%
#441665000000
1!
1%
#441670000000
0!
0%
#441675000000
1!
1%
#441680000000
0!
0%
#441685000000
1!
1%
#441690000000
0!
0%
#441695000000
1!
1%
#441700000000
0!
0%
#441705000000
1!
1%
#441710000000
0!
0%
#441715000000
1!
1%
#441720000000
0!
0%
#441725000000
1!
1%
#441730000000
0!
0%
#441735000000
1!
1%
#441740000000
0!
0%
#441745000000
1!
1%
#441750000000
0!
0%
#441755000000
1!
1%
#441760000000
0!
0%
#441765000000
1!
1%
#441770000000
0!
0%
#441775000000
1!
1%
#441780000000
0!
0%
#441785000000
1!
1%
#441790000000
0!
0%
#441795000000
1!
1%
#441800000000
0!
0%
#441805000000
1!
1%
#441810000000
0!
0%
#441815000000
1!
1%
#441820000000
0!
0%
#441825000000
1!
1%
#441830000000
0!
0%
#441835000000
1!
1%
#441840000000
0!
0%
#441845000000
1!
1%
#441850000000
0!
0%
#441855000000
1!
1%
#441860000000
0!
0%
#441865000000
1!
1%
#441870000000
0!
0%
#441875000000
1!
1%
#441880000000
0!
0%
#441885000000
1!
1%
#441890000000
0!
0%
#441895000000
1!
1%
#441900000000
0!
0%
#441905000000
1!
1%
#441910000000
0!
0%
#441915000000
1!
1%
#441920000000
0!
0%
#441925000000
1!
1%
#441930000000
0!
0%
#441935000000
1!
1%
#441940000000
0!
0%
#441945000000
1!
1%
#441950000000
0!
0%
#441955000000
1!
1%
#441960000000
0!
0%
#441965000000
1!
1%
#441970000000
0!
0%
#441975000000
1!
1%
#441980000000
0!
0%
#441985000000
1!
1%
#441990000000
0!
0%
#441995000000
1!
1%
#442000000000
0!
0%
#442005000000
1!
1%
#442010000000
0!
0%
#442015000000
1!
1%
#442020000000
0!
0%
#442025000000
1!
1%
#442030000000
0!
0%
#442035000000
1!
1%
#442040000000
0!
0%
#442045000000
1!
1%
#442050000000
0!
0%
#442055000000
1!
1%
#442060000000
0!
0%
#442065000000
1!
1%
#442070000000
0!
0%
#442075000000
1!
1%
#442080000000
0!
0%
#442085000000
1!
1%
#442090000000
0!
0%
#442095000000
1!
1%
#442100000000
0!
0%
#442105000000
1!
1%
#442110000000
0!
0%
#442115000000
1!
1%
#442120000000
0!
0%
#442125000000
1!
1%
#442130000000
0!
0%
#442135000000
1!
1%
#442140000000
0!
0%
#442145000000
1!
1%
#442150000000
0!
0%
#442155000000
1!
1%
#442160000000
0!
0%
#442165000000
1!
1%
#442170000000
0!
0%
#442175000000
1!
1%
#442180000000
0!
0%
#442185000000
1!
1%
#442190000000
0!
0%
#442195000000
1!
1%
#442200000000
0!
0%
#442205000000
1!
1%
#442210000000
0!
0%
#442215000000
1!
1%
#442220000000
0!
0%
#442225000000
1!
1%
#442230000000
0!
0%
#442235000000
1!
1%
#442240000000
0!
0%
#442245000000
1!
1%
#442250000000
0!
0%
#442255000000
1!
1%
#442260000000
0!
0%
#442265000000
1!
1%
#442270000000
0!
0%
#442275000000
1!
1%
#442280000000
0!
0%
#442285000000
1!
1%
#442290000000
0!
0%
#442295000000
1!
1%
#442300000000
0!
0%
#442305000000
1!
1%
#442310000000
0!
0%
#442315000000
1!
1%
#442320000000
0!
0%
#442325000000
1!
1%
#442330000000
0!
0%
#442335000000
1!
1%
#442340000000
0!
0%
#442345000000
1!
1%
#442350000000
0!
0%
#442355000000
1!
1%
#442360000000
0!
0%
#442365000000
1!
1%
#442370000000
0!
0%
#442375000000
1!
1%
#442380000000
0!
0%
#442385000000
1!
1%
#442390000000
0!
0%
#442395000000
1!
1%
#442400000000
0!
0%
#442405000000
1!
1%
#442410000000
0!
0%
#442415000000
1!
1%
#442420000000
0!
0%
#442425000000
1!
1%
#442430000000
0!
0%
#442435000000
1!
1%
#442440000000
0!
0%
#442445000000
1!
1%
#442450000000
0!
0%
#442455000000
1!
1%
#442460000000
0!
0%
#442465000000
1!
1%
#442470000000
0!
0%
#442475000000
1!
1%
#442480000000
0!
0%
#442485000000
1!
1%
#442490000000
0!
0%
#442495000000
1!
1%
#442500000000
0!
0%
#442505000000
1!
1%
#442510000000
0!
0%
#442515000000
1!
1%
#442520000000
0!
0%
#442525000000
1!
1%
#442530000000
0!
0%
#442535000000
1!
1%
#442540000000
0!
0%
#442545000000
1!
1%
#442550000000
0!
0%
#442555000000
1!
1%
#442560000000
0!
0%
#442565000000
1!
1%
#442570000000
0!
0%
#442575000000
1!
1%
#442580000000
0!
0%
#442585000000
1!
1%
#442590000000
0!
0%
#442595000000
1!
1%
#442600000000
0!
0%
#442605000000
1!
1%
#442610000000
0!
0%
#442615000000
1!
1%
#442620000000
0!
0%
#442625000000
1!
1%
#442630000000
0!
0%
#442635000000
1!
1%
#442640000000
0!
0%
#442645000000
1!
1%
#442650000000
0!
0%
#442655000000
1!
1%
#442660000000
0!
0%
#442665000000
1!
1%
#442670000000
0!
0%
#442675000000
1!
1%
#442680000000
0!
0%
#442685000000
1!
1%
#442690000000
0!
0%
#442695000000
1!
1%
#442700000000
0!
0%
#442705000000
1!
1%
#442710000000
0!
0%
#442715000000
1!
1%
#442720000000
0!
0%
#442725000000
1!
1%
#442730000000
0!
0%
#442735000000
1!
1%
#442740000000
0!
0%
#442745000000
1!
1%
#442750000000
0!
0%
#442755000000
1!
1%
#442760000000
0!
0%
#442765000000
1!
1%
#442770000000
0!
0%
#442775000000
1!
1%
#442780000000
0!
0%
#442785000000
1!
1%
#442790000000
0!
0%
#442795000000
1!
1%
#442800000000
0!
0%
#442805000000
1!
1%
#442810000000
0!
0%
#442815000000
1!
1%
#442820000000
0!
0%
#442825000000
1!
1%
#442830000000
0!
0%
#442835000000
1!
1%
#442840000000
0!
0%
#442845000000
1!
1%
#442850000000
0!
0%
#442855000000
1!
1%
#442860000000
0!
0%
#442865000000
1!
1%
#442870000000
0!
0%
#442875000000
1!
1%
#442880000000
0!
0%
#442885000000
1!
1%
#442890000000
0!
0%
#442895000000
1!
1%
#442900000000
0!
0%
#442905000000
1!
1%
#442910000000
0!
0%
#442915000000
1!
1%
#442920000000
0!
0%
#442925000000
1!
1%
#442930000000
0!
0%
#442935000000
1!
1%
#442940000000
0!
0%
#442945000000
1!
1%
#442950000000
0!
0%
#442955000000
1!
1%
#442960000000
0!
0%
#442965000000
1!
1%
#442970000000
0!
0%
#442975000000
1!
1%
#442980000000
0!
0%
#442985000000
1!
1%
#442990000000
0!
0%
#442995000000
1!
1%
#443000000000
0!
0%
#443005000000
1!
1%
#443010000000
0!
0%
#443015000000
1!
1%
#443020000000
0!
0%
#443025000000
1!
1%
#443030000000
0!
0%
#443035000000
1!
1%
#443040000000
0!
0%
#443045000000
1!
1%
#443050000000
0!
0%
#443055000000
1!
1%
#443060000000
0!
0%
#443065000000
1!
1%
#443070000000
0!
0%
#443075000000
1!
1%
#443080000000
0!
0%
#443085000000
1!
1%
#443090000000
0!
0%
#443095000000
1!
1%
#443100000000
0!
0%
#443105000000
1!
1%
#443110000000
0!
0%
#443115000000
1!
1%
#443120000000
0!
0%
#443125000000
1!
1%
#443130000000
0!
0%
#443135000000
1!
1%
#443140000000
0!
0%
#443145000000
1!
1%
#443150000000
0!
0%
#443155000000
1!
1%
#443160000000
0!
0%
#443165000000
1!
1%
#443170000000
0!
0%
#443175000000
1!
1%
#443180000000
0!
0%
#443185000000
1!
1%
#443190000000
0!
0%
#443195000000
1!
1%
#443200000000
0!
0%
#443205000000
1!
1%
#443210000000
0!
0%
#443215000000
1!
1%
#443220000000
0!
0%
#443225000000
1!
1%
#443230000000
0!
0%
#443235000000
1!
1%
#443240000000
0!
0%
#443245000000
1!
1%
#443250000000
0!
0%
#443255000000
1!
1%
#443260000000
0!
0%
#443265000000
1!
1%
#443270000000
0!
0%
#443275000000
1!
1%
#443280000000
0!
0%
#443285000000
1!
1%
#443290000000
0!
0%
#443295000000
1!
1%
#443300000000
0!
0%
#443305000000
1!
1%
#443310000000
0!
0%
#443315000000
1!
1%
#443320000000
0!
0%
#443325000000
1!
1%
#443330000000
0!
0%
#443335000000
1!
1%
#443340000000
0!
0%
#443345000000
1!
1%
#443350000000
0!
0%
#443355000000
1!
1%
#443360000000
0!
0%
#443365000000
1!
1%
#443370000000
0!
0%
#443375000000
1!
1%
#443380000000
0!
0%
#443385000000
1!
1%
#443390000000
0!
0%
#443395000000
1!
1%
#443400000000
0!
0%
#443405000000
1!
1%
#443410000000
0!
0%
#443415000000
1!
1%
#443420000000
0!
0%
#443425000000
1!
1%
#443430000000
0!
0%
#443435000000
1!
1%
#443440000000
0!
0%
#443445000000
1!
1%
#443450000000
0!
0%
#443455000000
1!
1%
#443460000000
0!
0%
#443465000000
1!
1%
#443470000000
0!
0%
#443475000000
1!
1%
#443480000000
0!
0%
#443485000000
1!
1%
#443490000000
0!
0%
#443495000000
1!
1%
#443500000000
0!
0%
#443505000000
1!
1%
#443510000000
0!
0%
#443515000000
1!
1%
#443520000000
0!
0%
#443525000000
1!
1%
#443530000000
0!
0%
#443535000000
1!
1%
#443540000000
0!
0%
#443545000000
1!
1%
#443550000000
0!
0%
#443555000000
1!
1%
#443560000000
0!
0%
#443565000000
1!
1%
#443570000000
0!
0%
#443575000000
1!
1%
#443580000000
0!
0%
#443585000000
1!
1%
#443590000000
0!
0%
#443595000000
1!
1%
#443600000000
0!
0%
#443605000000
1!
1%
#443610000000
0!
0%
#443615000000
1!
1%
#443620000000
0!
0%
#443625000000
1!
1%
#443630000000
0!
0%
#443635000000
1!
1%
#443640000000
0!
0%
#443645000000
1!
1%
#443650000000
0!
0%
#443655000000
1!
1%
#443660000000
0!
0%
#443665000000
1!
1%
#443670000000
0!
0%
#443675000000
1!
1%
#443680000000
0!
0%
#443685000000
1!
1%
#443690000000
0!
0%
#443695000000
1!
1%
#443700000000
0!
0%
#443705000000
1!
1%
#443710000000
0!
0%
#443715000000
1!
1%
#443720000000
0!
0%
#443725000000
1!
1%
#443730000000
0!
0%
#443735000000
1!
1%
#443740000000
0!
0%
#443745000000
1!
1%
#443750000000
0!
0%
#443755000000
1!
1%
#443760000000
0!
0%
#443765000000
1!
1%
#443770000000
0!
0%
#443775000000
1!
1%
#443780000000
0!
0%
#443785000000
1!
1%
#443790000000
0!
0%
#443795000000
1!
1%
#443800000000
0!
0%
#443805000000
1!
1%
#443810000000
0!
0%
#443815000000
1!
1%
#443820000000
0!
0%
#443825000000
1!
1%
#443830000000
0!
0%
#443835000000
1!
1%
#443840000000
0!
0%
#443845000000
1!
1%
#443850000000
0!
0%
#443855000000
1!
1%
#443860000000
0!
0%
#443865000000
1!
1%
#443870000000
0!
0%
#443875000000
1!
1%
#443880000000
0!
0%
#443885000000
1!
1%
#443890000000
0!
0%
#443895000000
1!
1%
#443900000000
0!
0%
#443905000000
1!
1%
#443910000000
0!
0%
#443915000000
1!
1%
#443920000000
0!
0%
#443925000000
1!
1%
#443930000000
0!
0%
#443935000000
1!
1%
#443940000000
0!
0%
#443945000000
1!
1%
#443950000000
0!
0%
#443955000000
1!
1%
#443960000000
0!
0%
#443965000000
1!
1%
#443970000000
0!
0%
#443975000000
1!
1%
#443980000000
0!
0%
#443985000000
1!
1%
#443990000000
0!
0%
#443995000000
1!
1%
#444000000000
0!
0%
#444005000000
1!
1%
#444010000000
0!
0%
#444015000000
1!
1%
#444020000000
0!
0%
#444025000000
1!
1%
#444030000000
0!
0%
#444035000000
1!
1%
#444040000000
0!
0%
#444045000000
1!
1%
#444050000000
0!
0%
#444055000000
1!
1%
#444060000000
0!
0%
#444065000000
1!
1%
#444070000000
0!
0%
#444075000000
1!
1%
#444080000000
0!
0%
#444085000000
1!
1%
#444090000000
0!
0%
#444095000000
1!
1%
#444100000000
0!
0%
#444105000000
1!
1%
#444110000000
0!
0%
#444115000000
1!
1%
#444120000000
0!
0%
#444125000000
1!
1%
#444130000000
0!
0%
#444135000000
1!
1%
#444140000000
0!
0%
#444145000000
1!
1%
#444150000000
0!
0%
#444155000000
1!
1%
#444160000000
0!
0%
#444165000000
1!
1%
#444170000000
0!
0%
#444175000000
1!
1%
#444180000000
0!
0%
#444185000000
1!
1%
#444190000000
0!
0%
#444195000000
1!
1%
#444200000000
0!
0%
#444205000000
1!
1%
#444210000000
0!
0%
#444215000000
1!
1%
#444220000000
0!
0%
#444225000000
1!
1%
#444230000000
0!
0%
#444235000000
1!
1%
#444240000000
0!
0%
#444245000000
1!
1%
#444250000000
0!
0%
#444255000000
1!
1%
#444260000000
0!
0%
#444265000000
1!
1%
#444270000000
0!
0%
#444275000000
1!
1%
#444280000000
0!
0%
#444285000000
1!
1%
#444290000000
0!
0%
#444295000000
1!
1%
#444300000000
0!
0%
#444305000000
1!
1%
#444310000000
0!
0%
#444315000000
1!
1%
#444320000000
0!
0%
#444325000000
1!
1%
#444330000000
0!
0%
#444335000000
1!
1%
#444340000000
0!
0%
#444345000000
1!
1%
#444350000000
0!
0%
#444355000000
1!
1%
#444360000000
0!
0%
#444365000000
1!
1%
#444370000000
0!
0%
#444375000000
1!
1%
#444380000000
0!
0%
#444385000000
1!
1%
#444390000000
0!
0%
#444395000000
1!
1%
#444400000000
0!
0%
#444405000000
1!
1%
#444410000000
0!
0%
#444415000000
1!
1%
#444420000000
0!
0%
#444425000000
1!
1%
#444430000000
0!
0%
#444435000000
1!
1%
#444440000000
0!
0%
#444445000000
1!
1%
#444450000000
0!
0%
#444455000000
1!
1%
#444460000000
0!
0%
#444465000000
1!
1%
#444470000000
0!
0%
#444475000000
1!
1%
#444480000000
0!
0%
#444485000000
1!
1%
#444490000000
0!
0%
#444495000000
1!
1%
#444500000000
0!
0%
#444505000000
1!
1%
#444510000000
0!
0%
#444515000000
1!
1%
#444520000000
0!
0%
#444525000000
1!
1%
#444530000000
0!
0%
#444535000000
1!
1%
#444540000000
0!
0%
#444545000000
1!
1%
#444550000000
0!
0%
#444555000000
1!
1%
#444560000000
0!
0%
#444565000000
1!
1%
#444570000000
0!
0%
#444575000000
1!
1%
#444580000000
0!
0%
#444585000000
1!
1%
#444590000000
0!
0%
#444595000000
1!
1%
#444600000000
0!
0%
#444605000000
1!
1%
#444610000000
0!
0%
#444615000000
1!
1%
#444620000000
0!
0%
#444625000000
1!
1%
#444630000000
0!
0%
#444635000000
1!
1%
#444640000000
0!
0%
#444645000000
1!
1%
#444650000000
0!
0%
#444655000000
1!
1%
#444660000000
0!
0%
#444665000000
1!
1%
#444670000000
0!
0%
#444675000000
1!
1%
#444680000000
0!
0%
#444685000000
1!
1%
#444690000000
0!
0%
#444695000000
1!
1%
#444700000000
0!
0%
#444705000000
1!
1%
#444710000000
0!
0%
#444715000000
1!
1%
#444720000000
0!
0%
#444725000000
1!
1%
#444730000000
0!
0%
#444735000000
1!
1%
#444740000000
0!
0%
#444745000000
1!
1%
#444750000000
0!
0%
#444755000000
1!
1%
#444760000000
0!
0%
#444765000000
1!
1%
#444770000000
0!
0%
#444775000000
1!
1%
#444780000000
0!
0%
#444785000000
1!
1%
#444790000000
0!
0%
#444795000000
1!
1%
#444800000000
0!
0%
#444805000000
1!
1%
#444810000000
0!
0%
#444815000000
1!
1%
#444820000000
0!
0%
#444825000000
1!
1%
#444830000000
0!
0%
#444835000000
1!
1%
#444840000000
0!
0%
#444845000000
1!
1%
#444850000000
0!
0%
#444855000000
1!
1%
#444860000000
0!
0%
#444865000000
1!
1%
#444870000000
0!
0%
#444875000000
1!
1%
#444880000000
0!
0%
#444885000000
1!
1%
#444890000000
0!
0%
#444895000000
1!
1%
#444900000000
0!
0%
#444905000000
1!
1%
#444910000000
0!
0%
#444915000000
1!
1%
#444920000000
0!
0%
#444925000000
1!
1%
#444930000000
0!
0%
#444935000000
1!
1%
#444940000000
0!
0%
#444945000000
1!
1%
#444950000000
0!
0%
#444955000000
1!
1%
#444960000000
0!
0%
#444965000000
1!
1%
#444970000000
0!
0%
#444975000000
1!
1%
#444980000000
0!
0%
#444985000000
1!
1%
#444990000000
0!
0%
#444995000000
1!
1%
#445000000000
0!
0%
#445005000000
1!
1%
#445010000000
0!
0%
#445015000000
1!
1%
#445020000000
0!
0%
#445025000000
1!
1%
#445030000000
0!
0%
#445035000000
1!
1%
#445040000000
0!
0%
#445045000000
1!
1%
#445050000000
0!
0%
#445055000000
1!
1%
#445060000000
0!
0%
#445065000000
1!
1%
#445070000000
0!
0%
#445075000000
1!
1%
#445080000000
0!
0%
#445085000000
1!
1%
#445090000000
0!
0%
#445095000000
1!
1%
#445100000000
0!
0%
#445105000000
1!
1%
#445110000000
0!
0%
#445115000000
1!
1%
#445120000000
0!
0%
#445125000000
1!
1%
#445130000000
0!
0%
#445135000000
1!
1%
#445140000000
0!
0%
#445145000000
1!
1%
#445150000000
0!
0%
#445155000000
1!
1%
#445160000000
0!
0%
#445165000000
1!
1%
#445170000000
0!
0%
#445175000000
1!
1%
#445180000000
0!
0%
#445185000000
1!
1%
#445190000000
0!
0%
#445195000000
1!
1%
#445200000000
0!
0%
#445205000000
1!
1%
#445210000000
0!
0%
#445215000000
1!
1%
#445220000000
0!
0%
#445225000000
1!
1%
#445230000000
0!
0%
#445235000000
1!
1%
#445240000000
0!
0%
#445245000000
1!
1%
#445250000000
0!
0%
#445255000000
1!
1%
#445260000000
0!
0%
#445265000000
1!
1%
#445270000000
0!
0%
#445275000000
1!
1%
#445280000000
0!
0%
#445285000000
1!
1%
#445290000000
0!
0%
#445295000000
1!
1%
#445300000000
0!
0%
#445305000000
1!
1%
#445310000000
0!
0%
#445315000000
1!
1%
#445320000000
0!
0%
#445325000000
1!
1%
#445330000000
0!
0%
#445335000000
1!
1%
#445340000000
0!
0%
#445345000000
1!
1%
#445350000000
0!
0%
#445355000000
1!
1%
#445360000000
0!
0%
#445365000000
1!
1%
#445370000000
0!
0%
#445375000000
1!
1%
#445380000000
0!
0%
#445385000000
1!
1%
#445390000000
0!
0%
#445395000000
1!
1%
#445400000000
0!
0%
#445405000000
1!
1%
#445410000000
0!
0%
#445415000000
1!
1%
#445420000000
0!
0%
#445425000000
1!
1%
#445430000000
0!
0%
#445435000000
1!
1%
#445440000000
0!
0%
#445445000000
1!
1%
#445450000000
0!
0%
#445455000000
1!
1%
#445460000000
0!
0%
#445465000000
1!
1%
#445470000000
0!
0%
#445475000000
1!
1%
#445480000000
0!
0%
#445485000000
1!
1%
#445490000000
0!
0%
#445495000000
1!
1%
#445500000000
0!
0%
#445505000000
1!
1%
#445510000000
0!
0%
#445515000000
1!
1%
#445520000000
0!
0%
#445525000000
1!
1%
#445530000000
0!
0%
#445535000000
1!
1%
#445540000000
0!
0%
#445545000000
1!
1%
#445550000000
0!
0%
#445555000000
1!
1%
#445560000000
0!
0%
#445565000000
1!
1%
#445570000000
0!
0%
#445575000000
1!
1%
#445580000000
0!
0%
#445585000000
1!
1%
#445590000000
0!
0%
#445595000000
1!
1%
#445600000000
0!
0%
#445605000000
1!
1%
#445610000000
0!
0%
#445615000000
1!
1%
#445620000000
0!
0%
#445625000000
1!
1%
#445630000000
0!
0%
#445635000000
1!
1%
#445640000000
0!
0%
#445645000000
1!
1%
#445650000000
0!
0%
#445655000000
1!
1%
#445660000000
0!
0%
#445665000000
1!
1%
#445670000000
0!
0%
#445675000000
1!
1%
#445680000000
0!
0%
#445685000000
1!
1%
#445690000000
0!
0%
#445695000000
1!
1%
#445700000000
0!
0%
#445705000000
1!
1%
#445710000000
0!
0%
#445715000000
1!
1%
#445720000000
0!
0%
#445725000000
1!
1%
#445730000000
0!
0%
#445735000000
1!
1%
#445740000000
0!
0%
#445745000000
1!
1%
#445750000000
0!
0%
#445755000000
1!
1%
#445760000000
0!
0%
#445765000000
1!
1%
#445770000000
0!
0%
#445775000000
1!
1%
#445780000000
0!
0%
#445785000000
1!
1%
#445790000000
0!
0%
#445795000000
1!
1%
#445800000000
0!
0%
#445805000000
1!
1%
#445810000000
0!
0%
#445815000000
1!
1%
#445820000000
0!
0%
#445825000000
1!
1%
#445830000000
0!
0%
#445835000000
1!
1%
#445840000000
0!
0%
#445845000000
1!
1%
#445850000000
0!
0%
#445855000000
1!
1%
#445860000000
0!
0%
#445865000000
1!
1%
#445870000000
0!
0%
#445875000000
1!
1%
#445880000000
0!
0%
#445885000000
1!
1%
#445890000000
0!
0%
#445895000000
1!
1%
#445900000000
0!
0%
#445905000000
1!
1%
#445910000000
0!
0%
#445915000000
1!
1%
#445920000000
0!
0%
#445925000000
1!
1%
#445930000000
0!
0%
#445935000000
1!
1%
#445940000000
0!
0%
#445945000000
1!
1%
#445950000000
0!
0%
#445955000000
1!
1%
#445960000000
0!
0%
#445965000000
1!
1%
#445970000000
0!
0%
#445975000000
1!
1%
#445980000000
0!
0%
#445985000000
1!
1%
#445990000000
0!
0%
#445995000000
1!
1%
#446000000000
0!
0%
#446005000000
1!
1%
#446010000000
0!
0%
#446015000000
1!
1%
#446020000000
0!
0%
#446025000000
1!
1%
#446030000000
0!
0%
#446035000000
1!
1%
#446040000000
0!
0%
#446045000000
1!
1%
#446050000000
0!
0%
#446055000000
1!
1%
#446060000000
0!
0%
#446065000000
1!
1%
#446070000000
0!
0%
#446075000000
1!
1%
#446080000000
0!
0%
#446085000000
1!
1%
#446090000000
0!
0%
#446095000000
1!
1%
#446100000000
0!
0%
#446105000000
1!
1%
#446110000000
0!
0%
#446115000000
1!
1%
#446120000000
0!
0%
#446125000000
1!
1%
#446130000000
0!
0%
#446135000000
1!
1%
#446140000000
0!
0%
#446145000000
1!
1%
#446150000000
0!
0%
#446155000000
1!
1%
#446160000000
0!
0%
#446165000000
1!
1%
#446170000000
0!
0%
#446175000000
1!
1%
#446180000000
0!
0%
#446185000000
1!
1%
#446190000000
0!
0%
#446195000000
1!
1%
#446200000000
0!
0%
#446205000000
1!
1%
#446210000000
0!
0%
#446215000000
1!
1%
#446220000000
0!
0%
#446225000000
1!
1%
#446230000000
0!
0%
#446235000000
1!
1%
#446240000000
0!
0%
#446245000000
1!
1%
#446250000000
0!
0%
#446255000000
1!
1%
#446260000000
0!
0%
#446265000000
1!
1%
#446270000000
0!
0%
#446275000000
1!
1%
#446280000000
0!
0%
#446285000000
1!
1%
#446290000000
0!
0%
#446295000000
1!
1%
#446300000000
0!
0%
#446305000000
1!
1%
#446310000000
0!
0%
#446315000000
1!
1%
#446320000000
0!
0%
#446325000000
1!
1%
#446330000000
0!
0%
#446335000000
1!
1%
#446340000000
0!
0%
#446345000000
1!
1%
#446350000000
0!
0%
#446355000000
1!
1%
#446360000000
0!
0%
#446365000000
1!
1%
#446370000000
0!
0%
#446375000000
1!
1%
#446380000000
0!
0%
#446385000000
1!
1%
#446390000000
0!
0%
#446395000000
1!
1%
#446400000000
0!
0%
#446405000000
1!
1%
#446410000000
0!
0%
#446415000000
1!
1%
#446420000000
0!
0%
#446425000000
1!
1%
#446430000000
0!
0%
#446435000000
1!
1%
#446440000000
0!
0%
#446445000000
1!
1%
#446450000000
0!
0%
#446455000000
1!
1%
#446460000000
0!
0%
#446465000000
1!
1%
#446470000000
0!
0%
#446475000000
1!
1%
#446480000000
0!
0%
#446485000000
1!
1%
#446490000000
0!
0%
#446495000000
1!
1%
#446500000000
0!
0%
#446505000000
1!
1%
#446510000000
0!
0%
#446515000000
1!
1%
#446520000000
0!
0%
#446525000000
1!
1%
#446530000000
0!
0%
#446535000000
1!
1%
#446540000000
0!
0%
#446545000000
1!
1%
#446550000000
0!
0%
#446555000000
1!
1%
#446560000000
0!
0%
#446565000000
1!
1%
#446570000000
0!
0%
#446575000000
1!
1%
#446580000000
0!
0%
#446585000000
1!
1%
#446590000000
0!
0%
#446595000000
1!
1%
#446600000000
0!
0%
#446605000000
1!
1%
#446610000000
0!
0%
#446615000000
1!
1%
#446620000000
0!
0%
#446625000000
1!
1%
#446630000000
0!
0%
#446635000000
1!
1%
#446640000000
0!
0%
#446645000000
1!
1%
#446650000000
0!
0%
#446655000000
1!
1%
#446660000000
0!
0%
#446665000000
1!
1%
#446670000000
0!
0%
#446675000000
1!
1%
#446680000000
0!
0%
#446685000000
1!
1%
#446690000000
0!
0%
#446695000000
1!
1%
#446700000000
0!
0%
#446705000000
1!
1%
#446710000000
0!
0%
#446715000000
1!
1%
#446720000000
0!
0%
#446725000000
1!
1%
#446730000000
0!
0%
#446735000000
1!
1%
#446740000000
0!
0%
#446745000000
1!
1%
#446750000000
0!
0%
#446755000000
1!
1%
#446760000000
0!
0%
#446765000000
1!
1%
#446770000000
0!
0%
#446775000000
1!
1%
#446780000000
0!
0%
#446785000000
1!
1%
#446790000000
0!
0%
#446795000000
1!
1%
#446800000000
0!
0%
#446805000000
1!
1%
#446810000000
0!
0%
#446815000000
1!
1%
#446820000000
0!
0%
#446825000000
1!
1%
#446830000000
0!
0%
#446835000000
1!
1%
#446840000000
0!
0%
#446845000000
1!
1%
#446850000000
0!
0%
#446855000000
1!
1%
#446860000000
0!
0%
#446865000000
1!
1%
#446870000000
0!
0%
#446875000000
1!
1%
#446880000000
0!
0%
#446885000000
1!
1%
#446890000000
0!
0%
#446895000000
1!
1%
#446900000000
0!
0%
#446905000000
1!
1%
#446910000000
0!
0%
#446915000000
1!
1%
#446920000000
0!
0%
#446925000000
1!
1%
#446930000000
0!
0%
#446935000000
1!
1%
#446940000000
0!
0%
#446945000000
1!
1%
#446950000000
0!
0%
#446955000000
1!
1%
#446960000000
0!
0%
#446965000000
1!
1%
#446970000000
0!
0%
#446975000000
1!
1%
#446980000000
0!
0%
#446985000000
1!
1%
#446990000000
0!
0%
#446995000000
1!
1%
#447000000000
0!
0%
#447005000000
1!
1%
#447010000000
0!
0%
#447015000000
1!
1%
#447020000000
0!
0%
#447025000000
1!
1%
#447030000000
0!
0%
#447035000000
1!
1%
#447040000000
0!
0%
#447045000000
1!
1%
#447050000000
0!
0%
#447055000000
1!
1%
#447060000000
0!
0%
#447065000000
1!
1%
#447070000000
0!
0%
#447075000000
1!
1%
#447080000000
0!
0%
#447085000000
1!
1%
#447090000000
0!
0%
#447095000000
1!
1%
#447100000000
0!
0%
#447105000000
1!
1%
#447110000000
0!
0%
#447115000000
1!
1%
#447120000000
0!
0%
#447125000000
1!
1%
#447130000000
0!
0%
#447135000000
1!
1%
#447140000000
0!
0%
#447145000000
1!
1%
#447150000000
0!
0%
#447155000000
1!
1%
#447160000000
0!
0%
#447165000000
1!
1%
#447170000000
0!
0%
#447175000000
1!
1%
#447180000000
0!
0%
#447185000000
1!
1%
#447190000000
0!
0%
#447195000000
1!
1%
#447200000000
0!
0%
#447205000000
1!
1%
#447210000000
0!
0%
#447215000000
1!
1%
#447220000000
0!
0%
#447225000000
1!
1%
#447230000000
0!
0%
#447235000000
1!
1%
#447240000000
0!
0%
#447245000000
1!
1%
#447250000000
0!
0%
#447255000000
1!
1%
#447260000000
0!
0%
#447265000000
1!
1%
#447270000000
0!
0%
#447275000000
1!
1%
#447280000000
0!
0%
#447285000000
1!
1%
#447290000000
0!
0%
#447295000000
1!
1%
#447300000000
0!
0%
#447305000000
1!
1%
#447310000000
0!
0%
#447315000000
1!
1%
#447320000000
0!
0%
#447325000000
1!
1%
#447330000000
0!
0%
#447335000000
1!
1%
#447340000000
0!
0%
#447345000000
1!
1%
#447350000000
0!
0%
#447355000000
1!
1%
#447360000000
0!
0%
#447365000000
1!
1%
#447370000000
0!
0%
#447375000000
1!
1%
#447380000000
0!
0%
#447385000000
1!
1%
#447390000000
0!
0%
#447395000000
1!
1%
#447400000000
0!
0%
#447405000000
1!
1%
#447410000000
0!
0%
#447415000000
1!
1%
#447420000000
0!
0%
#447425000000
1!
1%
#447430000000
0!
0%
#447435000000
1!
1%
#447440000000
0!
0%
#447445000000
1!
1%
#447450000000
0!
0%
#447455000000
1!
1%
#447460000000
0!
0%
#447465000000
1!
1%
#447470000000
0!
0%
#447475000000
1!
1%
#447480000000
0!
0%
#447485000000
1!
1%
#447490000000
0!
0%
#447495000000
1!
1%
#447500000000
0!
0%
#447505000000
1!
1%
#447510000000
0!
0%
#447515000000
1!
1%
#447520000000
0!
0%
#447525000000
1!
1%
#447530000000
0!
0%
#447535000000
1!
1%
#447540000000
0!
0%
#447545000000
1!
1%
#447550000000
0!
0%
#447555000000
1!
1%
#447560000000
0!
0%
#447565000000
1!
1%
#447570000000
0!
0%
#447575000000
1!
1%
#447580000000
0!
0%
#447585000000
1!
1%
#447590000000
0!
0%
#447595000000
1!
1%
#447600000000
0!
0%
#447605000000
1!
1%
#447610000000
0!
0%
#447615000000
1!
1%
#447620000000
0!
0%
#447625000000
1!
1%
#447630000000
0!
0%
#447635000000
1!
1%
#447640000000
0!
0%
#447645000000
1!
1%
#447650000000
0!
0%
#447655000000
1!
1%
#447660000000
0!
0%
#447665000000
1!
1%
#447670000000
0!
0%
#447675000000
1!
1%
#447680000000
0!
0%
#447685000000
1!
1%
#447690000000
0!
0%
#447695000000
1!
1%
#447700000000
0!
0%
#447705000000
1!
1%
#447710000000
0!
0%
#447715000000
1!
1%
#447720000000
0!
0%
#447725000000
1!
1%
#447730000000
0!
0%
#447735000000
1!
1%
#447740000000
0!
0%
#447745000000
1!
1%
#447750000000
0!
0%
#447755000000
1!
1%
#447760000000
0!
0%
#447765000000
1!
1%
#447770000000
0!
0%
#447775000000
1!
1%
#447780000000
0!
0%
#447785000000
1!
1%
#447790000000
0!
0%
#447795000000
1!
1%
#447800000000
0!
0%
#447805000000
1!
1%
#447810000000
0!
0%
#447815000000
1!
1%
#447820000000
0!
0%
#447825000000
1!
1%
#447830000000
0!
0%
#447835000000
1!
1%
#447840000000
0!
0%
#447845000000
1!
1%
#447850000000
0!
0%
#447855000000
1!
1%
#447860000000
0!
0%
#447865000000
1!
1%
#447870000000
0!
0%
#447875000000
1!
1%
#447880000000
0!
0%
#447885000000
1!
1%
#447890000000
0!
0%
#447895000000
1!
1%
#447900000000
0!
0%
#447905000000
1!
1%
#447910000000
0!
0%
#447915000000
1!
1%
#447920000000
0!
0%
#447925000000
1!
1%
#447930000000
0!
0%
#447935000000
1!
1%
#447940000000
0!
0%
#447945000000
1!
1%
#447950000000
0!
0%
#447955000000
1!
1%
#447960000000
0!
0%
#447965000000
1!
1%
#447970000000
0!
0%
#447975000000
1!
1%
#447980000000
0!
0%
#447985000000
1!
1%
#447990000000
0!
0%
#447995000000
1!
1%
#448000000000
0!
0%
#448005000000
1!
1%
#448010000000
0!
0%
#448015000000
1!
1%
#448020000000
0!
0%
#448025000000
1!
1%
#448030000000
0!
0%
#448035000000
1!
1%
#448040000000
0!
0%
#448045000000
1!
1%
#448050000000
0!
0%
#448055000000
1!
1%
#448060000000
0!
0%
#448065000000
1!
1%
#448070000000
0!
0%
#448075000000
1!
1%
#448080000000
0!
0%
#448085000000
1!
1%
#448090000000
0!
0%
#448095000000
1!
1%
#448100000000
0!
0%
#448105000000
1!
1%
#448110000000
0!
0%
#448115000000
1!
1%
#448120000000
0!
0%
#448125000000
1!
1%
#448130000000
0!
0%
#448135000000
1!
1%
#448140000000
0!
0%
#448145000000
1!
1%
#448150000000
0!
0%
#448155000000
1!
1%
#448160000000
0!
0%
#448165000000
1!
1%
#448170000000
0!
0%
#448175000000
1!
1%
#448180000000
0!
0%
#448185000000
1!
1%
#448190000000
0!
0%
#448195000000
1!
1%
#448200000000
0!
0%
#448205000000
1!
1%
#448210000000
0!
0%
#448215000000
1!
1%
#448220000000
0!
0%
#448225000000
1!
1%
#448230000000
0!
0%
#448235000000
1!
1%
#448240000000
0!
0%
#448245000000
1!
1%
#448250000000
0!
0%
#448255000000
1!
1%
#448260000000
0!
0%
#448265000000
1!
1%
#448270000000
0!
0%
#448275000000
1!
1%
#448280000000
0!
0%
#448285000000
1!
1%
#448290000000
0!
0%
#448295000000
1!
1%
#448300000000
0!
0%
#448305000000
1!
1%
#448310000000
0!
0%
#448315000000
1!
1%
#448320000000
0!
0%
#448325000000
1!
1%
#448330000000
0!
0%
#448335000000
1!
1%
#448340000000
0!
0%
#448345000000
1!
1%
#448350000000
0!
0%
#448355000000
1!
1%
#448360000000
0!
0%
#448365000000
1!
1%
#448370000000
0!
0%
#448375000000
1!
1%
#448380000000
0!
0%
#448385000000
1!
1%
#448390000000
0!
0%
#448395000000
1!
1%
#448400000000
0!
0%
#448405000000
1!
1%
#448410000000
0!
0%
#448415000000
1!
1%
#448420000000
0!
0%
#448425000000
1!
1%
#448430000000
0!
0%
#448435000000
1!
1%
#448440000000
0!
0%
#448445000000
1!
1%
#448450000000
0!
0%
#448455000000
1!
1%
#448460000000
0!
0%
#448465000000
1!
1%
#448470000000
0!
0%
#448475000000
1!
1%
#448480000000
0!
0%
#448485000000
1!
1%
#448490000000
0!
0%
#448495000000
1!
1%
#448500000000
0!
0%
#448505000000
1!
1%
#448510000000
0!
0%
#448515000000
1!
1%
#448520000000
0!
0%
#448525000000
1!
1%
#448530000000
0!
0%
#448535000000
1!
1%
#448540000000
0!
0%
#448545000000
1!
1%
#448550000000
0!
0%
#448555000000
1!
1%
#448560000000
0!
0%
#448565000000
1!
1%
#448570000000
0!
0%
#448575000000
1!
1%
#448580000000
0!
0%
#448585000000
1!
1%
#448590000000
0!
0%
#448595000000
1!
1%
#448600000000
0!
0%
#448605000000
1!
1%
#448610000000
0!
0%
#448615000000
1!
1%
#448620000000
0!
0%
#448625000000
1!
1%
#448630000000
0!
0%
#448635000000
1!
1%
#448640000000
0!
0%
#448645000000
1!
1%
#448650000000
0!
0%
#448655000000
1!
1%
#448660000000
0!
0%
#448665000000
1!
1%
#448670000000
0!
0%
#448675000000
1!
1%
#448680000000
0!
0%
#448685000000
1!
1%
#448690000000
0!
0%
#448695000000
1!
1%
#448700000000
0!
0%
#448705000000
1!
1%
#448710000000
0!
0%
#448715000000
1!
1%
#448720000000
0!
0%
#448725000000
1!
1%
#448730000000
0!
0%
#448735000000
1!
1%
#448740000000
0!
0%
#448745000000
1!
1%
#448750000000
0!
0%
#448755000000
1!
1%
#448760000000
0!
0%
#448765000000
1!
1%
#448770000000
0!
0%
#448775000000
1!
1%
#448780000000
0!
0%
#448785000000
1!
1%
#448790000000
0!
0%
#448795000000
1!
1%
#448800000000
0!
0%
#448805000000
1!
1%
#448810000000
0!
0%
#448815000000
1!
1%
#448820000000
0!
0%
#448825000000
1!
1%
#448830000000
0!
0%
#448835000000
1!
1%
#448840000000
0!
0%
#448845000000
1!
1%
#448850000000
0!
0%
#448855000000
1!
1%
#448860000000
0!
0%
#448865000000
1!
1%
#448870000000
0!
0%
#448875000000
1!
1%
#448880000000
0!
0%
#448885000000
1!
1%
#448890000000
0!
0%
#448895000000
1!
1%
#448900000000
0!
0%
#448905000000
1!
1%
#448910000000
0!
0%
#448915000000
1!
1%
#448920000000
0!
0%
#448925000000
1!
1%
#448930000000
0!
0%
#448935000000
1!
1%
#448940000000
0!
0%
#448945000000
1!
1%
#448950000000
0!
0%
#448955000000
1!
1%
#448960000000
0!
0%
#448965000000
1!
1%
#448970000000
0!
0%
#448975000000
1!
1%
#448980000000
0!
0%
#448985000000
1!
1%
#448990000000
0!
0%
#448995000000
1!
1%
#449000000000
0!
0%
#449005000000
1!
1%
#449010000000
0!
0%
#449015000000
1!
1%
#449020000000
0!
0%
#449025000000
1!
1%
#449030000000
0!
0%
#449035000000
1!
1%
#449040000000
0!
0%
#449045000000
1!
1%
#449050000000
0!
0%
#449055000000
1!
1%
#449060000000
0!
0%
#449065000000
1!
1%
#449070000000
0!
0%
#449075000000
1!
1%
#449080000000
0!
0%
#449085000000
1!
1%
#449090000000
0!
0%
#449095000000
1!
1%
#449100000000
0!
0%
#449105000000
1!
1%
#449110000000
0!
0%
#449115000000
1!
1%
#449120000000
0!
0%
#449125000000
1!
1%
#449130000000
0!
0%
#449135000000
1!
1%
#449140000000
0!
0%
#449145000000
1!
1%
#449150000000
0!
0%
#449155000000
1!
1%
#449160000000
0!
0%
#449165000000
1!
1%
#449170000000
0!
0%
#449175000000
1!
1%
#449180000000
0!
0%
#449185000000
1!
1%
#449190000000
0!
0%
#449195000000
1!
1%
#449200000000
0!
0%
#449205000000
1!
1%
#449210000000
0!
0%
#449215000000
1!
1%
#449220000000
0!
0%
#449225000000
1!
1%
#449230000000
0!
0%
#449235000000
1!
1%
#449240000000
0!
0%
#449245000000
1!
1%
#449250000000
0!
0%
#449255000000
1!
1%
#449260000000
0!
0%
#449265000000
1!
1%
#449270000000
0!
0%
#449275000000
1!
1%
#449280000000
0!
0%
#449285000000
1!
1%
#449290000000
0!
0%
#449295000000
1!
1%
#449300000000
0!
0%
#449305000000
1!
1%
#449310000000
0!
0%
#449315000000
1!
1%
#449320000000
0!
0%
#449325000000
1!
1%
#449330000000
0!
0%
#449335000000
1!
1%
#449340000000
0!
0%
#449345000000
1!
1%
#449350000000
0!
0%
#449355000000
1!
1%
#449360000000
0!
0%
#449365000000
1!
1%
#449370000000
0!
0%
#449375000000
1!
1%
#449380000000
0!
0%
#449385000000
1!
1%
#449390000000
0!
0%
#449395000000
1!
1%
#449400000000
0!
0%
#449405000000
1!
1%
#449410000000
0!
0%
#449415000000
1!
1%
#449420000000
0!
0%
#449425000000
1!
1%
#449430000000
0!
0%
#449435000000
1!
1%
#449440000000
0!
0%
#449445000000
1!
1%
#449450000000
0!
0%
#449455000000
1!
1%
#449460000000
0!
0%
#449465000000
1!
1%
#449470000000
0!
0%
#449475000000
1!
1%
#449480000000
0!
0%
#449485000000
1!
1%
#449490000000
0!
0%
#449495000000
1!
1%
#449500000000
0!
0%
#449505000000
1!
1%
#449510000000
0!
0%
#449515000000
1!
1%
#449520000000
0!
0%
#449525000000
1!
1%
#449530000000
0!
0%
#449535000000
1!
1%
#449540000000
0!
0%
#449545000000
1!
1%
#449550000000
0!
0%
#449555000000
1!
1%
#449560000000
0!
0%
#449565000000
1!
1%
#449570000000
0!
0%
#449575000000
1!
1%
#449580000000
0!
0%
#449585000000
1!
1%
#449590000000
0!
0%
#449595000000
1!
1%
#449600000000
0!
0%
#449605000000
1!
1%
#449610000000
0!
0%
#449615000000
1!
1%
#449620000000
0!
0%
#449625000000
1!
1%
#449630000000
0!
0%
#449635000000
1!
1%
#449640000000
0!
0%
#449645000000
1!
1%
#449650000000
0!
0%
#449655000000
1!
1%
#449660000000
0!
0%
#449665000000
1!
1%
#449670000000
0!
0%
#449675000000
1!
1%
#449680000000
0!
0%
#449685000000
1!
1%
#449690000000
0!
0%
#449695000000
1!
1%
#449700000000
0!
0%
#449705000000
1!
1%
#449710000000
0!
0%
#449715000000
1!
1%
#449720000000
0!
0%
#449725000000
1!
1%
#449730000000
0!
0%
#449735000000
1!
1%
#449740000000
0!
0%
#449745000000
1!
1%
#449750000000
0!
0%
#449755000000
1!
1%
#449760000000
0!
0%
#449765000000
1!
1%
#449770000000
0!
0%
#449775000000
1!
1%
#449780000000
0!
0%
#449785000000
1!
1%
#449790000000
0!
0%
#449795000000
1!
1%
#449800000000
0!
0%
#449805000000
1!
1%
#449810000000
0!
0%
#449815000000
1!
1%
#449820000000
0!
0%
#449825000000
1!
1%
#449830000000
0!
0%
#449835000000
1!
1%
#449840000000
0!
0%
#449845000000
1!
1%
#449850000000
0!
0%
#449855000000
1!
1%
#449860000000
0!
0%
#449865000000
1!
1%
#449870000000
0!
0%
#449875000000
1!
1%
#449880000000
0!
0%
#449885000000
1!
1%
#449890000000
0!
0%
#449895000000
1!
1%
#449900000000
0!
0%
#449905000000
1!
1%
#449910000000
0!
0%
#449915000000
1!
1%
#449920000000
0!
0%
#449925000000
1!
1%
#449930000000
0!
0%
#449935000000
1!
1%
#449940000000
0!
0%
#449945000000
1!
1%
#449950000000
0!
0%
#449955000000
1!
1%
#449960000000
0!
0%
#449965000000
1!
1%
#449970000000
0!
0%
#449975000000
1!
1%
#449980000000
0!
0%
#449985000000
1!
1%
#449990000000
0!
0%
#449995000000
1!
1%
#450000000000
0!
0%
#450005000000
1!
1%
#450010000000
0!
0%
#450015000000
1!
1%
#450020000000
0!
0%
#450025000000
1!
1%
#450030000000
0!
0%
#450035000000
1!
1%
#450040000000
0!
0%
#450045000000
1!
1%
#450050000000
0!
0%
#450055000000
1!
1%
#450060000000
0!
0%
#450065000000
1!
1%
#450070000000
0!
0%
#450075000000
1!
1%
#450080000000
0!
0%
#450085000000
1!
1%
#450090000000
0!
0%
#450095000000
1!
1%
#450100000000
0!
0%
#450105000000
1!
1%
#450110000000
0!
0%
#450115000000
1!
1%
#450120000000
0!
0%
#450125000000
1!
1%
#450130000000
0!
0%
#450135000000
1!
1%
#450140000000
0!
0%
#450145000000
1!
1%
#450150000000
0!
0%
#450155000000
1!
1%
#450160000000
0!
0%
#450165000000
1!
1%
#450170000000
0!
0%
#450175000000
1!
1%
#450180000000
0!
0%
#450185000000
1!
1%
#450190000000
0!
0%
#450195000000
1!
1%
#450200000000
0!
0%
#450205000000
1!
1%
#450210000000
0!
0%
#450215000000
1!
1%
#450220000000
0!
0%
#450225000000
1!
1%
#450230000000
0!
0%
#450235000000
1!
1%
#450240000000
0!
0%
#450245000000
1!
1%
#450250000000
0!
0%
#450255000000
1!
1%
#450260000000
0!
0%
#450265000000
1!
1%
#450270000000
0!
0%
#450275000000
1!
1%
#450280000000
0!
0%
#450285000000
1!
1%
#450290000000
0!
0%
#450295000000
1!
1%
#450300000000
0!
0%
#450305000000
1!
1%
#450310000000
0!
0%
#450315000000
1!
1%
#450320000000
0!
0%
#450325000000
1!
1%
#450330000000
0!
0%
#450335000000
1!
1%
#450340000000
0!
0%
#450345000000
1!
1%
#450350000000
0!
0%
#450355000000
1!
1%
#450360000000
0!
0%
#450365000000
1!
1%
#450370000000
0!
0%
#450375000000
1!
1%
#450380000000
0!
0%
#450385000000
1!
1%
#450390000000
0!
0%
#450395000000
1!
1%
#450400000000
0!
0%
#450405000000
1!
1%
#450410000000
0!
0%
#450415000000
1!
1%
#450420000000
0!
0%
#450425000000
1!
1%
#450430000000
0!
0%
#450435000000
1!
1%
#450440000000
0!
0%
#450445000000
1!
1%
#450450000000
0!
0%
#450455000000
1!
1%
#450460000000
0!
0%
#450465000000
1!
1%
#450470000000
0!
0%
#450475000000
1!
1%
#450480000000
0!
0%
#450485000000
1!
1%
#450490000000
0!
0%
#450495000000
1!
1%
#450500000000
0!
0%
#450505000000
1!
1%
#450510000000
0!
0%
#450515000000
1!
1%
#450520000000
0!
0%
#450525000000
1!
1%
#450530000000
0!
0%
#450535000000
1!
1%
#450540000000
0!
0%
#450545000000
1!
1%
#450550000000
0!
0%
#450555000000
1!
1%
#450560000000
0!
0%
#450565000000
1!
1%
#450570000000
0!
0%
#450575000000
1!
1%
#450580000000
0!
0%
#450585000000
1!
1%
#450590000000
0!
0%
#450595000000
1!
1%
#450600000000
0!
0%
#450605000000
1!
1%
#450610000000
0!
0%
#450615000000
1!
1%
#450620000000
0!
0%
#450625000000
1!
1%
#450630000000
0!
0%
#450635000000
1!
1%
#450640000000
0!
0%
#450645000000
1!
1%
#450650000000
0!
0%
#450655000000
1!
1%
#450660000000
0!
0%
#450665000000
1!
1%
#450670000000
0!
0%
#450675000000
1!
1%
#450680000000
0!
0%
#450685000000
1!
1%
#450690000000
0!
0%
#450695000000
1!
1%
#450700000000
0!
0%
#450705000000
1!
1%
#450710000000
0!
0%
#450715000000
1!
1%
#450720000000
0!
0%
#450725000000
1!
1%
#450730000000
0!
0%
#450735000000
1!
1%
#450740000000
0!
0%
#450745000000
1!
1%
#450750000000
0!
0%
#450755000000
1!
1%
#450760000000
0!
0%
#450765000000
1!
1%
#450770000000
0!
0%
#450775000000
1!
1%
#450780000000
0!
0%
#450785000000
1!
1%
#450790000000
0!
0%
#450795000000
1!
1%
#450800000000
0!
0%
#450805000000
1!
1%
#450810000000
0!
0%
#450815000000
1!
1%
#450820000000
0!
0%
#450825000000
1!
1%
#450830000000
0!
0%
#450835000000
1!
1%
#450840000000
0!
0%
#450845000000
1!
1%
#450850000000
0!
0%
#450855000000
1!
1%
#450860000000
0!
0%
#450865000000
1!
1%
#450870000000
0!
0%
#450875000000
1!
1%
#450880000000
0!
0%
#450885000000
1!
1%
#450890000000
0!
0%
#450895000000
1!
1%
#450900000000
0!
0%
#450905000000
1!
1%
#450910000000
0!
0%
#450915000000
1!
1%
#450920000000
0!
0%
#450925000000
1!
1%
#450930000000
0!
0%
#450935000000
1!
1%
#450940000000
0!
0%
#450945000000
1!
1%
#450950000000
0!
0%
#450955000000
1!
1%
#450960000000
0!
0%
#450965000000
1!
1%
#450970000000
0!
0%
#450975000000
1!
1%
#450980000000
0!
0%
#450985000000
1!
1%
#450990000000
0!
0%
#450995000000
1!
1%
#451000000000
0!
0%
#451005000000
1!
1%
#451010000000
0!
0%
#451015000000
1!
1%
#451020000000
0!
0%
#451025000000
1!
1%
#451030000000
0!
0%
#451035000000
1!
1%
#451040000000
0!
0%
#451045000000
1!
1%
#451050000000
0!
0%
#451055000000
1!
1%
#451060000000
0!
0%
#451065000000
1!
1%
#451070000000
0!
0%
#451075000000
1!
1%
#451080000000
0!
0%
#451085000000
1!
1%
#451090000000
0!
0%
#451095000000
1!
1%
#451100000000
0!
0%
#451105000000
1!
1%
#451110000000
0!
0%
#451115000000
1!
1%
#451120000000
0!
0%
#451125000000
1!
1%
#451130000000
0!
0%
#451135000000
1!
1%
#451140000000
0!
0%
#451145000000
1!
1%
#451150000000
0!
0%
#451155000000
1!
1%
#451160000000
0!
0%
#451165000000
1!
1%
#451170000000
0!
0%
#451175000000
1!
1%
#451180000000
0!
0%
#451185000000
1!
1%
#451190000000
0!
0%
#451195000000
1!
1%
#451200000000
0!
0%
#451205000000
1!
1%
#451210000000
0!
0%
#451215000000
1!
1%
#451220000000
0!
0%
#451225000000
1!
1%
#451230000000
0!
0%
#451235000000
1!
1%
#451240000000
0!
0%
#451245000000
1!
1%
#451250000000
0!
0%
#451255000000
1!
1%
#451260000000
0!
0%
#451265000000
1!
1%
#451270000000
0!
0%
#451275000000
1!
1%
#451280000000
0!
0%
#451285000000
1!
1%
#451290000000
0!
0%
#451295000000
1!
1%
#451300000000
0!
0%
#451305000000
1!
1%
#451310000000
0!
0%
#451315000000
1!
1%
#451320000000
0!
0%
#451325000000
1!
1%
#451330000000
0!
0%
#451335000000
1!
1%
#451340000000
0!
0%
#451345000000
1!
1%
#451350000000
0!
0%
#451355000000
1!
1%
#451360000000
0!
0%
#451365000000
1!
1%
#451370000000
0!
0%
#451375000000
1!
1%
#451380000000
0!
0%
#451385000000
1!
1%
#451390000000
0!
0%
#451395000000
1!
1%
#451400000000
0!
0%
#451405000000
1!
1%
#451410000000
0!
0%
#451415000000
1!
1%
#451420000000
0!
0%
#451425000000
1!
1%
#451430000000
0!
0%
#451435000000
1!
1%
#451440000000
0!
0%
#451445000000
1!
1%
#451450000000
0!
0%
#451455000000
1!
1%
#451460000000
0!
0%
#451465000000
1!
1%
#451470000000
0!
0%
#451475000000
1!
1%
#451480000000
0!
0%
#451485000000
1!
1%
#451490000000
0!
0%
#451495000000
1!
1%
#451500000000
0!
0%
#451505000000
1!
1%
#451510000000
0!
0%
#451515000000
1!
1%
#451520000000
0!
0%
#451525000000
1!
1%
#451530000000
0!
0%
#451535000000
1!
1%
#451540000000
0!
0%
#451545000000
1!
1%
#451550000000
0!
0%
#451555000000
1!
1%
#451560000000
0!
0%
#451565000000
1!
1%
#451570000000
0!
0%
#451575000000
1!
1%
#451580000000
0!
0%
#451585000000
1!
1%
#451590000000
0!
0%
#451595000000
1!
1%
#451600000000
0!
0%
#451605000000
1!
1%
#451610000000
0!
0%
#451615000000
1!
1%
#451620000000
0!
0%
#451625000000
1!
1%
#451630000000
0!
0%
#451635000000
1!
1%
#451640000000
0!
0%
#451645000000
1!
1%
#451650000000
0!
0%
#451655000000
1!
1%
#451660000000
0!
0%
#451665000000
1!
1%
#451670000000
0!
0%
#451675000000
1!
1%
#451680000000
0!
0%
#451685000000
1!
1%
#451690000000
0!
0%
#451695000000
1!
1%
#451700000000
0!
0%
#451705000000
1!
1%
#451710000000
0!
0%
#451715000000
1!
1%
#451720000000
0!
0%
#451725000000
1!
1%
#451730000000
0!
0%
#451735000000
1!
1%
#451740000000
0!
0%
#451745000000
1!
1%
#451750000000
0!
0%
#451755000000
1!
1%
#451760000000
0!
0%
#451765000000
1!
1%
#451770000000
0!
0%
#451775000000
1!
1%
#451780000000
0!
0%
#451785000000
1!
1%
#451790000000
0!
0%
#451795000000
1!
1%
#451800000000
0!
0%
#451805000000
1!
1%
#451810000000
0!
0%
#451815000000
1!
1%
#451820000000
0!
0%
#451825000000
1!
1%
#451830000000
0!
0%
#451835000000
1!
1%
#451840000000
0!
0%
#451845000000
1!
1%
#451850000000
0!
0%
#451855000000
1!
1%
#451860000000
0!
0%
#451865000000
1!
1%
#451870000000
0!
0%
#451875000000
1!
1%
#451880000000
0!
0%
#451885000000
1!
1%
#451890000000
0!
0%
#451895000000
1!
1%
#451900000000
0!
0%
#451905000000
1!
1%
#451910000000
0!
0%
#451915000000
1!
1%
#451920000000
0!
0%
#451925000000
1!
1%
#451930000000
0!
0%
#451935000000
1!
1%
#451940000000
0!
0%
#451945000000
1!
1%
#451950000000
0!
0%
#451955000000
1!
1%
#451960000000
0!
0%
#451965000000
1!
1%
#451970000000
0!
0%
#451975000000
1!
1%
#451980000000
0!
0%
#451985000000
1!
1%
#451990000000
0!
0%
#451995000000
1!
1%
#452000000000
0!
0%
#452005000000
1!
1%
#452010000000
0!
0%
#452015000000
1!
1%
#452020000000
0!
0%
#452025000000
1!
1%
#452030000000
0!
0%
#452035000000
1!
1%
#452040000000
0!
0%
#452045000000
1!
1%
#452050000000
0!
0%
#452055000000
1!
1%
#452060000000
0!
0%
#452065000000
1!
1%
#452070000000
0!
0%
#452075000000
1!
1%
#452080000000
0!
0%
#452085000000
1!
1%
#452090000000
0!
0%
#452095000000
1!
1%
#452100000000
0!
0%
#452105000000
1!
1%
#452110000000
0!
0%
#452115000000
1!
1%
#452120000000
0!
0%
#452125000000
1!
1%
#452130000000
0!
0%
#452135000000
1!
1%
#452140000000
0!
0%
#452145000000
1!
1%
#452150000000
0!
0%
#452155000000
1!
1%
#452160000000
0!
0%
#452165000000
1!
1%
#452170000000
0!
0%
#452175000000
1!
1%
#452180000000
0!
0%
#452185000000
1!
1%
#452190000000
0!
0%
#452195000000
1!
1%
#452200000000
0!
0%
#452205000000
1!
1%
#452210000000
0!
0%
#452215000000
1!
1%
#452220000000
0!
0%
#452225000000
1!
1%
#452230000000
0!
0%
#452235000000
1!
1%
#452240000000
0!
0%
#452245000000
1!
1%
#452250000000
0!
0%
#452255000000
1!
1%
#452260000000
0!
0%
#452265000000
1!
1%
#452270000000
0!
0%
#452275000000
1!
1%
#452280000000
0!
0%
#452285000000
1!
1%
#452290000000
0!
0%
#452295000000
1!
1%
#452300000000
0!
0%
#452305000000
1!
1%
#452310000000
0!
0%
#452315000000
1!
1%
#452320000000
0!
0%
#452325000000
1!
1%
#452330000000
0!
0%
#452335000000
1!
1%
#452340000000
0!
0%
#452345000000
1!
1%
#452350000000
0!
0%
#452355000000
1!
1%
#452360000000
0!
0%
#452365000000
1!
1%
#452370000000
0!
0%
#452375000000
1!
1%
#452380000000
0!
0%
#452385000000
1!
1%
#452390000000
0!
0%
#452395000000
1!
1%
#452400000000
0!
0%
#452405000000
1!
1%
#452410000000
0!
0%
#452415000000
1!
1%
#452420000000
0!
0%
#452425000000
1!
1%
#452430000000
0!
0%
#452435000000
1!
1%
#452440000000
0!
0%
#452445000000
1!
1%
#452450000000
0!
0%
#452455000000
1!
1%
#452460000000
0!
0%
#452465000000
1!
1%
#452470000000
0!
0%
#452475000000
1!
1%
#452480000000
0!
0%
#452485000000
1!
1%
#452490000000
0!
0%
#452495000000
1!
1%
#452500000000
0!
0%
#452505000000
1!
1%
#452510000000
0!
0%
#452515000000
1!
1%
#452520000000
0!
0%
#452525000000
1!
1%
#452530000000
0!
0%
#452535000000
1!
1%
#452540000000
0!
0%
#452545000000
1!
1%
#452550000000
0!
0%
#452555000000
1!
1%
#452560000000
0!
0%
#452565000000
1!
1%
#452570000000
0!
0%
#452575000000
1!
1%
#452580000000
0!
0%
#452585000000
1!
1%
#452590000000
0!
0%
#452595000000
1!
1%
#452600000000
0!
0%
#452605000000
1!
1%
#452610000000
0!
0%
#452615000000
1!
1%
#452620000000
0!
0%
#452625000000
1!
1%
#452630000000
0!
0%
#452635000000
1!
1%
#452640000000
0!
0%
#452645000000
1!
1%
#452650000000
0!
0%
#452655000000
1!
1%
#452660000000
0!
0%
#452665000000
1!
1%
#452670000000
0!
0%
#452675000000
1!
1%
#452680000000
0!
0%
#452685000000
1!
1%
#452690000000
0!
0%
#452695000000
1!
1%
#452700000000
0!
0%
#452705000000
1!
1%
#452710000000
0!
0%
#452715000000
1!
1%
#452720000000
0!
0%
#452725000000
1!
1%
#452730000000
0!
0%
#452735000000
1!
1%
#452740000000
0!
0%
#452745000000
1!
1%
#452750000000
0!
0%
#452755000000
1!
1%
#452760000000
0!
0%
#452765000000
1!
1%
#452770000000
0!
0%
#452775000000
1!
1%
#452780000000
0!
0%
#452785000000
1!
1%
#452790000000
0!
0%
#452795000000
1!
1%
#452800000000
0!
0%
#452805000000
1!
1%
#452810000000
0!
0%
#452815000000
1!
1%
#452820000000
0!
0%
#452825000000
1!
1%
#452830000000
0!
0%
#452835000000
1!
1%
#452840000000
0!
0%
#452845000000
1!
1%
#452850000000
0!
0%
#452855000000
1!
1%
#452860000000
0!
0%
#452865000000
1!
1%
#452870000000
0!
0%
#452875000000
1!
1%
#452880000000
0!
0%
#452885000000
1!
1%
#452890000000
0!
0%
#452895000000
1!
1%
#452900000000
0!
0%
#452905000000
1!
1%
#452910000000
0!
0%
#452915000000
1!
1%
#452920000000
0!
0%
#452925000000
1!
1%
#452930000000
0!
0%
#452935000000
1!
1%
#452940000000
0!
0%
#452945000000
1!
1%
#452950000000
0!
0%
#452955000000
1!
1%
#452960000000
0!
0%
#452965000000
1!
1%
#452970000000
0!
0%
#452975000000
1!
1%
#452980000000
0!
0%
#452985000000
1!
1%
#452990000000
0!
0%
#452995000000
1!
1%
#453000000000
0!
0%
#453005000000
1!
1%
#453010000000
0!
0%
#453015000000
1!
1%
#453020000000
0!
0%
#453025000000
1!
1%
#453030000000
0!
0%
#453035000000
1!
1%
#453040000000
0!
0%
#453045000000
1!
1%
#453050000000
0!
0%
#453055000000
1!
1%
#453060000000
0!
0%
#453065000000
1!
1%
#453070000000
0!
0%
#453075000000
1!
1%
#453080000000
0!
0%
#453085000000
1!
1%
#453090000000
0!
0%
#453095000000
1!
1%
#453100000000
0!
0%
#453105000000
1!
1%
#453110000000
0!
0%
#453115000000
1!
1%
#453120000000
0!
0%
#453125000000
1!
1%
#453130000000
0!
0%
#453135000000
1!
1%
#453140000000
0!
0%
#453145000000
1!
1%
#453150000000
0!
0%
#453155000000
1!
1%
#453160000000
0!
0%
#453165000000
1!
1%
#453170000000
0!
0%
#453175000000
1!
1%
#453180000000
0!
0%
#453185000000
1!
1%
#453190000000
0!
0%
#453195000000
1!
1%
#453200000000
0!
0%
#453205000000
1!
1%
#453210000000
0!
0%
#453215000000
1!
1%
#453220000000
0!
0%
#453225000000
1!
1%
#453230000000
0!
0%
#453235000000
1!
1%
#453240000000
0!
0%
#453245000000
1!
1%
#453250000000
0!
0%
#453255000000
1!
1%
#453260000000
0!
0%
#453265000000
1!
1%
#453270000000
0!
0%
#453275000000
1!
1%
#453280000000
0!
0%
#453285000000
1!
1%
#453290000000
0!
0%
#453295000000
1!
1%
#453300000000
0!
0%
#453305000000
1!
1%
#453310000000
0!
0%
#453315000000
1!
1%
#453320000000
0!
0%
#453325000000
1!
1%
#453330000000
0!
0%
#453335000000
1!
1%
#453340000000
0!
0%
#453345000000
1!
1%
#453350000000
0!
0%
#453355000000
1!
1%
#453360000000
0!
0%
#453365000000
1!
1%
#453370000000
0!
0%
#453375000000
1!
1%
#453380000000
0!
0%
#453385000000
1!
1%
#453390000000
0!
0%
#453395000000
1!
1%
#453400000000
0!
0%
#453405000000
1!
1%
#453410000000
0!
0%
#453415000000
1!
1%
#453420000000
0!
0%
#453425000000
1!
1%
#453430000000
0!
0%
#453435000000
1!
1%
#453440000000
0!
0%
#453445000000
1!
1%
#453450000000
0!
0%
#453455000000
1!
1%
#453460000000
0!
0%
#453465000000
1!
1%
#453470000000
0!
0%
#453475000000
1!
1%
#453480000000
0!
0%
#453485000000
1!
1%
#453490000000
0!
0%
#453495000000
1!
1%
#453500000000
0!
0%
#453505000000
1!
1%
#453510000000
0!
0%
#453515000000
1!
1%
#453520000000
0!
0%
#453525000000
1!
1%
#453530000000
0!
0%
#453535000000
1!
1%
#453540000000
0!
0%
#453545000000
1!
1%
#453550000000
0!
0%
#453555000000
1!
1%
#453560000000
0!
0%
#453565000000
1!
1%
#453570000000
0!
0%
#453575000000
1!
1%
#453580000000
0!
0%
#453585000000
1!
1%
#453590000000
0!
0%
#453595000000
1!
1%
#453600000000
0!
0%
#453605000000
1!
1%
#453610000000
0!
0%
#453615000000
1!
1%
#453620000000
0!
0%
#453625000000
1!
1%
#453630000000
0!
0%
#453635000000
1!
1%
#453640000000
0!
0%
#453645000000
1!
1%
#453650000000
0!
0%
#453655000000
1!
1%
#453660000000
0!
0%
#453665000000
1!
1%
#453670000000
0!
0%
#453675000000
1!
1%
#453680000000
0!
0%
#453685000000
1!
1%
#453690000000
0!
0%
#453695000000
1!
1%
#453700000000
0!
0%
#453705000000
1!
1%
#453710000000
0!
0%
#453715000000
1!
1%
#453720000000
0!
0%
#453725000000
1!
1%
#453730000000
0!
0%
#453735000000
1!
1%
#453740000000
0!
0%
#453745000000
1!
1%
#453750000000
0!
0%
#453755000000
1!
1%
#453760000000
0!
0%
#453765000000
1!
1%
#453770000000
0!
0%
#453775000000
1!
1%
#453780000000
0!
0%
#453785000000
1!
1%
#453790000000
0!
0%
#453795000000
1!
1%
#453800000000
0!
0%
#453805000000
1!
1%
#453810000000
0!
0%
#453815000000
1!
1%
#453820000000
0!
0%
#453825000000
1!
1%
#453830000000
0!
0%
#453835000000
1!
1%
#453840000000
0!
0%
#453845000000
1!
1%
#453850000000
0!
0%
#453855000000
1!
1%
#453860000000
0!
0%
#453865000000
1!
1%
#453870000000
0!
0%
#453875000000
1!
1%
#453880000000
0!
0%
#453885000000
1!
1%
#453890000000
0!
0%
#453895000000
1!
1%
#453900000000
0!
0%
#453905000000
1!
1%
#453910000000
0!
0%
#453915000000
1!
1%
#453920000000
0!
0%
#453925000000
1!
1%
#453930000000
0!
0%
#453935000000
1!
1%
#453940000000
0!
0%
#453945000000
1!
1%
#453950000000
0!
0%
#453955000000
1!
1%
#453960000000
0!
0%
#453965000000
1!
1%
#453970000000
0!
0%
#453975000000
1!
1%
#453980000000
0!
0%
#453985000000
1!
1%
#453990000000
0!
0%
#453995000000
1!
1%
#454000000000
0!
0%
#454005000000
1!
1%
#454010000000
0!
0%
#454015000000
1!
1%
#454020000000
0!
0%
#454025000000
1!
1%
#454030000000
0!
0%
#454035000000
1!
1%
#454040000000
0!
0%
#454045000000
1!
1%
#454050000000
0!
0%
#454055000000
1!
1%
#454060000000
0!
0%
#454065000000
1!
1%
#454070000000
0!
0%
#454075000000
1!
1%
#454080000000
0!
0%
#454085000000
1!
1%
#454090000000
0!
0%
#454095000000
1!
1%
#454100000000
0!
0%
#454105000000
1!
1%
#454110000000
0!
0%
#454115000000
1!
1%
#454120000000
0!
0%
#454125000000
1!
1%
#454130000000
0!
0%
#454135000000
1!
1%
#454140000000
0!
0%
#454145000000
1!
1%
#454150000000
0!
0%
#454155000000
1!
1%
#454160000000
0!
0%
#454165000000
1!
1%
#454170000000
0!
0%
#454175000000
1!
1%
#454180000000
0!
0%
#454185000000
1!
1%
#454190000000
0!
0%
#454195000000
1!
1%
#454200000000
0!
0%
#454205000000
1!
1%
#454210000000
0!
0%
#454215000000
1!
1%
#454220000000
0!
0%
#454225000000
1!
1%
#454230000000
0!
0%
#454235000000
1!
1%
#454240000000
0!
0%
#454245000000
1!
1%
#454250000000
0!
0%
#454255000000
1!
1%
#454260000000
0!
0%
#454265000000
1!
1%
#454270000000
0!
0%
#454275000000
1!
1%
#454280000000
0!
0%
#454285000000
1!
1%
#454290000000
0!
0%
#454295000000
1!
1%
#454300000000
0!
0%
#454305000000
1!
1%
#454310000000
0!
0%
#454315000000
1!
1%
#454320000000
0!
0%
#454325000000
1!
1%
#454330000000
0!
0%
#454335000000
1!
1%
#454340000000
0!
0%
#454345000000
1!
1%
#454350000000
0!
0%
#454355000000
1!
1%
#454360000000
0!
0%
#454365000000
1!
1%
#454370000000
0!
0%
#454375000000
1!
1%
#454380000000
0!
0%
#454385000000
1!
1%
#454390000000
0!
0%
#454395000000
1!
1%
#454400000000
0!
0%
#454405000000
1!
1%
#454410000000
0!
0%
#454415000000
1!
1%
#454420000000
0!
0%
#454425000000
1!
1%
#454430000000
0!
0%
#454435000000
1!
1%
#454440000000
0!
0%
#454445000000
1!
1%
#454450000000
0!
0%
#454455000000
1!
1%
#454460000000
0!
0%
#454465000000
1!
1%
#454470000000
0!
0%
#454475000000
1!
1%
#454480000000
0!
0%
#454485000000
1!
1%
#454490000000
0!
0%
#454495000000
1!
1%
#454500000000
0!
0%
#454505000000
1!
1%
#454510000000
0!
0%
#454515000000
1!
1%
#454520000000
0!
0%
#454525000000
1!
1%
#454530000000
0!
0%
#454535000000
1!
1%
#454540000000
0!
0%
#454545000000
1!
1%
#454550000000
0!
0%
#454555000000
1!
1%
#454560000000
0!
0%
#454565000000
1!
1%
#454570000000
0!
0%
#454575000000
1!
1%
#454580000000
0!
0%
#454585000000
1!
1%
#454590000000
0!
0%
#454595000000
1!
1%
#454600000000
0!
0%
#454605000000
1!
1%
#454610000000
0!
0%
#454615000000
1!
1%
#454620000000
0!
0%
#454625000000
1!
1%
#454630000000
0!
0%
#454635000000
1!
1%
#454640000000
0!
0%
#454645000000
1!
1%
#454650000000
0!
0%
#454655000000
1!
1%
#454660000000
0!
0%
#454665000000
1!
1%
#454670000000
0!
0%
#454675000000
1!
1%
#454680000000
0!
0%
#454685000000
1!
1%
#454690000000
0!
0%
#454695000000
1!
1%
#454700000000
0!
0%
#454705000000
1!
1%
#454710000000
0!
0%
#454715000000
1!
1%
#454720000000
0!
0%
#454725000000
1!
1%
#454730000000
0!
0%
#454735000000
1!
1%
#454740000000
0!
0%
#454745000000
1!
1%
#454750000000
0!
0%
#454755000000
1!
1%
#454760000000
0!
0%
#454765000000
1!
1%
#454770000000
0!
0%
#454775000000
1!
1%
#454780000000
0!
0%
#454785000000
1!
1%
#454790000000
0!
0%
#454795000000
1!
1%
#454800000000
0!
0%
#454805000000
1!
1%
#454810000000
0!
0%
#454815000000
1!
1%
#454820000000
0!
0%
#454825000000
1!
1%
#454830000000
0!
0%
#454835000000
1!
1%
#454840000000
0!
0%
#454845000000
1!
1%
#454850000000
0!
0%
#454855000000
1!
1%
#454860000000
0!
0%
#454865000000
1!
1%
#454870000000
0!
0%
#454875000000
1!
1%
#454880000000
0!
0%
#454885000000
1!
1%
#454890000000
0!
0%
#454895000000
1!
1%
#454900000000
0!
0%
#454905000000
1!
1%
#454910000000
0!
0%
#454915000000
1!
1%
#454920000000
0!
0%
#454925000000
1!
1%
#454930000000
0!
0%
#454935000000
1!
1%
#454940000000
0!
0%
#454945000000
1!
1%
#454950000000
0!
0%
#454955000000
1!
1%
#454960000000
0!
0%
#454965000000
1!
1%
#454970000000
0!
0%
#454975000000
1!
1%
#454980000000
0!
0%
#454985000000
1!
1%
#454990000000
0!
0%
#454995000000
1!
1%
#455000000000
0!
0%
#455005000000
1!
1%
#455010000000
0!
0%
#455015000000
1!
1%
#455020000000
0!
0%
#455025000000
1!
1%
#455030000000
0!
0%
#455035000000
1!
1%
#455040000000
0!
0%
#455045000000
1!
1%
#455050000000
0!
0%
#455055000000
1!
1%
#455060000000
0!
0%
#455065000000
1!
1%
#455070000000
0!
0%
#455075000000
1!
1%
#455080000000
0!
0%
#455085000000
1!
1%
#455090000000
0!
0%
#455095000000
1!
1%
#455100000000
0!
0%
#455105000000
1!
1%
#455110000000
0!
0%
#455115000000
1!
1%
#455120000000
0!
0%
#455125000000
1!
1%
#455130000000
0!
0%
#455135000000
1!
1%
#455140000000
0!
0%
#455145000000
1!
1%
#455150000000
0!
0%
#455155000000
1!
1%
#455160000000
0!
0%
#455165000000
1!
1%
#455170000000
0!
0%
#455175000000
1!
1%
#455180000000
0!
0%
#455185000000
1!
1%
#455190000000
0!
0%
#455195000000
1!
1%
#455200000000
0!
0%
#455205000000
1!
1%
#455210000000
0!
0%
#455215000000
1!
1%
#455220000000
0!
0%
#455225000000
1!
1%
#455230000000
0!
0%
#455235000000
1!
1%
#455240000000
0!
0%
#455245000000
1!
1%
#455250000000
0!
0%
#455255000000
1!
1%
#455260000000
0!
0%
#455265000000
1!
1%
#455270000000
0!
0%
#455275000000
1!
1%
#455280000000
0!
0%
#455285000000
1!
1%
#455290000000
0!
0%
#455295000000
1!
1%
#455300000000
0!
0%
#455305000000
1!
1%
#455310000000
0!
0%
#455315000000
1!
1%
#455320000000
0!
0%
#455325000000
1!
1%
#455330000000
0!
0%
#455335000000
1!
1%
#455340000000
0!
0%
#455345000000
1!
1%
#455350000000
0!
0%
#455355000000
1!
1%
#455360000000
0!
0%
#455365000000
1!
1%
#455370000000
0!
0%
#455375000000
1!
1%
#455380000000
0!
0%
#455385000000
1!
1%
#455390000000
0!
0%
#455395000000
1!
1%
#455400000000
0!
0%
#455405000000
1!
1%
#455410000000
0!
0%
#455415000000
1!
1%
#455420000000
0!
0%
#455425000000
1!
1%
#455430000000
0!
0%
#455435000000
1!
1%
#455440000000
0!
0%
#455445000000
1!
1%
#455450000000
0!
0%
#455455000000
1!
1%
#455460000000
0!
0%
#455465000000
1!
1%
#455470000000
0!
0%
#455475000000
1!
1%
#455480000000
0!
0%
#455485000000
1!
1%
#455490000000
0!
0%
#455495000000
1!
1%
#455500000000
0!
0%
#455505000000
1!
1%
#455510000000
0!
0%
#455515000000
1!
1%
#455520000000
0!
0%
#455525000000
1!
1%
#455530000000
0!
0%
#455535000000
1!
1%
#455540000000
0!
0%
#455545000000
1!
1%
#455550000000
0!
0%
#455555000000
1!
1%
#455560000000
0!
0%
#455565000000
1!
1%
#455570000000
0!
0%
#455575000000
1!
1%
#455580000000
0!
0%
#455585000000
1!
1%
#455590000000
0!
0%
#455595000000
1!
1%
#455600000000
0!
0%
#455605000000
1!
1%
#455610000000
0!
0%
#455615000000
1!
1%
#455620000000
0!
0%
#455625000000
1!
1%
#455630000000
0!
0%
#455635000000
1!
1%
#455640000000
0!
0%
#455645000000
1!
1%
#455650000000
0!
0%
#455655000000
1!
1%
#455660000000
0!
0%
#455665000000
1!
1%
#455670000000
0!
0%
#455675000000
1!
1%
#455680000000
0!
0%
#455685000000
1!
1%
#455690000000
0!
0%
#455695000000
1!
1%
#455700000000
0!
0%
#455705000000
1!
1%
#455710000000
0!
0%
#455715000000
1!
1%
#455720000000
0!
0%
#455725000000
1!
1%
#455730000000
0!
0%
#455735000000
1!
1%
#455740000000
0!
0%
#455745000000
1!
1%
#455750000000
0!
0%
#455755000000
1!
1%
#455760000000
0!
0%
#455765000000
1!
1%
#455770000000
0!
0%
#455775000000
1!
1%
#455780000000
0!
0%
#455785000000
1!
1%
#455790000000
0!
0%
#455795000000
1!
1%
#455800000000
0!
0%
#455805000000
1!
1%
#455810000000
0!
0%
#455815000000
1!
1%
#455820000000
0!
0%
#455825000000
1!
1%
#455830000000
0!
0%
#455835000000
1!
1%
#455840000000
0!
0%
#455845000000
1!
1%
#455850000000
0!
0%
#455855000000
1!
1%
#455860000000
0!
0%
#455865000000
1!
1%
#455870000000
0!
0%
#455875000000
1!
1%
#455880000000
0!
0%
#455885000000
1!
1%
#455890000000
0!
0%
#455895000000
1!
1%
#455900000000
0!
0%
#455905000000
1!
1%
#455910000000
0!
0%
#455915000000
1!
1%
#455920000000
0!
0%
#455925000000
1!
1%
#455930000000
0!
0%
#455935000000
1!
1%
#455940000000
0!
0%
#455945000000
1!
1%
#455950000000
0!
0%
#455955000000
1!
1%
#455960000000
0!
0%
#455965000000
1!
1%
#455970000000
0!
0%
#455975000000
1!
1%
#455980000000
0!
0%
#455985000000
1!
1%
#455990000000
0!
0%
#455995000000
1!
1%
#456000000000
0!
0%
#456005000000
1!
1%
#456010000000
0!
0%
#456015000000
1!
1%
#456020000000
0!
0%
#456025000000
1!
1%
#456030000000
0!
0%
#456035000000
1!
1%
#456040000000
0!
0%
#456045000000
1!
1%
#456050000000
0!
0%
#456055000000
1!
1%
#456060000000
0!
0%
#456065000000
1!
1%
#456070000000
0!
0%
#456075000000
1!
1%
#456080000000
0!
0%
#456085000000
1!
1%
#456090000000
0!
0%
#456095000000
1!
1%
#456100000000
0!
0%
#456105000000
1!
1%
#456110000000
0!
0%
#456115000000
1!
1%
#456120000000
0!
0%
#456125000000
1!
1%
#456130000000
0!
0%
#456135000000
1!
1%
#456140000000
0!
0%
#456145000000
1!
1%
#456150000000
0!
0%
#456155000000
1!
1%
#456160000000
0!
0%
#456165000000
1!
1%
#456170000000
0!
0%
#456175000000
1!
1%
#456180000000
0!
0%
#456185000000
1!
1%
#456190000000
0!
0%
#456195000000
1!
1%
#456200000000
0!
0%
#456205000000
1!
1%
#456210000000
0!
0%
#456215000000
1!
1%
#456220000000
0!
0%
#456225000000
1!
1%
#456230000000
0!
0%
#456235000000
1!
1%
#456240000000
0!
0%
#456245000000
1!
1%
#456250000000
0!
0%
#456255000000
1!
1%
#456260000000
0!
0%
#456265000000
1!
1%
#456270000000
0!
0%
#456275000000
1!
1%
#456280000000
0!
0%
#456285000000
1!
1%
#456290000000
0!
0%
#456295000000
1!
1%
#456300000000
0!
0%
#456305000000
1!
1%
#456310000000
0!
0%
#456315000000
1!
1%
#456320000000
0!
0%
#456325000000
1!
1%
#456330000000
0!
0%
#456335000000
1!
1%
#456340000000
0!
0%
#456345000000
1!
1%
#456350000000
0!
0%
#456355000000
1!
1%
#456360000000
0!
0%
#456365000000
1!
1%
#456370000000
0!
0%
#456375000000
1!
1%
#456380000000
0!
0%
#456385000000
1!
1%
#456390000000
0!
0%
#456395000000
1!
1%
#456400000000
0!
0%
#456405000000
1!
1%
#456410000000
0!
0%
#456415000000
1!
1%
#456420000000
0!
0%
#456425000000
1!
1%
#456430000000
0!
0%
#456435000000
1!
1%
#456440000000
0!
0%
#456445000000
1!
1%
#456450000000
0!
0%
#456455000000
1!
1%
#456460000000
0!
0%
#456465000000
1!
1%
#456470000000
0!
0%
#456475000000
1!
1%
#456480000000
0!
0%
#456485000000
1!
1%
#456490000000
0!
0%
#456495000000
1!
1%
#456500000000
0!
0%
#456505000000
1!
1%
#456510000000
0!
0%
#456515000000
1!
1%
#456520000000
0!
0%
#456525000000
1!
1%
#456530000000
0!
0%
#456535000000
1!
1%
#456540000000
0!
0%
#456545000000
1!
1%
#456550000000
0!
0%
#456555000000
1!
1%
#456560000000
0!
0%
#456565000000
1!
1%
#456570000000
0!
0%
#456575000000
1!
1%
#456580000000
0!
0%
#456585000000
1!
1%
#456590000000
0!
0%
#456595000000
1!
1%
#456600000000
0!
0%
#456605000000
1!
1%
#456610000000
0!
0%
#456615000000
1!
1%
#456620000000
0!
0%
#456625000000
1!
1%
#456630000000
0!
0%
#456635000000
1!
1%
#456640000000
0!
0%
#456645000000
1!
1%
#456650000000
0!
0%
#456655000000
1!
1%
#456660000000
0!
0%
#456665000000
1!
1%
#456670000000
0!
0%
#456675000000
1!
1%
#456680000000
0!
0%
#456685000000
1!
1%
#456690000000
0!
0%
#456695000000
1!
1%
#456700000000
0!
0%
#456705000000
1!
1%
#456710000000
0!
0%
#456715000000
1!
1%
#456720000000
0!
0%
#456725000000
1!
1%
#456730000000
0!
0%
#456735000000
1!
1%
#456740000000
0!
0%
#456745000000
1!
1%
#456750000000
0!
0%
#456755000000
1!
1%
#456760000000
0!
0%
#456765000000
1!
1%
#456770000000
0!
0%
#456775000000
1!
1%
#456780000000
0!
0%
#456785000000
1!
1%
#456790000000
0!
0%
#456795000000
1!
1%
#456800000000
0!
0%
#456805000000
1!
1%
#456810000000
0!
0%
#456815000000
1!
1%
#456820000000
0!
0%
#456825000000
1!
1%
#456830000000
0!
0%
#456835000000
1!
1%
#456840000000
0!
0%
#456845000000
1!
1%
#456850000000
0!
0%
#456855000000
1!
1%
#456860000000
0!
0%
#456865000000
1!
1%
#456870000000
0!
0%
#456875000000
1!
1%
#456880000000
0!
0%
#456885000000
1!
1%
#456890000000
0!
0%
#456895000000
1!
1%
#456900000000
0!
0%
#456905000000
1!
1%
#456910000000
0!
0%
#456915000000
1!
1%
#456920000000
0!
0%
#456925000000
1!
1%
#456930000000
0!
0%
#456935000000
1!
1%
#456940000000
0!
0%
#456945000000
1!
1%
#456950000000
0!
0%
#456955000000
1!
1%
#456960000000
0!
0%
#456965000000
1!
1%
#456970000000
0!
0%
#456975000000
1!
1%
#456980000000
0!
0%
#456985000000
1!
1%
#456990000000
0!
0%
#456995000000
1!
1%
#457000000000
0!
0%
#457005000000
1!
1%
#457010000000
0!
0%
#457015000000
1!
1%
#457020000000
0!
0%
#457025000000
1!
1%
#457030000000
0!
0%
#457035000000
1!
1%
#457040000000
0!
0%
#457045000000
1!
1%
#457050000000
0!
0%
#457055000000
1!
1%
#457060000000
0!
0%
#457065000000
1!
1%
#457070000000
0!
0%
#457075000000
1!
1%
#457080000000
0!
0%
#457085000000
1!
1%
#457090000000
0!
0%
#457095000000
1!
1%
#457100000000
0!
0%
#457105000000
1!
1%
#457110000000
0!
0%
#457115000000
1!
1%
#457120000000
0!
0%
#457125000000
1!
1%
#457130000000
0!
0%
#457135000000
1!
1%
#457140000000
0!
0%
#457145000000
1!
1%
#457150000000
0!
0%
#457155000000
1!
1%
#457160000000
0!
0%
#457165000000
1!
1%
#457170000000
0!
0%
#457175000000
1!
1%
#457180000000
0!
0%
#457185000000
1!
1%
#457190000000
0!
0%
#457195000000
1!
1%
#457200000000
0!
0%
#457205000000
1!
1%
#457210000000
0!
0%
#457215000000
1!
1%
#457220000000
0!
0%
#457225000000
1!
1%
#457230000000
0!
0%
#457235000000
1!
1%
#457240000000
0!
0%
#457245000000
1!
1%
#457250000000
0!
0%
#457255000000
1!
1%
#457260000000
0!
0%
#457265000000
1!
1%
#457270000000
0!
0%
#457275000000
1!
1%
#457280000000
0!
0%
#457285000000
1!
1%
#457290000000
0!
0%
#457295000000
1!
1%
#457300000000
0!
0%
#457305000000
1!
1%
#457310000000
0!
0%
#457315000000
1!
1%
#457320000000
0!
0%
#457325000000
1!
1%
#457330000000
0!
0%
#457335000000
1!
1%
#457340000000
0!
0%
#457345000000
1!
1%
#457350000000
0!
0%
#457355000000
1!
1%
#457360000000
0!
0%
#457365000000
1!
1%
#457370000000
0!
0%
#457375000000
1!
1%
#457380000000
0!
0%
#457385000000
1!
1%
#457390000000
0!
0%
#457395000000
1!
1%
#457400000000
0!
0%
#457405000000
1!
1%
#457410000000
0!
0%
#457415000000
1!
1%
#457420000000
0!
0%
#457425000000
1!
1%
#457430000000
0!
0%
#457435000000
1!
1%
#457440000000
0!
0%
#457445000000
1!
1%
#457450000000
0!
0%
#457455000000
1!
1%
#457460000000
0!
0%
#457465000000
1!
1%
#457470000000
0!
0%
#457475000000
1!
1%
#457480000000
0!
0%
#457485000000
1!
1%
#457490000000
0!
0%
#457495000000
1!
1%
#457500000000
0!
0%
#457505000000
1!
1%
#457510000000
0!
0%
#457515000000
1!
1%
#457520000000
0!
0%
#457525000000
1!
1%
#457530000000
0!
0%
#457535000000
1!
1%
#457540000000
0!
0%
#457545000000
1!
1%
#457550000000
0!
0%
#457555000000
1!
1%
#457560000000
0!
0%
#457565000000
1!
1%
#457570000000
0!
0%
#457575000000
1!
1%
#457580000000
0!
0%
#457585000000
1!
1%
#457590000000
0!
0%
#457595000000
1!
1%
#457600000000
0!
0%
#457605000000
1!
1%
#457610000000
0!
0%
#457615000000
1!
1%
#457620000000
0!
0%
#457625000000
1!
1%
#457630000000
0!
0%
#457635000000
1!
1%
#457640000000
0!
0%
#457645000000
1!
1%
#457650000000
0!
0%
#457655000000
1!
1%
#457660000000
0!
0%
#457665000000
1!
1%
#457670000000
0!
0%
#457675000000
1!
1%
#457680000000
0!
0%
#457685000000
1!
1%
#457690000000
0!
0%
#457695000000
1!
1%
#457700000000
0!
0%
#457705000000
1!
1%
#457710000000
0!
0%
#457715000000
1!
1%
#457720000000
0!
0%
#457725000000
1!
1%
#457730000000
0!
0%
#457735000000
1!
1%
#457740000000
0!
0%
#457745000000
1!
1%
#457750000000
0!
0%
#457755000000
1!
1%
#457760000000
0!
0%
#457765000000
1!
1%
#457770000000
0!
0%
#457775000000
1!
1%
#457780000000
0!
0%
#457785000000
1!
1%
#457790000000
0!
0%
#457795000000
1!
1%
#457800000000
0!
0%
#457805000000
1!
1%
#457810000000
0!
0%
#457815000000
1!
1%
#457820000000
0!
0%
#457825000000
1!
1%
#457830000000
0!
0%
#457835000000
1!
1%
#457840000000
0!
0%
#457845000000
1!
1%
#457850000000
0!
0%
#457855000000
1!
1%
#457860000000
0!
0%
#457865000000
1!
1%
#457870000000
0!
0%
#457875000000
1!
1%
#457880000000
0!
0%
#457885000000
1!
1%
#457890000000
0!
0%
#457895000000
1!
1%
#457900000000
0!
0%
#457905000000
1!
1%
#457910000000
0!
0%
#457915000000
1!
1%
#457920000000
0!
0%
#457925000000
1!
1%
#457930000000
0!
0%
#457935000000
1!
1%
#457940000000
0!
0%
#457945000000
1!
1%
#457950000000
0!
0%
#457955000000
1!
1%
#457960000000
0!
0%
#457965000000
1!
1%
#457970000000
0!
0%
#457975000000
1!
1%
#457980000000
0!
0%
#457985000000
1!
1%
#457990000000
0!
0%
#457995000000
1!
1%
#458000000000
0!
0%
#458005000000
1!
1%
#458010000000
0!
0%
#458015000000
1!
1%
#458020000000
0!
0%
#458025000000
1!
1%
#458030000000
0!
0%
#458035000000
1!
1%
#458040000000
0!
0%
#458045000000
1!
1%
#458050000000
0!
0%
#458055000000
1!
1%
#458060000000
0!
0%
#458065000000
1!
1%
#458070000000
0!
0%
#458075000000
1!
1%
#458080000000
0!
0%
#458085000000
1!
1%
#458090000000
0!
0%
#458095000000
1!
1%
#458100000000
0!
0%
#458105000000
1!
1%
#458110000000
0!
0%
#458115000000
1!
1%
#458120000000
0!
0%
#458125000000
1!
1%
#458130000000
0!
0%
#458135000000
1!
1%
#458140000000
0!
0%
#458145000000
1!
1%
#458150000000
0!
0%
#458155000000
1!
1%
#458160000000
0!
0%
#458165000000
1!
1%
#458170000000
0!
0%
#458175000000
1!
1%
#458180000000
0!
0%
#458185000000
1!
1%
#458190000000
0!
0%
#458195000000
1!
1%
#458200000000
0!
0%
#458205000000
1!
1%
#458210000000
0!
0%
#458215000000
1!
1%
#458220000000
0!
0%
#458225000000
1!
1%
#458230000000
0!
0%
#458235000000
1!
1%
#458240000000
0!
0%
#458245000000
1!
1%
#458250000000
0!
0%
#458255000000
1!
1%
#458260000000
0!
0%
#458265000000
1!
1%
#458270000000
0!
0%
#458275000000
1!
1%
#458280000000
0!
0%
#458285000000
1!
1%
#458290000000
0!
0%
#458295000000
1!
1%
#458300000000
0!
0%
#458305000000
1!
1%
#458310000000
0!
0%
#458315000000
1!
1%
#458320000000
0!
0%
#458325000000
1!
1%
#458330000000
0!
0%
#458335000000
1!
1%
#458340000000
0!
0%
#458345000000
1!
1%
#458350000000
0!
0%
#458355000000
1!
1%
#458360000000
0!
0%
#458365000000
1!
1%
#458370000000
0!
0%
#458375000000
1!
1%
#458380000000
0!
0%
#458385000000
1!
1%
#458390000000
0!
0%
#458395000000
1!
1%
#458400000000
0!
0%
#458405000000
1!
1%
#458410000000
0!
0%
#458415000000
1!
1%
#458420000000
0!
0%
#458425000000
1!
1%
#458430000000
0!
0%
#458435000000
1!
1%
#458440000000
0!
0%
#458445000000
1!
1%
#458450000000
0!
0%
#458455000000
1!
1%
#458460000000
0!
0%
#458465000000
1!
1%
#458470000000
0!
0%
#458475000000
1!
1%
#458480000000
0!
0%
#458485000000
1!
1%
#458490000000
0!
0%
#458495000000
1!
1%
#458500000000
0!
0%
#458505000000
1!
1%
#458510000000
0!
0%
#458515000000
1!
1%
#458520000000
0!
0%
#458525000000
1!
1%
#458530000000
0!
0%
#458535000000
1!
1%
#458540000000
0!
0%
#458545000000
1!
1%
#458550000000
0!
0%
#458555000000
1!
1%
#458560000000
0!
0%
#458565000000
1!
1%
#458570000000
0!
0%
#458575000000
1!
1%
#458580000000
0!
0%
#458585000000
1!
1%
#458590000000
0!
0%
#458595000000
1!
1%
#458600000000
0!
0%
#458605000000
1!
1%
#458610000000
0!
0%
#458615000000
1!
1%
#458620000000
0!
0%
#458625000000
1!
1%
#458630000000
0!
0%
#458635000000
1!
1%
#458640000000
0!
0%
#458645000000
1!
1%
#458650000000
0!
0%
#458655000000
1!
1%
#458660000000
0!
0%
#458665000000
1!
1%
#458670000000
0!
0%
#458675000000
1!
1%
#458680000000
0!
0%
#458685000000
1!
1%
#458690000000
0!
0%
#458695000000
1!
1%
#458700000000
0!
0%
#458705000000
1!
1%
#458710000000
0!
0%
#458715000000
1!
1%
#458720000000
0!
0%
#458725000000
1!
1%
#458730000000
0!
0%
#458735000000
1!
1%
#458740000000
0!
0%
#458745000000
1!
1%
#458750000000
0!
0%
#458755000000
1!
1%
#458760000000
0!
0%
#458765000000
1!
1%
#458770000000
0!
0%
#458775000000
1!
1%
#458780000000
0!
0%
#458785000000
1!
1%
#458790000000
0!
0%
#458795000000
1!
1%
#458800000000
0!
0%
#458805000000
1!
1%
#458810000000
0!
0%
#458815000000
1!
1%
#458820000000
0!
0%
#458825000000
1!
1%
#458830000000
0!
0%
#458835000000
1!
1%
#458840000000
0!
0%
#458845000000
1!
1%
#458850000000
0!
0%
#458855000000
1!
1%
#458860000000
0!
0%
#458865000000
1!
1%
#458870000000
0!
0%
#458875000000
1!
1%
#458880000000
0!
0%
#458885000000
1!
1%
#458890000000
0!
0%
#458895000000
1!
1%
#458900000000
0!
0%
#458905000000
1!
1%
#458910000000
0!
0%
#458915000000
1!
1%
#458920000000
0!
0%
#458925000000
1!
1%
#458930000000
0!
0%
#458935000000
1!
1%
#458940000000
0!
0%
#458945000000
1!
1%
#458950000000
0!
0%
#458955000000
1!
1%
#458960000000
0!
0%
#458965000000
1!
1%
#458970000000
0!
0%
#458975000000
1!
1%
#458980000000
0!
0%
#458985000000
1!
1%
#458990000000
0!
0%
#458995000000
1!
1%
#459000000000
0!
0%
#459005000000
1!
1%
#459010000000
0!
0%
#459015000000
1!
1%
#459020000000
0!
0%
#459025000000
1!
1%
#459030000000
0!
0%
#459035000000
1!
1%
#459040000000
0!
0%
#459045000000
1!
1%
#459050000000
0!
0%
#459055000000
1!
1%
#459060000000
0!
0%
#459065000000
1!
1%
#459070000000
0!
0%
#459075000000
1!
1%
#459080000000
0!
0%
#459085000000
1!
1%
#459090000000
0!
0%
#459095000000
1!
1%
#459100000000
0!
0%
#459105000000
1!
1%
#459110000000
0!
0%
#459115000000
1!
1%
#459120000000
0!
0%
#459125000000
1!
1%
#459130000000
0!
0%
#459135000000
1!
1%
#459140000000
0!
0%
#459145000000
1!
1%
#459150000000
0!
0%
#459155000000
1!
1%
#459160000000
0!
0%
#459165000000
1!
1%
#459170000000
0!
0%
#459175000000
1!
1%
#459180000000
0!
0%
#459185000000
1!
1%
#459190000000
0!
0%
#459195000000
1!
1%
#459200000000
0!
0%
#459205000000
1!
1%
#459210000000
0!
0%
#459215000000
1!
1%
#459220000000
0!
0%
#459225000000
1!
1%
#459230000000
0!
0%
#459235000000
1!
1%
#459240000000
0!
0%
#459245000000
1!
1%
#459250000000
0!
0%
#459255000000
1!
1%
#459260000000
0!
0%
#459265000000
1!
1%
#459270000000
0!
0%
#459275000000
1!
1%
#459280000000
0!
0%
#459285000000
1!
1%
#459290000000
0!
0%
#459295000000
1!
1%
#459300000000
0!
0%
#459305000000
1!
1%
#459310000000
0!
0%
#459315000000
1!
1%
#459320000000
0!
0%
#459325000000
1!
1%
#459330000000
0!
0%
#459335000000
1!
1%
#459340000000
0!
0%
#459345000000
1!
1%
#459350000000
0!
0%
#459355000000
1!
1%
#459360000000
0!
0%
#459365000000
1!
1%
#459370000000
0!
0%
#459375000000
1!
1%
#459380000000
0!
0%
#459385000000
1!
1%
#459390000000
0!
0%
#459395000000
1!
1%
#459400000000
0!
0%
#459405000000
1!
1%
#459410000000
0!
0%
#459415000000
1!
1%
#459420000000
0!
0%
#459425000000
1!
1%
#459430000000
0!
0%
#459435000000
1!
1%
#459440000000
0!
0%
#459445000000
1!
1%
#459450000000
0!
0%
#459455000000
1!
1%
#459460000000
0!
0%
#459465000000
1!
1%
#459470000000
0!
0%
#459475000000
1!
1%
#459480000000
0!
0%
#459485000000
1!
1%
#459490000000
0!
0%
#459495000000
1!
1%
#459500000000
0!
0%
#459505000000
1!
1%
#459510000000
0!
0%
#459515000000
1!
1%
#459520000000
0!
0%
#459525000000
1!
1%
#459530000000
0!
0%
#459535000000
1!
1%
#459540000000
0!
0%
#459545000000
1!
1%
#459550000000
0!
0%
#459555000000
1!
1%
#459560000000
0!
0%
#459565000000
1!
1%
#459570000000
0!
0%
#459575000000
1!
1%
#459580000000
0!
0%
#459585000000
1!
1%
#459590000000
0!
0%
#459595000000
1!
1%
#459600000000
0!
0%
#459605000000
1!
1%
#459610000000
0!
0%
#459615000000
1!
1%
#459620000000
0!
0%
#459625000000
1!
1%
#459630000000
0!
0%
#459635000000
1!
1%
#459640000000
0!
0%
#459645000000
1!
1%
#459650000000
0!
0%
#459655000000
1!
1%
#459660000000
0!
0%
#459665000000
1!
1%
#459670000000
0!
0%
#459675000000
1!
1%
#459680000000
0!
0%
#459685000000
1!
1%
#459690000000
0!
0%
#459695000000
1!
1%
#459700000000
0!
0%
#459705000000
1!
1%
#459710000000
0!
0%
#459715000000
1!
1%
#459720000000
0!
0%
#459725000000
1!
1%
#459730000000
0!
0%
#459735000000
1!
1%
#459740000000
0!
0%
#459745000000
1!
1%
#459750000000
0!
0%
#459755000000
1!
1%
#459760000000
0!
0%
#459765000000
1!
1%
#459770000000
0!
0%
#459775000000
1!
1%
#459780000000
0!
0%
#459785000000
1!
1%
#459790000000
0!
0%
#459795000000
1!
1%
#459800000000
0!
0%
#459805000000
1!
1%
#459810000000
0!
0%
#459815000000
1!
1%
#459820000000
0!
0%
#459825000000
1!
1%
#459830000000
0!
0%
#459835000000
1!
1%
#459840000000
0!
0%
#459845000000
1!
1%
#459850000000
0!
0%
#459855000000
1!
1%
#459860000000
0!
0%
#459865000000
1!
1%
#459870000000
0!
0%
#459875000000
1!
1%
#459880000000
0!
0%
#459885000000
1!
1%
#459890000000
0!
0%
#459895000000
1!
1%
#459900000000
0!
0%
#459905000000
1!
1%
#459910000000
0!
0%
#459915000000
1!
1%
#459920000000
0!
0%
#459925000000
1!
1%
#459930000000
0!
0%
#459935000000
1!
1%
#459940000000
0!
0%
#459945000000
1!
1%
#459950000000
0!
0%
#459955000000
1!
1%
#459960000000
0!
0%
#459965000000
1!
1%
#459970000000
0!
0%
#459975000000
1!
1%
#459980000000
0!
0%
#459985000000
1!
1%
#459990000000
0!
0%
#459995000000
1!
1%
#460000000000
0!
0%
#460005000000
1!
1%
#460010000000
0!
0%
#460015000000
1!
1%
#460020000000
0!
0%
#460025000000
1!
1%
#460030000000
0!
0%
#460035000000
1!
1%
#460040000000
0!
0%
#460045000000
1!
1%
#460050000000
0!
0%
#460055000000
1!
1%
#460060000000
0!
0%
#460065000000
1!
1%
#460070000000
0!
0%
#460075000000
1!
1%
#460080000000
0!
0%
#460085000000
1!
1%
#460090000000
0!
0%
#460095000000
1!
1%
#460100000000
0!
0%
#460105000000
1!
1%
#460110000000
0!
0%
#460115000000
1!
1%
#460120000000
0!
0%
#460125000000
1!
1%
#460130000000
0!
0%
#460135000000
1!
1%
#460140000000
0!
0%
#460145000000
1!
1%
#460150000000
0!
0%
#460155000000
1!
1%
#460160000000
0!
0%
#460165000000
1!
1%
#460170000000
0!
0%
#460175000000
1!
1%
#460180000000
0!
0%
#460185000000
1!
1%
#460190000000
0!
0%
#460195000000
1!
1%
#460200000000
0!
0%
#460205000000
1!
1%
#460210000000
0!
0%
#460215000000
1!
1%
#460220000000
0!
0%
#460225000000
1!
1%
#460230000000
0!
0%
#460235000000
1!
1%
#460240000000
0!
0%
#460245000000
1!
1%
#460250000000
0!
0%
#460255000000
1!
1%
#460260000000
0!
0%
#460265000000
1!
1%
#460270000000
0!
0%
#460275000000
1!
1%
#460280000000
0!
0%
#460285000000
1!
1%
#460290000000
0!
0%
#460295000000
1!
1%
#460300000000
0!
0%
#460305000000
1!
1%
#460310000000
0!
0%
#460315000000
1!
1%
#460320000000
0!
0%
#460325000000
1!
1%
#460330000000
0!
0%
#460335000000
1!
1%
#460340000000
0!
0%
#460345000000
1!
1%
#460350000000
0!
0%
#460355000000
1!
1%
#460360000000
0!
0%
#460365000000
1!
1%
#460370000000
0!
0%
#460375000000
1!
1%
#460380000000
0!
0%
#460385000000
1!
1%
#460390000000
0!
0%
#460395000000
1!
1%
#460400000000
0!
0%
#460405000000
1!
1%
#460410000000
0!
0%
#460415000000
1!
1%
#460420000000
0!
0%
#460425000000
1!
1%
#460430000000
0!
0%
#460435000000
1!
1%
#460440000000
0!
0%
#460445000000
1!
1%
#460450000000
0!
0%
#460455000000
1!
1%
#460460000000
0!
0%
#460465000000
1!
1%
#460470000000
0!
0%
#460475000000
1!
1%
#460480000000
0!
0%
#460485000000
1!
1%
#460490000000
0!
0%
#460495000000
1!
1%
#460500000000
0!
0%
#460505000000
1!
1%
#460510000000
0!
0%
#460515000000
1!
1%
#460520000000
0!
0%
#460525000000
1!
1%
#460530000000
0!
0%
#460535000000
1!
1%
#460540000000
0!
0%
#460545000000
1!
1%
#460550000000
0!
0%
#460555000000
1!
1%
#460560000000
0!
0%
#460565000000
1!
1%
#460570000000
0!
0%
#460575000000
1!
1%
#460580000000
0!
0%
#460585000000
1!
1%
#460590000000
0!
0%
#460595000000
1!
1%
#460600000000
0!
0%
#460605000000
1!
1%
#460610000000
0!
0%
#460615000000
1!
1%
#460620000000
0!
0%
#460625000000
1!
1%
#460630000000
0!
0%
#460635000000
1!
1%
#460640000000
0!
0%
#460645000000
1!
1%
#460650000000
0!
0%
#460655000000
1!
1%
#460660000000
0!
0%
#460665000000
1!
1%
#460670000000
0!
0%
#460675000000
1!
1%
#460680000000
0!
0%
#460685000000
1!
1%
#460690000000
0!
0%
#460695000000
1!
1%
#460700000000
0!
0%
#460705000000
1!
1%
#460710000000
0!
0%
#460715000000
1!
1%
#460720000000
0!
0%
#460725000000
1!
1%
#460730000000
0!
0%
#460735000000
1!
1%
#460740000000
0!
0%
#460745000000
1!
1%
#460750000000
0!
0%
#460755000000
1!
1%
#460760000000
0!
0%
#460765000000
1!
1%
#460770000000
0!
0%
#460775000000
1!
1%
#460780000000
0!
0%
#460785000000
1!
1%
#460790000000
0!
0%
#460795000000
1!
1%
#460800000000
0!
0%
#460805000000
1!
1%
#460810000000
0!
0%
#460815000000
1!
1%
#460820000000
0!
0%
#460825000000
1!
1%
#460830000000
0!
0%
#460835000000
1!
1%
#460840000000
0!
0%
#460845000000
1!
1%
#460850000000
0!
0%
#460855000000
1!
1%
#460860000000
0!
0%
#460865000000
1!
1%
#460870000000
0!
0%
#460875000000
1!
1%
#460880000000
0!
0%
#460885000000
1!
1%
#460890000000
0!
0%
#460895000000
1!
1%
#460900000000
0!
0%
#460905000000
1!
1%
#460910000000
0!
0%
#460915000000
1!
1%
#460920000000
0!
0%
#460925000000
1!
1%
#460930000000
0!
0%
#460935000000
1!
1%
#460940000000
0!
0%
#460945000000
1!
1%
#460950000000
0!
0%
#460955000000
1!
1%
#460960000000
0!
0%
#460965000000
1!
1%
#460970000000
0!
0%
#460975000000
1!
1%
#460980000000
0!
0%
#460985000000
1!
1%
#460990000000
0!
0%
#460995000000
1!
1%
#461000000000
0!
0%
#461005000000
1!
1%
#461010000000
0!
0%
#461015000000
1!
1%
#461020000000
0!
0%
#461025000000
1!
1%
#461030000000
0!
0%
#461035000000
1!
1%
#461040000000
0!
0%
#461045000000
1!
1%
#461050000000
0!
0%
#461055000000
1!
1%
#461060000000
0!
0%
#461065000000
1!
1%
#461070000000
0!
0%
#461075000000
1!
1%
#461080000000
0!
0%
#461085000000
1!
1%
#461090000000
0!
0%
#461095000000
1!
1%
#461100000000
0!
0%
#461105000000
1!
1%
#461110000000
0!
0%
#461115000000
1!
1%
#461120000000
0!
0%
#461125000000
1!
1%
#461130000000
0!
0%
#461135000000
1!
1%
#461140000000
0!
0%
#461145000000
1!
1%
#461150000000
0!
0%
#461155000000
1!
1%
#461160000000
0!
0%
#461165000000
1!
1%
#461170000000
0!
0%
#461175000000
1!
1%
#461180000000
0!
0%
#461185000000
1!
1%
#461190000000
0!
0%
#461195000000
1!
1%
#461200000000
0!
0%
#461205000000
1!
1%
#461210000000
0!
0%
#461215000000
1!
1%
#461220000000
0!
0%
#461225000000
1!
1%
#461230000000
0!
0%
#461235000000
1!
1%
#461240000000
0!
0%
#461245000000
1!
1%
#461250000000
0!
0%
#461255000000
1!
1%
#461260000000
0!
0%
#461265000000
1!
1%
#461270000000
0!
0%
#461275000000
1!
1%
#461280000000
0!
0%
#461285000000
1!
1%
#461290000000
0!
0%
#461295000000
1!
1%
#461300000000
0!
0%
#461305000000
1!
1%
#461310000000
0!
0%
#461315000000
1!
1%
#461320000000
0!
0%
#461325000000
1!
1%
#461330000000
0!
0%
#461335000000
1!
1%
#461340000000
0!
0%
#461345000000
1!
1%
#461350000000
0!
0%
#461355000000
1!
1%
#461360000000
0!
0%
#461365000000
1!
1%
#461370000000
0!
0%
#461375000000
1!
1%
#461380000000
0!
0%
#461385000000
1!
1%
#461390000000
0!
0%
#461395000000
1!
1%
#461400000000
0!
0%
#461405000000
1!
1%
#461410000000
0!
0%
#461415000000
1!
1%
#461420000000
0!
0%
#461425000000
1!
1%
#461430000000
0!
0%
#461435000000
1!
1%
#461440000000
0!
0%
#461445000000
1!
1%
#461450000000
0!
0%
#461455000000
1!
1%
#461460000000
0!
0%
#461465000000
1!
1%
#461470000000
0!
0%
#461475000000
1!
1%
#461480000000
0!
0%
#461485000000
1!
1%
#461490000000
0!
0%
#461495000000
1!
1%
#461500000000
0!
0%
#461505000000
1!
1%
#461510000000
0!
0%
#461515000000
1!
1%
#461520000000
0!
0%
#461525000000
1!
1%
#461530000000
0!
0%
#461535000000
1!
1%
#461540000000
0!
0%
#461545000000
1!
1%
#461550000000
0!
0%
#461555000000
1!
1%
#461560000000
0!
0%
#461565000000
1!
1%
#461570000000
0!
0%
#461575000000
1!
1%
#461580000000
0!
0%
#461585000000
1!
1%
#461590000000
0!
0%
#461595000000
1!
1%
#461600000000
0!
0%
#461605000000
1!
1%
#461610000000
0!
0%
#461615000000
1!
1%
#461620000000
0!
0%
#461625000000
1!
1%
#461630000000
0!
0%
#461635000000
1!
1%
#461640000000
0!
0%
#461645000000
1!
1%
#461650000000
0!
0%
#461655000000
1!
1%
#461660000000
0!
0%
#461665000000
1!
1%
#461670000000
0!
0%
#461675000000
1!
1%
#461680000000
0!
0%
#461685000000
1!
1%
#461690000000
0!
0%
#461695000000
1!
1%
#461700000000
0!
0%
#461705000000
1!
1%
#461710000000
0!
0%
#461715000000
1!
1%
#461720000000
0!
0%
#461725000000
1!
1%
#461730000000
0!
0%
#461735000000
1!
1%
#461740000000
0!
0%
#461745000000
1!
1%
#461750000000
0!
0%
#461755000000
1!
1%
#461760000000
0!
0%
#461765000000
1!
1%
#461770000000
0!
0%
#461775000000
1!
1%
#461780000000
0!
0%
#461785000000
1!
1%
#461790000000
0!
0%
#461795000000
1!
1%
#461800000000
0!
0%
#461805000000
1!
1%
#461810000000
0!
0%
#461815000000
1!
1%
#461820000000
0!
0%
#461825000000
1!
1%
#461830000000
0!
0%
#461835000000
1!
1%
#461840000000
0!
0%
#461845000000
1!
1%
#461850000000
0!
0%
#461855000000
1!
1%
#461860000000
0!
0%
#461865000000
1!
1%
#461870000000
0!
0%
#461875000000
1!
1%
#461880000000
0!
0%
#461885000000
1!
1%
#461890000000
0!
0%
#461895000000
1!
1%
#461900000000
0!
0%
#461905000000
1!
1%
#461910000000
0!
0%
#461915000000
1!
1%
#461920000000
0!
0%
#461925000000
1!
1%
#461930000000
0!
0%
#461935000000
1!
1%
#461940000000
0!
0%
#461945000000
1!
1%
#461950000000
0!
0%
#461955000000
1!
1%
#461960000000
0!
0%
#461965000000
1!
1%
#461970000000
0!
0%
#461975000000
1!
1%
#461980000000
0!
0%
#461985000000
1!
1%
#461990000000
0!
0%
#461995000000
1!
1%
#462000000000
0!
0%
#462005000000
1!
1%
#462010000000
0!
0%
#462015000000
1!
1%
#462020000000
0!
0%
#462025000000
1!
1%
#462030000000
0!
0%
#462035000000
1!
1%
#462040000000
0!
0%
#462045000000
1!
1%
#462050000000
0!
0%
#462055000000
1!
1%
#462060000000
0!
0%
#462065000000
1!
1%
#462070000000
0!
0%
#462075000000
1!
1%
#462080000000
0!
0%
#462085000000
1!
1%
#462090000000
0!
0%
#462095000000
1!
1%
#462100000000
0!
0%
#462105000000
1!
1%
#462110000000
0!
0%
#462115000000
1!
1%
#462120000000
0!
0%
#462125000000
1!
1%
#462130000000
0!
0%
#462135000000
1!
1%
#462140000000
0!
0%
#462145000000
1!
1%
#462150000000
0!
0%
#462155000000
1!
1%
#462160000000
0!
0%
#462165000000
1!
1%
#462170000000
0!
0%
#462175000000
1!
1%
#462180000000
0!
0%
#462185000000
1!
1%
#462190000000
0!
0%
#462195000000
1!
1%
#462200000000
0!
0%
#462205000000
1!
1%
#462210000000
0!
0%
#462215000000
1!
1%
#462220000000
0!
0%
#462225000000
1!
1%
#462230000000
0!
0%
#462235000000
1!
1%
#462240000000
0!
0%
#462245000000
1!
1%
#462250000000
0!
0%
#462255000000
1!
1%
#462260000000
0!
0%
#462265000000
1!
1%
#462270000000
0!
0%
#462275000000
1!
1%
#462280000000
0!
0%
#462285000000
1!
1%
#462290000000
0!
0%
#462295000000
1!
1%
#462300000000
0!
0%
#462305000000
1!
1%
#462310000000
0!
0%
#462315000000
1!
1%
#462320000000
0!
0%
#462325000000
1!
1%
#462330000000
0!
0%
#462335000000
1!
1%
#462340000000
0!
0%
#462345000000
1!
1%
#462350000000
0!
0%
#462355000000
1!
1%
#462360000000
0!
0%
#462365000000
1!
1%
#462370000000
0!
0%
#462375000000
1!
1%
#462380000000
0!
0%
#462385000000
1!
1%
#462390000000
0!
0%
#462395000000
1!
1%
#462400000000
0!
0%
#462405000000
1!
1%
#462410000000
0!
0%
#462415000000
1!
1%
#462420000000
0!
0%
#462425000000
1!
1%
#462430000000
0!
0%
#462435000000
1!
1%
#462440000000
0!
0%
#462445000000
1!
1%
#462450000000
0!
0%
#462455000000
1!
1%
#462460000000
0!
0%
#462465000000
1!
1%
#462470000000
0!
0%
#462475000000
1!
1%
#462480000000
0!
0%
#462485000000
1!
1%
#462490000000
0!
0%
#462495000000
1!
1%
#462500000000
0!
0%
#462505000000
1!
1%
#462510000000
0!
0%
#462515000000
1!
1%
#462520000000
0!
0%
#462525000000
1!
1%
#462530000000
0!
0%
#462535000000
1!
1%
#462540000000
0!
0%
#462545000000
1!
1%
#462550000000
0!
0%
#462555000000
1!
1%
#462560000000
0!
0%
#462565000000
1!
1%
#462570000000
0!
0%
#462575000000
1!
1%
#462580000000
0!
0%
#462585000000
1!
1%
#462590000000
0!
0%
#462595000000
1!
1%
#462600000000
0!
0%
#462605000000
1!
1%
#462610000000
0!
0%
#462615000000
1!
1%
#462620000000
0!
0%
#462625000000
1!
1%
#462630000000
0!
0%
#462635000000
1!
1%
#462640000000
0!
0%
#462645000000
1!
1%
#462650000000
0!
0%
#462655000000
1!
1%
#462660000000
0!
0%
#462665000000
1!
1%
#462670000000
0!
0%
#462675000000
1!
1%
#462680000000
0!
0%
#462685000000
1!
1%
#462690000000
0!
0%
#462695000000
1!
1%
#462700000000
0!
0%
#462705000000
1!
1%
#462710000000
0!
0%
#462715000000
1!
1%
#462720000000
0!
0%
#462725000000
1!
1%
#462730000000
0!
0%
#462735000000
1!
1%
#462740000000
0!
0%
#462745000000
1!
1%
#462750000000
0!
0%
#462755000000
1!
1%
#462760000000
0!
0%
#462765000000
1!
1%
#462770000000
0!
0%
#462775000000
1!
1%
#462780000000
0!
0%
#462785000000
1!
1%
#462790000000
0!
0%
#462795000000
1!
1%
#462800000000
0!
0%
#462805000000
1!
1%
#462810000000
0!
0%
#462815000000
1!
1%
#462820000000
0!
0%
#462825000000
1!
1%
#462830000000
0!
0%
#462835000000
1!
1%
#462840000000
0!
0%
#462845000000
1!
1%
#462850000000
0!
0%
#462855000000
1!
1%
#462860000000
0!
0%
#462865000000
1!
1%
#462870000000
0!
0%
#462875000000
1!
1%
#462880000000
0!
0%
#462885000000
1!
1%
#462890000000
0!
0%
#462895000000
1!
1%
#462900000000
0!
0%
#462905000000
1!
1%
#462910000000
0!
0%
#462915000000
1!
1%
#462920000000
0!
0%
#462925000000
1!
1%
#462930000000
0!
0%
#462935000000
1!
1%
#462940000000
0!
0%
#462945000000
1!
1%
#462950000000
0!
0%
#462955000000
1!
1%
#462960000000
0!
0%
#462965000000
1!
1%
#462970000000
0!
0%
#462975000000
1!
1%
#462980000000
0!
0%
#462985000000
1!
1%
#462990000000
0!
0%
#462995000000
1!
1%
#463000000000
0!
0%
#463005000000
1!
1%
#463010000000
0!
0%
#463015000000
1!
1%
#463020000000
0!
0%
#463025000000
1!
1%
#463030000000
0!
0%
#463035000000
1!
1%
#463040000000
0!
0%
#463045000000
1!
1%
#463050000000
0!
0%
#463055000000
1!
1%
#463060000000
0!
0%
#463065000000
1!
1%
#463070000000
0!
0%
#463075000000
1!
1%
#463080000000
0!
0%
#463085000000
1!
1%
#463090000000
0!
0%
#463095000000
1!
1%
#463100000000
0!
0%
#463105000000
1!
1%
#463110000000
0!
0%
#463115000000
1!
1%
#463120000000
0!
0%
#463125000000
1!
1%
#463130000000
0!
0%
#463135000000
1!
1%
#463140000000
0!
0%
#463145000000
1!
1%
#463150000000
0!
0%
#463155000000
1!
1%
#463160000000
0!
0%
#463165000000
1!
1%
#463170000000
0!
0%
#463175000000
1!
1%
#463180000000
0!
0%
#463185000000
1!
1%
#463190000000
0!
0%
#463195000000
1!
1%
#463200000000
0!
0%
#463205000000
1!
1%
#463210000000
0!
0%
#463215000000
1!
1%
#463220000000
0!
0%
#463225000000
1!
1%
#463230000000
0!
0%
#463235000000
1!
1%
#463240000000
0!
0%
#463245000000
1!
1%
#463250000000
0!
0%
#463255000000
1!
1%
#463260000000
0!
0%
#463265000000
1!
1%
#463270000000
0!
0%
#463275000000
1!
1%
#463280000000
0!
0%
#463285000000
1!
1%
#463290000000
0!
0%
#463295000000
1!
1%
#463300000000
0!
0%
#463305000000
1!
1%
#463310000000
0!
0%
#463315000000
1!
1%
#463320000000
0!
0%
#463325000000
1!
1%
#463330000000
0!
0%
#463335000000
1!
1%
#463340000000
0!
0%
#463345000000
1!
1%
#463350000000
0!
0%
#463355000000
1!
1%
#463360000000
0!
0%
#463365000000
1!
1%
#463370000000
0!
0%
#463375000000
1!
1%
#463380000000
0!
0%
#463385000000
1!
1%
#463390000000
0!
0%
#463395000000
1!
1%
#463400000000
0!
0%
#463405000000
1!
1%
#463410000000
0!
0%
#463415000000
1!
1%
#463420000000
0!
0%
#463425000000
1!
1%
#463430000000
0!
0%
#463435000000
1!
1%
#463440000000
0!
0%
#463445000000
1!
1%
#463450000000
0!
0%
#463455000000
1!
1%
#463460000000
0!
0%
#463465000000
1!
1%
#463470000000
0!
0%
#463475000000
1!
1%
#463480000000
0!
0%
#463485000000
1!
1%
#463490000000
0!
0%
#463495000000
1!
1%
#463500000000
0!
0%
#463505000000
1!
1%
#463510000000
0!
0%
#463515000000
1!
1%
#463520000000
0!
0%
#463525000000
1!
1%
#463530000000
0!
0%
#463535000000
1!
1%
#463540000000
0!
0%
#463545000000
1!
1%
#463550000000
0!
0%
#463555000000
1!
1%
#463560000000
0!
0%
#463565000000
1!
1%
#463570000000
0!
0%
#463575000000
1!
1%
#463580000000
0!
0%
#463585000000
1!
1%
#463590000000
0!
0%
#463595000000
1!
1%
#463600000000
0!
0%
#463605000000
1!
1%
#463610000000
0!
0%
#463615000000
1!
1%
#463620000000
0!
0%
#463625000000
1!
1%
#463630000000
0!
0%
#463635000000
1!
1%
#463640000000
0!
0%
#463645000000
1!
1%
#463650000000
0!
0%
#463655000000
1!
1%
#463660000000
0!
0%
#463665000000
1!
1%
#463670000000
0!
0%
#463675000000
1!
1%
#463680000000
0!
0%
#463685000000
1!
1%
#463690000000
0!
0%
#463695000000
1!
1%
#463700000000
0!
0%
#463705000000
1!
1%
#463710000000
0!
0%
#463715000000
1!
1%
#463720000000
0!
0%
#463725000000
1!
1%
#463730000000
0!
0%
#463735000000
1!
1%
#463740000000
0!
0%
#463745000000
1!
1%
#463750000000
0!
0%
#463755000000
1!
1%
#463760000000
0!
0%
#463765000000
1!
1%
#463770000000
0!
0%
#463775000000
1!
1%
#463780000000
0!
0%
#463785000000
1!
1%
#463790000000
0!
0%
#463795000000
1!
1%
#463800000000
0!
0%
#463805000000
1!
1%
#463810000000
0!
0%
#463815000000
1!
1%
#463820000000
0!
0%
#463825000000
1!
1%
#463830000000
0!
0%
#463835000000
1!
1%
#463840000000
0!
0%
#463845000000
1!
1%
#463850000000
0!
0%
#463855000000
1!
1%
#463860000000
0!
0%
#463865000000
1!
1%
#463870000000
0!
0%
#463875000000
1!
1%
#463880000000
0!
0%
#463885000000
1!
1%
#463890000000
0!
0%
#463895000000
1!
1%
#463900000000
0!
0%
#463905000000
1!
1%
#463910000000
0!
0%
#463915000000
1!
1%
#463920000000
0!
0%
#463925000000
1!
1%
#463930000000
0!
0%
#463935000000
1!
1%
#463940000000
0!
0%
#463945000000
1!
1%
#463950000000
0!
0%
#463955000000
1!
1%
#463960000000
0!
0%
#463965000000
1!
1%
#463970000000
0!
0%
#463975000000
1!
1%
#463980000000
0!
0%
#463985000000
1!
1%
#463990000000
0!
0%
#463995000000
1!
1%
#464000000000
0!
0%
#464005000000
1!
1%
#464010000000
0!
0%
#464015000000
1!
1%
#464020000000
0!
0%
#464025000000
1!
1%
#464030000000
0!
0%
#464035000000
1!
1%
#464040000000
0!
0%
#464045000000
1!
1%
#464050000000
0!
0%
#464055000000
1!
1%
#464060000000
0!
0%
#464065000000
1!
1%
#464070000000
0!
0%
#464075000000
1!
1%
#464080000000
0!
0%
#464085000000
1!
1%
#464090000000
0!
0%
#464095000000
1!
1%
#464100000000
0!
0%
#464105000000
1!
1%
#464110000000
0!
0%
#464115000000
1!
1%
#464120000000
0!
0%
#464125000000
1!
1%
#464130000000
0!
0%
#464135000000
1!
1%
#464140000000
0!
0%
#464145000000
1!
1%
#464150000000
0!
0%
#464155000000
1!
1%
#464160000000
0!
0%
#464165000000
1!
1%
#464170000000
0!
0%
#464175000000
1!
1%
#464180000000
0!
0%
#464185000000
1!
1%
#464190000000
0!
0%
#464195000000
1!
1%
#464200000000
0!
0%
#464205000000
1!
1%
#464210000000
0!
0%
#464215000000
1!
1%
#464220000000
0!
0%
#464225000000
1!
1%
#464230000000
0!
0%
#464235000000
1!
1%
#464240000000
0!
0%
#464245000000
1!
1%
#464250000000
0!
0%
#464255000000
1!
1%
#464260000000
0!
0%
#464265000000
1!
1%
#464270000000
0!
0%
#464275000000
1!
1%
#464280000000
0!
0%
#464285000000
1!
1%
#464290000000
0!
0%
#464295000000
1!
1%
#464300000000
0!
0%
#464305000000
1!
1%
#464310000000
0!
0%
#464315000000
1!
1%
#464320000000
0!
0%
#464325000000
1!
1%
#464330000000
0!
0%
#464335000000
1!
1%
#464340000000
0!
0%
#464345000000
1!
1%
#464350000000
0!
0%
#464355000000
1!
1%
#464360000000
0!
0%
#464365000000
1!
1%
#464370000000
0!
0%
#464375000000
1!
1%
#464380000000
0!
0%
#464385000000
1!
1%
#464390000000
0!
0%
#464395000000
1!
1%
#464400000000
0!
0%
#464405000000
1!
1%
#464410000000
0!
0%
#464415000000
1!
1%
#464420000000
0!
0%
#464425000000
1!
1%
#464430000000
0!
0%
#464435000000
1!
1%
#464440000000
0!
0%
#464445000000
1!
1%
#464450000000
0!
0%
#464455000000
1!
1%
#464460000000
0!
0%
#464465000000
1!
1%
#464470000000
0!
0%
#464475000000
1!
1%
#464480000000
0!
0%
#464485000000
1!
1%
#464490000000
0!
0%
#464495000000
1!
1%
#464500000000
0!
0%
#464505000000
1!
1%
#464510000000
0!
0%
#464515000000
1!
1%
#464520000000
0!
0%
#464525000000
1!
1%
#464530000000
0!
0%
#464535000000
1!
1%
#464540000000
0!
0%
#464545000000
1!
1%
#464550000000
0!
0%
#464555000000
1!
1%
#464560000000
0!
0%
#464565000000
1!
1%
#464570000000
0!
0%
#464575000000
1!
1%
#464580000000
0!
0%
#464585000000
1!
1%
#464590000000
0!
0%
#464595000000
1!
1%
#464600000000
0!
0%
#464605000000
1!
1%
#464610000000
0!
0%
#464615000000
1!
1%
#464620000000
0!
0%
#464625000000
1!
1%
#464630000000
0!
0%
#464635000000
1!
1%
#464640000000
0!
0%
#464645000000
1!
1%
#464650000000
0!
0%
#464655000000
1!
1%
#464660000000
0!
0%
#464665000000
1!
1%
#464670000000
0!
0%
#464675000000
1!
1%
#464680000000
0!
0%
#464685000000
1!
1%
#464690000000
0!
0%
#464695000000
1!
1%
#464700000000
0!
0%
#464705000000
1!
1%
#464710000000
0!
0%
#464715000000
1!
1%
#464720000000
0!
0%
#464725000000
1!
1%
#464730000000
0!
0%
#464735000000
1!
1%
#464740000000
0!
0%
#464745000000
1!
1%
#464750000000
0!
0%
#464755000000
1!
1%
#464760000000
0!
0%
#464765000000
1!
1%
#464770000000
0!
0%
#464775000000
1!
1%
#464780000000
0!
0%
#464785000000
1!
1%
#464790000000
0!
0%
#464795000000
1!
1%
#464800000000
0!
0%
#464805000000
1!
1%
#464810000000
0!
0%
#464815000000
1!
1%
#464820000000
0!
0%
#464825000000
1!
1%
#464830000000
0!
0%
#464835000000
1!
1%
#464840000000
0!
0%
#464845000000
1!
1%
#464850000000
0!
0%
#464855000000
1!
1%
#464860000000
0!
0%
#464865000000
1!
1%
#464870000000
0!
0%
#464875000000
1!
1%
#464880000000
0!
0%
#464885000000
1!
1%
#464890000000
0!
0%
#464895000000
1!
1%
#464900000000
0!
0%
#464905000000
1!
1%
#464910000000
0!
0%
#464915000000
1!
1%
#464920000000
0!
0%
#464925000000
1!
1%
#464930000000
0!
0%
#464935000000
1!
1%
#464940000000
0!
0%
#464945000000
1!
1%
#464950000000
0!
0%
#464955000000
1!
1%
#464960000000
0!
0%
#464965000000
1!
1%
#464970000000
0!
0%
#464975000000
1!
1%
#464980000000
0!
0%
#464985000000
1!
1%
#464990000000
0!
0%
#464995000000
1!
1%
#465000000000
0!
0%
#465005000000
1!
1%
#465010000000
0!
0%
#465015000000
1!
1%
#465020000000
0!
0%
#465025000000
1!
1%
#465030000000
0!
0%
#465035000000
1!
1%
#465040000000
0!
0%
#465045000000
1!
1%
#465050000000
0!
0%
#465055000000
1!
1%
#465060000000
0!
0%
#465065000000
1!
1%
#465070000000
0!
0%
#465075000000
1!
1%
#465080000000
0!
0%
#465085000000
1!
1%
#465090000000
0!
0%
#465095000000
1!
1%
#465100000000
0!
0%
#465105000000
1!
1%
#465110000000
0!
0%
#465115000000
1!
1%
#465120000000
0!
0%
#465125000000
1!
1%
#465130000000
0!
0%
#465135000000
1!
1%
#465140000000
0!
0%
#465145000000
1!
1%
#465150000000
0!
0%
#465155000000
1!
1%
#465160000000
0!
0%
#465165000000
1!
1%
#465170000000
0!
0%
#465175000000
1!
1%
#465180000000
0!
0%
#465185000000
1!
1%
#465190000000
0!
0%
#465195000000
1!
1%
#465200000000
0!
0%
#465205000000
1!
1%
#465210000000
0!
0%
#465215000000
1!
1%
#465220000000
0!
0%
#465225000000
1!
1%
#465230000000
0!
0%
#465235000000
1!
1%
#465240000000
0!
0%
#465245000000
1!
1%
#465250000000
0!
0%
#465255000000
1!
1%
#465260000000
0!
0%
#465265000000
1!
1%
#465270000000
0!
0%
#465275000000
1!
1%
#465280000000
0!
0%
#465285000000
1!
1%
#465290000000
0!
0%
#465295000000
1!
1%
#465300000000
0!
0%
#465305000000
1!
1%
#465310000000
0!
0%
#465315000000
1!
1%
#465320000000
0!
0%
#465325000000
1!
1%
#465330000000
0!
0%
#465335000000
1!
1%
#465340000000
0!
0%
#465345000000
1!
1%
#465350000000
0!
0%
#465355000000
1!
1%
#465360000000
0!
0%
#465365000000
1!
1%
#465370000000
0!
0%
#465375000000
1!
1%
#465380000000
0!
0%
#465385000000
1!
1%
#465390000000
0!
0%
#465395000000
1!
1%
#465400000000
0!
0%
#465405000000
1!
1%
#465410000000
0!
0%
#465415000000
1!
1%
#465420000000
0!
0%
#465425000000
1!
1%
#465430000000
0!
0%
#465435000000
1!
1%
#465440000000
0!
0%
#465445000000
1!
1%
#465450000000
0!
0%
#465455000000
1!
1%
#465460000000
0!
0%
#465465000000
1!
1%
#465470000000
0!
0%
#465475000000
1!
1%
#465480000000
0!
0%
#465485000000
1!
1%
#465490000000
0!
0%
#465495000000
1!
1%
#465500000000
0!
0%
#465505000000
1!
1%
#465510000000
0!
0%
#465515000000
1!
1%
#465520000000
0!
0%
#465525000000
1!
1%
#465530000000
0!
0%
#465535000000
1!
1%
#465540000000
0!
0%
#465545000000
1!
1%
#465550000000
0!
0%
#465555000000
1!
1%
#465560000000
0!
0%
#465565000000
1!
1%
#465570000000
0!
0%
#465575000000
1!
1%
#465580000000
0!
0%
#465585000000
1!
1%
#465590000000
0!
0%
#465595000000
1!
1%
#465600000000
0!
0%
#465605000000
1!
1%
#465610000000
0!
0%
#465615000000
1!
1%
#465620000000
0!
0%
#465625000000
1!
1%
#465630000000
0!
0%
#465635000000
1!
1%
#465640000000
0!
0%
#465645000000
1!
1%
#465650000000
0!
0%
#465655000000
1!
1%
#465660000000
0!
0%
#465665000000
1!
1%
#465670000000
0!
0%
#465675000000
1!
1%
#465680000000
0!
0%
#465685000000
1!
1%
#465690000000
0!
0%
#465695000000
1!
1%
#465700000000
0!
0%
#465705000000
1!
1%
#465710000000
0!
0%
#465715000000
1!
1%
#465720000000
0!
0%
#465725000000
1!
1%
#465730000000
0!
0%
#465735000000
1!
1%
#465740000000
0!
0%
#465745000000
1!
1%
#465750000000
0!
0%
#465755000000
1!
1%
#465760000000
0!
0%
#465765000000
1!
1%
#465770000000
0!
0%
#465775000000
1!
1%
#465780000000
0!
0%
#465785000000
1!
1%
#465790000000
0!
0%
#465795000000
1!
1%
#465800000000
0!
0%
#465805000000
1!
1%
#465810000000
0!
0%
#465815000000
1!
1%
#465820000000
0!
0%
#465825000000
1!
1%
#465830000000
0!
0%
#465835000000
1!
1%
#465840000000
0!
0%
#465845000000
1!
1%
#465850000000
0!
0%
#465855000000
1!
1%
#465860000000
0!
0%
#465865000000
1!
1%
#465870000000
0!
0%
#465875000000
1!
1%
#465880000000
0!
0%
#465885000000
1!
1%
#465890000000
0!
0%
#465895000000
1!
1%
#465900000000
0!
0%
#465905000000
1!
1%
#465910000000
0!
0%
#465915000000
1!
1%
#465920000000
0!
0%
#465925000000
1!
1%
#465930000000
0!
0%
#465935000000
1!
1%
#465940000000
0!
0%
#465945000000
1!
1%
#465950000000
0!
0%
#465955000000
1!
1%
#465960000000
0!
0%
#465965000000
1!
1%
#465970000000
0!
0%
#465975000000
1!
1%
#465980000000
0!
0%
#465985000000
1!
1%
#465990000000
0!
0%
#465995000000
1!
1%
#466000000000
0!
0%
#466005000000
1!
1%
#466010000000
0!
0%
#466015000000
1!
1%
#466020000000
0!
0%
#466025000000
1!
1%
#466030000000
0!
0%
#466035000000
1!
1%
#466040000000
0!
0%
#466045000000
1!
1%
#466050000000
0!
0%
#466055000000
1!
1%
#466060000000
0!
0%
#466065000000
1!
1%
#466070000000
0!
0%
#466075000000
1!
1%
#466080000000
0!
0%
#466085000000
1!
1%
#466090000000
0!
0%
#466095000000
1!
1%
#466100000000
0!
0%
#466105000000
1!
1%
#466110000000
0!
0%
#466115000000
1!
1%
#466120000000
0!
0%
#466125000000
1!
1%
#466130000000
0!
0%
#466135000000
1!
1%
#466140000000
0!
0%
#466145000000
1!
1%
#466150000000
0!
0%
#466155000000
1!
1%
#466160000000
0!
0%
#466165000000
1!
1%
#466170000000
0!
0%
#466175000000
1!
1%
#466180000000
0!
0%
#466185000000
1!
1%
#466190000000
0!
0%
#466195000000
1!
1%
#466200000000
0!
0%
#466205000000
1!
1%
#466210000000
0!
0%
#466215000000
1!
1%
#466220000000
0!
0%
#466225000000
1!
1%
#466230000000
0!
0%
#466235000000
1!
1%
#466240000000
0!
0%
#466245000000
1!
1%
#466250000000
0!
0%
#466255000000
1!
1%
#466260000000
0!
0%
#466265000000
1!
1%
#466270000000
0!
0%
#466275000000
1!
1%
#466280000000
0!
0%
#466285000000
1!
1%
#466290000000
0!
0%
#466295000000
1!
1%
#466300000000
0!
0%
#466305000000
1!
1%
#466310000000
0!
0%
#466315000000
1!
1%
#466320000000
0!
0%
#466325000000
1!
1%
#466330000000
0!
0%
#466335000000
1!
1%
#466340000000
0!
0%
#466345000000
1!
1%
#466350000000
0!
0%
#466355000000
1!
1%
#466360000000
0!
0%
#466365000000
1!
1%
#466370000000
0!
0%
#466375000000
1!
1%
#466380000000
0!
0%
#466385000000
1!
1%
#466390000000
0!
0%
#466395000000
1!
1%
#466400000000
0!
0%
#466405000000
1!
1%
#466410000000
0!
0%
#466415000000
1!
1%
#466420000000
0!
0%
#466425000000
1!
1%
#466430000000
0!
0%
#466435000000
1!
1%
#466440000000
0!
0%
#466445000000
1!
1%
#466450000000
0!
0%
#466455000000
1!
1%
#466460000000
0!
0%
#466465000000
1!
1%
#466470000000
0!
0%
#466475000000
1!
1%
#466480000000
0!
0%
#466485000000
1!
1%
#466490000000
0!
0%
#466495000000
1!
1%
#466500000000
0!
0%
#466505000000
1!
1%
#466510000000
0!
0%
#466515000000
1!
1%
#466520000000
0!
0%
#466525000000
1!
1%
#466530000000
0!
0%
#466535000000
1!
1%
#466540000000
0!
0%
#466545000000
1!
1%
#466550000000
0!
0%
#466555000000
1!
1%
#466560000000
0!
0%
#466565000000
1!
1%
#466570000000
0!
0%
#466575000000
1!
1%
#466580000000
0!
0%
#466585000000
1!
1%
#466590000000
0!
0%
#466595000000
1!
1%
#466600000000
0!
0%
#466605000000
1!
1%
#466610000000
0!
0%
#466615000000
1!
1%
#466620000000
0!
0%
#466625000000
1!
1%
#466630000000
0!
0%
#466635000000
1!
1%
#466640000000
0!
0%
#466645000000
1!
1%
#466650000000
0!
0%
#466655000000
1!
1%
#466660000000
0!
0%
#466665000000
1!
1%
#466670000000
0!
0%
#466675000000
1!
1%
#466680000000
0!
0%
#466685000000
1!
1%
#466690000000
0!
0%
#466695000000
1!
1%
#466700000000
0!
0%
#466705000000
1!
1%
#466710000000
0!
0%
#466715000000
1!
1%
#466720000000
0!
0%
#466725000000
1!
1%
#466730000000
0!
0%
#466735000000
1!
1%
#466740000000
0!
0%
#466745000000
1!
1%
#466750000000
0!
0%
#466755000000
1!
1%
#466760000000
0!
0%
#466765000000
1!
1%
#466770000000
0!
0%
#466775000000
1!
1%
#466780000000
0!
0%
#466785000000
1!
1%
#466790000000
0!
0%
#466795000000
1!
1%
#466800000000
0!
0%
#466805000000
1!
1%
#466810000000
0!
0%
#466815000000
1!
1%
#466820000000
0!
0%
#466825000000
1!
1%
#466830000000
0!
0%
#466835000000
1!
1%
#466840000000
0!
0%
#466845000000
1!
1%
#466850000000
0!
0%
#466855000000
1!
1%
#466860000000
0!
0%
#466865000000
1!
1%
#466870000000
0!
0%
#466875000000
1!
1%
#466880000000
0!
0%
#466885000000
1!
1%
#466890000000
0!
0%
#466895000000
1!
1%
#466900000000
0!
0%
#466905000000
1!
1%
#466910000000
0!
0%
#466915000000
1!
1%
#466920000000
0!
0%
#466925000000
1!
1%
#466930000000
0!
0%
#466935000000
1!
1%
#466940000000
0!
0%
#466945000000
1!
1%
#466950000000
0!
0%
#466955000000
1!
1%
#466960000000
0!
0%
#466965000000
1!
1%
#466970000000
0!
0%
#466975000000
1!
1%
#466980000000
0!
0%
#466985000000
1!
1%
#466990000000
0!
0%
#466995000000
1!
1%
#467000000000
0!
0%
#467005000000
1!
1%
#467010000000
0!
0%
#467015000000
1!
1%
#467020000000
0!
0%
#467025000000
1!
1%
#467030000000
0!
0%
#467035000000
1!
1%
#467040000000
0!
0%
#467045000000
1!
1%
#467050000000
0!
0%
#467055000000
1!
1%
#467060000000
0!
0%
#467065000000
1!
1%
#467070000000
0!
0%
#467075000000
1!
1%
#467080000000
0!
0%
#467085000000
1!
1%
#467090000000
0!
0%
#467095000000
1!
1%
#467100000000
0!
0%
#467105000000
1!
1%
#467110000000
0!
0%
#467115000000
1!
1%
#467120000000
0!
0%
#467125000000
1!
1%
#467130000000
0!
0%
#467135000000
1!
1%
#467140000000
0!
0%
#467145000000
1!
1%
#467150000000
0!
0%
#467155000000
1!
1%
#467160000000
0!
0%
#467165000000
1!
1%
#467170000000
0!
0%
#467175000000
1!
1%
#467180000000
0!
0%
#467185000000
1!
1%
#467190000000
0!
0%
#467195000000
1!
1%
#467200000000
0!
0%
#467205000000
1!
1%
#467210000000
0!
0%
#467215000000
1!
1%
#467220000000
0!
0%
#467225000000
1!
1%
#467230000000
0!
0%
#467235000000
1!
1%
#467240000000
0!
0%
#467245000000
1!
1%
#467250000000
0!
0%
#467255000000
1!
1%
#467260000000
0!
0%
#467265000000
1!
1%
#467270000000
0!
0%
#467275000000
1!
1%
#467280000000
0!
0%
#467285000000
1!
1%
#467290000000
0!
0%
#467295000000
1!
1%
#467300000000
0!
0%
#467305000000
1!
1%
#467310000000
0!
0%
#467315000000
1!
1%
#467320000000
0!
0%
#467325000000
1!
1%
#467330000000
0!
0%
#467335000000
1!
1%
#467340000000
0!
0%
#467345000000
1!
1%
#467350000000
0!
0%
#467355000000
1!
1%
#467360000000
0!
0%
#467365000000
1!
1%
#467370000000
0!
0%
#467375000000
1!
1%
#467380000000
0!
0%
#467385000000
1!
1%
#467390000000
0!
0%
#467395000000
1!
1%
#467400000000
0!
0%
#467405000000
1!
1%
#467410000000
0!
0%
#467415000000
1!
1%
#467420000000
0!
0%
#467425000000
1!
1%
#467430000000
0!
0%
#467435000000
1!
1%
#467440000000
0!
0%
#467445000000
1!
1%
#467450000000
0!
0%
#467455000000
1!
1%
#467460000000
0!
0%
#467465000000
1!
1%
#467470000000
0!
0%
#467475000000
1!
1%
#467480000000
0!
0%
#467485000000
1!
1%
#467490000000
0!
0%
#467495000000
1!
1%
#467500000000
0!
0%
#467505000000
1!
1%
#467510000000
0!
0%
#467515000000
1!
1%
#467520000000
0!
0%
#467525000000
1!
1%
#467530000000
0!
0%
#467535000000
1!
1%
#467540000000
0!
0%
#467545000000
1!
1%
#467550000000
0!
0%
#467555000000
1!
1%
#467560000000
0!
0%
#467565000000
1!
1%
#467570000000
0!
0%
#467575000000
1!
1%
#467580000000
0!
0%
#467585000000
1!
1%
#467590000000
0!
0%
#467595000000
1!
1%
#467600000000
0!
0%
#467605000000
1!
1%
#467610000000
0!
0%
#467615000000
1!
1%
#467620000000
0!
0%
#467625000000
1!
1%
#467630000000
0!
0%
#467635000000
1!
1%
#467640000000
0!
0%
#467645000000
1!
1%
#467650000000
0!
0%
#467655000000
1!
1%
#467660000000
0!
0%
#467665000000
1!
1%
#467670000000
0!
0%
#467675000000
1!
1%
#467680000000
0!
0%
#467685000000
1!
1%
#467690000000
0!
0%
#467695000000
1!
1%
#467700000000
0!
0%
#467705000000
1!
1%
#467710000000
0!
0%
#467715000000
1!
1%
#467720000000
0!
0%
#467725000000
1!
1%
#467730000000
0!
0%
#467735000000
1!
1%
#467740000000
0!
0%
#467745000000
1!
1%
#467750000000
0!
0%
#467755000000
1!
1%
#467760000000
0!
0%
#467765000000
1!
1%
#467770000000
0!
0%
#467775000000
1!
1%
#467780000000
0!
0%
#467785000000
1!
1%
#467790000000
0!
0%
#467795000000
1!
1%
#467800000000
0!
0%
#467805000000
1!
1%
#467810000000
0!
0%
#467815000000
1!
1%
#467820000000
0!
0%
#467825000000
1!
1%
#467830000000
0!
0%
#467835000000
1!
1%
#467840000000
0!
0%
#467845000000
1!
1%
#467850000000
0!
0%
#467855000000
1!
1%
#467860000000
0!
0%
#467865000000
1!
1%
#467870000000
0!
0%
#467875000000
1!
1%
#467880000000
0!
0%
#467885000000
1!
1%
#467890000000
0!
0%
#467895000000
1!
1%
#467900000000
0!
0%
#467905000000
1!
1%
#467910000000
0!
0%
#467915000000
1!
1%
#467920000000
0!
0%
#467925000000
1!
1%
#467930000000
0!
0%
#467935000000
1!
1%
#467940000000
0!
0%
#467945000000
1!
1%
#467950000000
0!
0%
#467955000000
1!
1%
#467960000000
0!
0%
#467965000000
1!
1%
#467970000000
0!
0%
#467975000000
1!
1%
#467980000000
0!
0%
#467985000000
1!
1%
#467990000000
0!
0%
#467995000000
1!
1%
#468000000000
0!
0%
#468005000000
1!
1%
#468010000000
0!
0%
#468015000000
1!
1%
#468020000000
0!
0%
#468025000000
1!
1%
#468030000000
0!
0%
#468035000000
1!
1%
#468040000000
0!
0%
#468045000000
1!
1%
#468050000000
0!
0%
#468055000000
1!
1%
#468060000000
0!
0%
#468065000000
1!
1%
#468070000000
0!
0%
#468075000000
1!
1%
#468080000000
0!
0%
#468085000000
1!
1%
#468090000000
0!
0%
#468095000000
1!
1%
#468100000000
0!
0%
#468105000000
1!
1%
#468110000000
0!
0%
#468115000000
1!
1%
#468120000000
0!
0%
#468125000000
1!
1%
#468130000000
0!
0%
#468135000000
1!
1%
#468140000000
0!
0%
#468145000000
1!
1%
#468150000000
0!
0%
#468155000000
1!
1%
#468160000000
0!
0%
#468165000000
1!
1%
#468170000000
0!
0%
#468175000000
1!
1%
#468180000000
0!
0%
#468185000000
1!
1%
#468190000000
0!
0%
#468195000000
1!
1%
#468200000000
0!
0%
#468205000000
1!
1%
#468210000000
0!
0%
#468215000000
1!
1%
#468220000000
0!
0%
#468225000000
1!
1%
#468230000000
0!
0%
#468235000000
1!
1%
#468240000000
0!
0%
#468245000000
1!
1%
#468250000000
0!
0%
#468255000000
1!
1%
#468260000000
0!
0%
#468265000000
1!
1%
#468270000000
0!
0%
#468275000000
1!
1%
#468280000000
0!
0%
#468285000000
1!
1%
#468290000000
0!
0%
#468295000000
1!
1%
#468300000000
0!
0%
#468305000000
1!
1%
#468310000000
0!
0%
#468315000000
1!
1%
#468320000000
0!
0%
#468325000000
1!
1%
#468330000000
0!
0%
#468335000000
1!
1%
#468340000000
0!
0%
#468345000000
1!
1%
#468350000000
0!
0%
#468355000000
1!
1%
#468360000000
0!
0%
#468365000000
1!
1%
#468370000000
0!
0%
#468375000000
1!
1%
#468380000000
0!
0%
#468385000000
1!
1%
#468390000000
0!
0%
#468395000000
1!
1%
#468400000000
0!
0%
#468405000000
1!
1%
#468410000000
0!
0%
#468415000000
1!
1%
#468420000000
0!
0%
#468425000000
1!
1%
#468430000000
0!
0%
#468435000000
1!
1%
#468440000000
0!
0%
#468445000000
1!
1%
#468450000000
0!
0%
#468455000000
1!
1%
#468460000000
0!
0%
#468465000000
1!
1%
#468470000000
0!
0%
#468475000000
1!
1%
#468480000000
0!
0%
#468485000000
1!
1%
#468490000000
0!
0%
#468495000000
1!
1%
#468500000000
0!
0%
#468505000000
1!
1%
#468510000000
0!
0%
#468515000000
1!
1%
#468520000000
0!
0%
#468525000000
1!
1%
#468530000000
0!
0%
#468535000000
1!
1%
#468540000000
0!
0%
#468545000000
1!
1%
#468550000000
0!
0%
#468555000000
1!
1%
#468560000000
0!
0%
#468565000000
1!
1%
#468570000000
0!
0%
#468575000000
1!
1%
#468580000000
0!
0%
#468585000000
1!
1%
#468590000000
0!
0%
#468595000000
1!
1%
#468600000000
0!
0%
#468605000000
1!
1%
#468610000000
0!
0%
#468615000000
1!
1%
#468620000000
0!
0%
#468625000000
1!
1%
#468630000000
0!
0%
#468635000000
1!
1%
#468640000000
0!
0%
#468645000000
1!
1%
#468650000000
0!
0%
#468655000000
1!
1%
#468660000000
0!
0%
#468665000000
1!
1%
#468670000000
0!
0%
#468675000000
1!
1%
#468680000000
0!
0%
#468685000000
1!
1%
#468690000000
0!
0%
#468695000000
1!
1%
#468700000000
0!
0%
#468705000000
1!
1%
#468710000000
0!
0%
#468715000000
1!
1%
#468720000000
0!
0%
#468725000000
1!
1%
#468730000000
0!
0%
#468735000000
1!
1%
#468740000000
0!
0%
#468745000000
1!
1%
#468750000000
0!
0%
#468755000000
1!
1%
#468760000000
0!
0%
#468765000000
1!
1%
#468770000000
0!
0%
#468775000000
1!
1%
#468780000000
0!
0%
#468785000000
1!
1%
#468790000000
0!
0%
#468795000000
1!
1%
#468800000000
0!
0%
#468805000000
1!
1%
#468810000000
0!
0%
#468815000000
1!
1%
#468820000000
0!
0%
#468825000000
1!
1%
#468830000000
0!
0%
#468835000000
1!
1%
#468840000000
0!
0%
#468845000000
1!
1%
#468850000000
0!
0%
#468855000000
1!
1%
#468860000000
0!
0%
#468865000000
1!
1%
#468870000000
0!
0%
#468875000000
1!
1%
#468880000000
0!
0%
#468885000000
1!
1%
#468890000000
0!
0%
#468895000000
1!
1%
#468900000000
0!
0%
#468905000000
1!
1%
#468910000000
0!
0%
#468915000000
1!
1%
#468920000000
0!
0%
#468925000000
1!
1%
#468930000000
0!
0%
#468935000000
1!
1%
#468940000000
0!
0%
#468945000000
1!
1%
#468950000000
0!
0%
#468955000000
1!
1%
#468960000000
0!
0%
#468965000000
1!
1%
#468970000000
0!
0%
#468975000000
1!
1%
#468980000000
0!
0%
#468985000000
1!
1%
#468990000000
0!
0%
#468995000000
1!
1%
#469000000000
0!
0%
#469005000000
1!
1%
#469010000000
0!
0%
#469015000000
1!
1%
#469020000000
0!
0%
#469025000000
1!
1%
#469030000000
0!
0%
#469035000000
1!
1%
#469040000000
0!
0%
#469045000000
1!
1%
#469050000000
0!
0%
#469055000000
1!
1%
#469060000000
0!
0%
#469065000000
1!
1%
#469070000000
0!
0%
#469075000000
1!
1%
#469080000000
0!
0%
#469085000000
1!
1%
#469090000000
0!
0%
#469095000000
1!
1%
#469100000000
0!
0%
#469105000000
1!
1%
#469110000000
0!
0%
#469115000000
1!
1%
#469120000000
0!
0%
#469125000000
1!
1%
#469130000000
0!
0%
#469135000000
1!
1%
#469140000000
0!
0%
#469145000000
1!
1%
#469150000000
0!
0%
#469155000000
1!
1%
#469160000000
0!
0%
#469165000000
1!
1%
#469170000000
0!
0%
#469175000000
1!
1%
#469180000000
0!
0%
#469185000000
1!
1%
#469190000000
0!
0%
#469195000000
1!
1%
#469200000000
0!
0%
#469205000000
1!
1%
#469210000000
0!
0%
#469215000000
1!
1%
#469220000000
0!
0%
#469225000000
1!
1%
#469230000000
0!
0%
#469235000000
1!
1%
#469240000000
0!
0%
#469245000000
1!
1%
#469250000000
0!
0%
#469255000000
1!
1%
#469260000000
0!
0%
#469265000000
1!
1%
#469270000000
0!
0%
#469275000000
1!
1%
#469280000000
0!
0%
#469285000000
1!
1%
#469290000000
0!
0%
#469295000000
1!
1%
#469300000000
0!
0%
#469305000000
1!
1%
#469310000000
0!
0%
#469315000000
1!
1%
#469320000000
0!
0%
#469325000000
1!
1%
#469330000000
0!
0%
#469335000000
1!
1%
#469340000000
0!
0%
#469345000000
1!
1%
#469350000000
0!
0%
#469355000000
1!
1%
#469360000000
0!
0%
#469365000000
1!
1%
#469370000000
0!
0%
#469375000000
1!
1%
#469380000000
0!
0%
#469385000000
1!
1%
#469390000000
0!
0%
#469395000000
1!
1%
#469400000000
0!
0%
#469405000000
1!
1%
#469410000000
0!
0%
#469415000000
1!
1%
#469420000000
0!
0%
#469425000000
1!
1%
#469430000000
0!
0%
#469435000000
1!
1%
#469440000000
0!
0%
#469445000000
1!
1%
#469450000000
0!
0%
#469455000000
1!
1%
#469460000000
0!
0%
#469465000000
1!
1%
#469470000000
0!
0%
#469475000000
1!
1%
#469480000000
0!
0%
#469485000000
1!
1%
#469490000000
0!
0%
#469495000000
1!
1%
#469500000000
0!
0%
#469505000000
1!
1%
#469510000000
0!
0%
#469515000000
1!
1%
#469520000000
0!
0%
#469525000000
1!
1%
#469530000000
0!
0%
#469535000000
1!
1%
#469540000000
0!
0%
#469545000000
1!
1%
#469550000000
0!
0%
#469555000000
1!
1%
#469560000000
0!
0%
#469565000000
1!
1%
#469570000000
0!
0%
#469575000000
1!
1%
#469580000000
0!
0%
#469585000000
1!
1%
#469590000000
0!
0%
#469595000000
1!
1%
#469600000000
0!
0%
#469605000000
1!
1%
#469610000000
0!
0%
#469615000000
1!
1%
#469620000000
0!
0%
#469625000000
1!
1%
#469630000000
0!
0%
#469635000000
1!
1%
#469640000000
0!
0%
#469645000000
1!
1%
#469650000000
0!
0%
#469655000000
1!
1%
#469660000000
0!
0%
#469665000000
1!
1%
#469670000000
0!
0%
#469675000000
1!
1%
#469680000000
0!
0%
#469685000000
1!
1%
#469690000000
0!
0%
#469695000000
1!
1%
#469700000000
0!
0%
#469705000000
1!
1%
#469710000000
0!
0%
#469715000000
1!
1%
#469720000000
0!
0%
#469725000000
1!
1%
#469730000000
0!
0%
#469735000000
1!
1%
#469740000000
0!
0%
#469745000000
1!
1%
#469750000000
0!
0%
#469755000000
1!
1%
#469760000000
0!
0%
#469765000000
1!
1%
#469770000000
0!
0%
#469775000000
1!
1%
#469780000000
0!
0%
#469785000000
1!
1%
#469790000000
0!
0%
#469795000000
1!
1%
#469800000000
0!
0%
#469805000000
1!
1%
#469810000000
0!
0%
#469815000000
1!
1%
#469820000000
0!
0%
#469825000000
1!
1%
#469830000000
0!
0%
#469835000000
1!
1%
#469840000000
0!
0%
#469845000000
1!
1%
#469850000000
0!
0%
#469855000000
1!
1%
#469860000000
0!
0%
#469865000000
1!
1%
#469870000000
0!
0%
#469875000000
1!
1%
#469880000000
0!
0%
#469885000000
1!
1%
#469890000000
0!
0%
#469895000000
1!
1%
#469900000000
0!
0%
#469905000000
1!
1%
#469910000000
0!
0%
#469915000000
1!
1%
#469920000000
0!
0%
#469925000000
1!
1%
#469930000000
0!
0%
#469935000000
1!
1%
#469940000000
0!
0%
#469945000000
1!
1%
#469950000000
0!
0%
#469955000000
1!
1%
#469960000000
0!
0%
#469965000000
1!
1%
#469970000000
0!
0%
#469975000000
1!
1%
#469980000000
0!
0%
#469985000000
1!
1%
#469990000000
0!
0%
#469995000000
1!
1%
#470000000000
0!
0%
#470005000000
1!
1%
#470010000000
0!
0%
#470015000000
1!
1%
#470020000000
0!
0%
#470025000000
1!
1%
#470030000000
0!
0%
#470035000000
1!
1%
#470040000000
0!
0%
#470045000000
1!
1%
#470050000000
0!
0%
#470055000000
1!
1%
#470060000000
0!
0%
#470065000000
1!
1%
#470070000000
0!
0%
#470075000000
1!
1%
#470080000000
0!
0%
#470085000000
1!
1%
#470090000000
0!
0%
#470095000000
1!
1%
#470100000000
0!
0%
#470105000000
1!
1%
#470110000000
0!
0%
#470115000000
1!
1%
#470120000000
0!
0%
#470125000000
1!
1%
#470130000000
0!
0%
#470135000000
1!
1%
#470140000000
0!
0%
#470145000000
1!
1%
#470150000000
0!
0%
#470155000000
1!
1%
#470160000000
0!
0%
#470165000000
1!
1%
#470170000000
0!
0%
#470175000000
1!
1%
#470180000000
0!
0%
#470185000000
1!
1%
#470190000000
0!
0%
#470195000000
1!
1%
#470200000000
0!
0%
#470205000000
1!
1%
#470210000000
0!
0%
#470215000000
1!
1%
#470220000000
0!
0%
#470225000000
1!
1%
#470230000000
0!
0%
#470235000000
1!
1%
#470240000000
0!
0%
#470245000000
1!
1%
#470250000000
0!
0%
#470255000000
1!
1%
#470260000000
0!
0%
#470265000000
1!
1%
#470270000000
0!
0%
#470275000000
1!
1%
#470280000000
0!
0%
#470285000000
1!
1%
#470290000000
0!
0%
#470295000000
1!
1%
#470300000000
0!
0%
#470305000000
1!
1%
#470310000000
0!
0%
#470315000000
1!
1%
#470320000000
0!
0%
#470325000000
1!
1%
#470330000000
0!
0%
#470335000000
1!
1%
#470340000000
0!
0%
#470345000000
1!
1%
#470350000000
0!
0%
#470355000000
1!
1%
#470360000000
0!
0%
#470365000000
1!
1%
#470370000000
0!
0%
#470375000000
1!
1%
#470380000000
0!
0%
#470385000000
1!
1%
#470390000000
0!
0%
#470395000000
1!
1%
#470400000000
0!
0%
#470405000000
1!
1%
#470410000000
0!
0%
#470415000000
1!
1%
#470420000000
0!
0%
#470425000000
1!
1%
#470430000000
0!
0%
#470435000000
1!
1%
#470440000000
0!
0%
#470445000000
1!
1%
#470450000000
0!
0%
#470455000000
1!
1%
#470460000000
0!
0%
#470465000000
1!
1%
#470470000000
0!
0%
#470475000000
1!
1%
#470480000000
0!
0%
#470485000000
1!
1%
#470490000000
0!
0%
#470495000000
1!
1%
#470500000000
0!
0%
#470505000000
1!
1%
#470510000000
0!
0%
#470515000000
1!
1%
#470520000000
0!
0%
#470525000000
1!
1%
#470530000000
0!
0%
#470535000000
1!
1%
#470540000000
0!
0%
#470545000000
1!
1%
#470550000000
0!
0%
#470555000000
1!
1%
#470560000000
0!
0%
#470565000000
1!
1%
#470570000000
0!
0%
#470575000000
1!
1%
#470580000000
0!
0%
#470585000000
1!
1%
#470590000000
0!
0%
#470595000000
1!
1%
#470600000000
0!
0%
#470605000000
1!
1%
#470610000000
0!
0%
#470615000000
1!
1%
#470620000000
0!
0%
#470625000000
1!
1%
#470630000000
0!
0%
#470635000000
1!
1%
#470640000000
0!
0%
#470645000000
1!
1%
#470650000000
0!
0%
#470655000000
1!
1%
#470660000000
0!
0%
#470665000000
1!
1%
#470670000000
0!
0%
#470675000000
1!
1%
#470680000000
0!
0%
#470685000000
1!
1%
#470690000000
0!
0%
#470695000000
1!
1%
#470700000000
0!
0%
#470705000000
1!
1%
#470710000000
0!
0%
#470715000000
1!
1%
#470720000000
0!
0%
#470725000000
1!
1%
#470730000000
0!
0%
#470735000000
1!
1%
#470740000000
0!
0%
#470745000000
1!
1%
#470750000000
0!
0%
#470755000000
1!
1%
#470760000000
0!
0%
#470765000000
1!
1%
#470770000000
0!
0%
#470775000000
1!
1%
#470780000000
0!
0%
#470785000000
1!
1%
#470790000000
0!
0%
#470795000000
1!
1%
#470800000000
0!
0%
#470805000000
1!
1%
#470810000000
0!
0%
#470815000000
1!
1%
#470820000000
0!
0%
#470825000000
1!
1%
#470830000000
0!
0%
#470835000000
1!
1%
#470840000000
0!
0%
#470845000000
1!
1%
#470850000000
0!
0%
#470855000000
1!
1%
#470860000000
0!
0%
#470865000000
1!
1%
#470870000000
0!
0%
#470875000000
1!
1%
#470880000000
0!
0%
#470885000000
1!
1%
#470890000000
0!
0%
#470895000000
1!
1%
#470900000000
0!
0%
#470905000000
1!
1%
#470910000000
0!
0%
#470915000000
1!
1%
#470920000000
0!
0%
#470925000000
1!
1%
#470930000000
0!
0%
#470935000000
1!
1%
#470940000000
0!
0%
#470945000000
1!
1%
#470950000000
0!
0%
#470955000000
1!
1%
#470960000000
0!
0%
#470965000000
1!
1%
#470970000000
0!
0%
#470975000000
1!
1%
#470980000000
0!
0%
#470985000000
1!
1%
#470990000000
0!
0%
#470995000000
1!
1%
#471000000000
0!
0%
#471005000000
1!
1%
#471010000000
0!
0%
#471015000000
1!
1%
#471020000000
0!
0%
#471025000000
1!
1%
#471030000000
0!
0%
#471035000000
1!
1%
#471040000000
0!
0%
#471045000000
1!
1%
#471050000000
0!
0%
#471055000000
1!
1%
#471060000000
0!
0%
#471065000000
1!
1%
#471070000000
0!
0%
#471075000000
1!
1%
#471080000000
0!
0%
#471085000000
1!
1%
#471090000000
0!
0%
#471095000000
1!
1%
#471100000000
0!
0%
#471105000000
1!
1%
#471110000000
0!
0%
#471115000000
1!
1%
#471120000000
0!
0%
#471125000000
1!
1%
#471130000000
0!
0%
#471135000000
1!
1%
#471140000000
0!
0%
#471145000000
1!
1%
#471150000000
0!
0%
#471155000000
1!
1%
#471160000000
0!
0%
#471165000000
1!
1%
#471170000000
0!
0%
#471175000000
1!
1%
#471180000000
0!
0%
#471185000000
1!
1%
#471190000000
0!
0%
#471195000000
1!
1%
#471200000000
0!
0%
#471205000000
1!
1%
#471210000000
0!
0%
#471215000000
1!
1%
#471220000000
0!
0%
#471225000000
1!
1%
#471230000000
0!
0%
#471235000000
1!
1%
#471240000000
0!
0%
#471245000000
1!
1%
#471250000000
0!
0%
#471255000000
1!
1%
#471260000000
0!
0%
#471265000000
1!
1%
#471270000000
0!
0%
#471275000000
1!
1%
#471280000000
0!
0%
#471285000000
1!
1%
#471290000000
0!
0%
#471295000000
1!
1%
#471300000000
0!
0%
#471305000000
1!
1%
#471310000000
0!
0%
#471315000000
1!
1%
#471320000000
0!
0%
#471325000000
1!
1%
#471330000000
0!
0%
#471335000000
1!
1%
#471340000000
0!
0%
#471345000000
1!
1%
#471350000000
0!
0%
#471355000000
1!
1%
#471360000000
0!
0%
#471365000000
1!
1%
#471370000000
0!
0%
#471375000000
1!
1%
#471380000000
0!
0%
#471385000000
1!
1%
#471390000000
0!
0%
#471395000000
1!
1%
#471400000000
0!
0%
#471405000000
1!
1%
#471410000000
0!
0%
#471415000000
1!
1%
#471420000000
0!
0%
#471425000000
1!
1%
#471430000000
0!
0%
#471435000000
1!
1%
#471440000000
0!
0%
#471445000000
1!
1%
#471450000000
0!
0%
#471455000000
1!
1%
#471460000000
0!
0%
#471465000000
1!
1%
#471470000000
0!
0%
#471475000000
1!
1%
#471480000000
0!
0%
#471485000000
1!
1%
#471490000000
0!
0%
#471495000000
1!
1%
#471500000000
0!
0%
#471505000000
1!
1%
#471510000000
0!
0%
#471515000000
1!
1%
#471520000000
0!
0%
#471525000000
1!
1%
#471530000000
0!
0%
#471535000000
1!
1%
#471540000000
0!
0%
#471545000000
1!
1%
#471550000000
0!
0%
#471555000000
1!
1%
#471560000000
0!
0%
#471565000000
1!
1%
#471570000000
0!
0%
#471575000000
1!
1%
#471580000000
0!
0%
#471585000000
1!
1%
#471590000000
0!
0%
#471595000000
1!
1%
#471600000000
0!
0%
#471605000000
1!
1%
#471610000000
0!
0%
#471615000000
1!
1%
#471620000000
0!
0%
#471625000000
1!
1%
#471630000000
0!
0%
#471635000000
1!
1%
#471640000000
0!
0%
#471645000000
1!
1%
#471650000000
0!
0%
#471655000000
1!
1%
#471660000000
0!
0%
#471665000000
1!
1%
#471670000000
0!
0%
#471675000000
1!
1%
#471680000000
0!
0%
#471685000000
1!
1%
#471690000000
0!
0%
#471695000000
1!
1%
#471700000000
0!
0%
#471705000000
1!
1%
#471710000000
0!
0%
#471715000000
1!
1%
#471720000000
0!
0%
#471725000000
1!
1%
#471730000000
0!
0%
#471735000000
1!
1%
#471740000000
0!
0%
#471745000000
1!
1%
#471750000000
0!
0%
#471755000000
1!
1%
#471760000000
0!
0%
#471765000000
1!
1%
#471770000000
0!
0%
#471775000000
1!
1%
#471780000000
0!
0%
#471785000000
1!
1%
#471790000000
0!
0%
#471795000000
1!
1%
#471800000000
0!
0%
#471805000000
1!
1%
#471810000000
0!
0%
#471815000000
1!
1%
#471820000000
0!
0%
#471825000000
1!
1%
#471830000000
0!
0%
#471835000000
1!
1%
#471840000000
0!
0%
#471845000000
1!
1%
#471850000000
0!
0%
#471855000000
1!
1%
#471860000000
0!
0%
#471865000000
1!
1%
#471870000000
0!
0%
#471875000000
1!
1%
#471880000000
0!
0%
#471885000000
1!
1%
#471890000000
0!
0%
#471895000000
1!
1%
#471900000000
0!
0%
#471905000000
1!
1%
#471910000000
0!
0%
#471915000000
1!
1%
#471920000000
0!
0%
#471925000000
1!
1%
#471930000000
0!
0%
#471935000000
1!
1%
#471940000000
0!
0%
#471945000000
1!
1%
#471950000000
0!
0%
#471955000000
1!
1%
#471960000000
0!
0%
#471965000000
1!
1%
#471970000000
0!
0%
#471975000000
1!
1%
#471980000000
0!
0%
#471985000000
1!
1%
#471990000000
0!
0%
#471995000000
1!
1%
#472000000000
0!
0%
#472005000000
1!
1%
#472010000000
0!
0%
#472015000000
1!
1%
#472020000000
0!
0%
#472025000000
1!
1%
#472030000000
0!
0%
#472035000000
1!
1%
#472040000000
0!
0%
#472045000000
1!
1%
#472050000000
0!
0%
#472055000000
1!
1%
#472060000000
0!
0%
#472065000000
1!
1%
#472070000000
0!
0%
#472075000000
1!
1%
#472080000000
0!
0%
#472085000000
1!
1%
#472090000000
0!
0%
#472095000000
1!
1%
#472100000000
0!
0%
#472105000000
1!
1%
#472110000000
0!
0%
#472115000000
1!
1%
#472120000000
0!
0%
#472125000000
1!
1%
#472130000000
0!
0%
#472135000000
1!
1%
#472140000000
0!
0%
#472145000000
1!
1%
#472150000000
0!
0%
#472155000000
1!
1%
#472160000000
0!
0%
#472165000000
1!
1%
#472170000000
0!
0%
#472175000000
1!
1%
#472180000000
0!
0%
#472185000000
1!
1%
#472190000000
0!
0%
#472195000000
1!
1%
#472200000000
0!
0%
#472205000000
1!
1%
#472210000000
0!
0%
#472215000000
1!
1%
#472220000000
0!
0%
#472225000000
1!
1%
#472230000000
0!
0%
#472235000000
1!
1%
#472240000000
0!
0%
#472245000000
1!
1%
#472250000000
0!
0%
#472255000000
1!
1%
#472260000000
0!
0%
#472265000000
1!
1%
#472270000000
0!
0%
#472275000000
1!
1%
#472280000000
0!
0%
#472285000000
1!
1%
#472290000000
0!
0%
#472295000000
1!
1%
#472300000000
0!
0%
#472305000000
1!
1%
#472310000000
0!
0%
#472315000000
1!
1%
#472320000000
0!
0%
#472325000000
1!
1%
#472330000000
0!
0%
#472335000000
1!
1%
#472340000000
0!
0%
#472345000000
1!
1%
#472350000000
0!
0%
#472355000000
1!
1%
#472360000000
0!
0%
#472365000000
1!
1%
#472370000000
0!
0%
#472375000000
1!
1%
#472380000000
0!
0%
#472385000000
1!
1%
#472390000000
0!
0%
#472395000000
1!
1%
#472400000000
0!
0%
#472405000000
1!
1%
#472410000000
0!
0%
#472415000000
1!
1%
#472420000000
0!
0%
#472425000000
1!
1%
#472430000000
0!
0%
#472435000000
1!
1%
#472440000000
0!
0%
#472445000000
1!
1%
#472450000000
0!
0%
#472455000000
1!
1%
#472460000000
0!
0%
#472465000000
1!
1%
#472470000000
0!
0%
#472475000000
1!
1%
#472480000000
0!
0%
#472485000000
1!
1%
#472490000000
0!
0%
#472495000000
1!
1%
#472500000000
0!
0%
#472505000000
1!
1%
#472510000000
0!
0%
#472515000000
1!
1%
#472520000000
0!
0%
#472525000000
1!
1%
#472530000000
0!
0%
#472535000000
1!
1%
#472540000000
0!
0%
#472545000000
1!
1%
#472550000000
0!
0%
#472555000000
1!
1%
#472560000000
0!
0%
#472565000000
1!
1%
#472570000000
0!
0%
#472575000000
1!
1%
#472580000000
0!
0%
#472585000000
1!
1%
#472590000000
0!
0%
#472595000000
1!
1%
#472600000000
0!
0%
#472605000000
1!
1%
#472610000000
0!
0%
#472615000000
1!
1%
#472620000000
0!
0%
#472625000000
1!
1%
#472630000000
0!
0%
#472635000000
1!
1%
#472640000000
0!
0%
#472645000000
1!
1%
#472650000000
0!
0%
#472655000000
1!
1%
#472660000000
0!
0%
#472665000000
1!
1%
#472670000000
0!
0%
#472675000000
1!
1%
#472680000000
0!
0%
#472685000000
1!
1%
#472690000000
0!
0%
#472695000000
1!
1%
#472700000000
0!
0%
#472705000000
1!
1%
#472710000000
0!
0%
#472715000000
1!
1%
#472720000000
0!
0%
#472725000000
1!
1%
#472730000000
0!
0%
#472735000000
1!
1%
#472740000000
0!
0%
#472745000000
1!
1%
#472750000000
0!
0%
#472755000000
1!
1%
#472760000000
0!
0%
#472765000000
1!
1%
#472770000000
0!
0%
#472775000000
1!
1%
#472780000000
0!
0%
#472785000000
1!
1%
#472790000000
0!
0%
#472795000000
1!
1%
#472800000000
0!
0%
#472805000000
1!
1%
#472810000000
0!
0%
#472815000000
1!
1%
#472820000000
0!
0%
#472825000000
1!
1%
#472830000000
0!
0%
#472835000000
1!
1%
#472840000000
0!
0%
#472845000000
1!
1%
#472850000000
0!
0%
#472855000000
1!
1%
#472860000000
0!
0%
#472865000000
1!
1%
#472870000000
0!
0%
#472875000000
1!
1%
#472880000000
0!
0%
#472885000000
1!
1%
#472890000000
0!
0%
#472895000000
1!
1%
#472900000000
0!
0%
#472905000000
1!
1%
#472910000000
0!
0%
#472915000000
1!
1%
#472920000000
0!
0%
#472925000000
1!
1%
#472930000000
0!
0%
#472935000000
1!
1%
#472940000000
0!
0%
#472945000000
1!
1%
#472950000000
0!
0%
#472955000000
1!
1%
#472960000000
0!
0%
#472965000000
1!
1%
#472970000000
0!
0%
#472975000000
1!
1%
#472980000000
0!
0%
#472985000000
1!
1%
#472990000000
0!
0%
#472995000000
1!
1%
#473000000000
0!
0%
#473005000000
1!
1%
#473010000000
0!
0%
#473015000000
1!
1%
#473020000000
0!
0%
#473025000000
1!
1%
#473030000000
0!
0%
#473035000000
1!
1%
#473040000000
0!
0%
#473045000000
1!
1%
#473050000000
0!
0%
#473055000000
1!
1%
#473060000000
0!
0%
#473065000000
1!
1%
#473070000000
0!
0%
#473075000000
1!
1%
#473080000000
0!
0%
#473085000000
1!
1%
#473090000000
0!
0%
#473095000000
1!
1%
#473100000000
0!
0%
#473105000000
1!
1%
#473110000000
0!
0%
#473115000000
1!
1%
#473120000000
0!
0%
#473125000000
1!
1%
#473130000000
0!
0%
#473135000000
1!
1%
#473140000000
0!
0%
#473145000000
1!
1%
#473150000000
0!
0%
#473155000000
1!
1%
#473160000000
0!
0%
#473165000000
1!
1%
#473170000000
0!
0%
#473175000000
1!
1%
#473180000000
0!
0%
#473185000000
1!
1%
#473190000000
0!
0%
#473195000000
1!
1%
#473200000000
0!
0%
#473205000000
1!
1%
#473210000000
0!
0%
#473215000000
1!
1%
#473220000000
0!
0%
#473225000000
1!
1%
#473230000000
0!
0%
#473235000000
1!
1%
#473240000000
0!
0%
#473245000000
1!
1%
#473250000000
0!
0%
#473255000000
1!
1%
#473260000000
0!
0%
#473265000000
1!
1%
#473270000000
0!
0%
#473275000000
1!
1%
#473280000000
0!
0%
#473285000000
1!
1%
#473290000000
0!
0%
#473295000000
1!
1%
#473300000000
0!
0%
#473305000000
1!
1%
#473310000000
0!
0%
#473315000000
1!
1%
#473320000000
0!
0%
#473325000000
1!
1%
#473330000000
0!
0%
#473335000000
1!
1%
#473340000000
0!
0%
#473345000000
1!
1%
#473350000000
0!
0%
#473355000000
1!
1%
#473360000000
0!
0%
#473365000000
1!
1%
#473370000000
0!
0%
#473375000000
1!
1%
#473380000000
0!
0%
#473385000000
1!
1%
#473390000000
0!
0%
#473395000000
1!
1%
#473400000000
0!
0%
#473405000000
1!
1%
#473410000000
0!
0%
#473415000000
1!
1%
#473420000000
0!
0%
#473425000000
1!
1%
#473430000000
0!
0%
#473435000000
1!
1%
#473440000000
0!
0%
#473445000000
1!
1%
#473450000000
0!
0%
#473455000000
1!
1%
#473460000000
0!
0%
#473465000000
1!
1%
#473470000000
0!
0%
#473475000000
1!
1%
#473480000000
0!
0%
#473485000000
1!
1%
#473490000000
0!
0%
#473495000000
1!
1%
#473500000000
0!
0%
#473505000000
1!
1%
#473510000000
0!
0%
#473515000000
1!
1%
#473520000000
0!
0%
#473525000000
1!
1%
#473530000000
0!
0%
#473535000000
1!
1%
#473540000000
0!
0%
#473545000000
1!
1%
#473550000000
0!
0%
#473555000000
1!
1%
#473560000000
0!
0%
#473565000000
1!
1%
#473570000000
0!
0%
#473575000000
1!
1%
#473580000000
0!
0%
#473585000000
1!
1%
#473590000000
0!
0%
#473595000000
1!
1%
#473600000000
0!
0%
#473605000000
1!
1%
#473610000000
0!
0%
#473615000000
1!
1%
#473620000000
0!
0%
#473625000000
1!
1%
#473630000000
0!
0%
#473635000000
1!
1%
#473640000000
0!
0%
#473645000000
1!
1%
#473650000000
0!
0%
#473655000000
1!
1%
#473660000000
0!
0%
#473665000000
1!
1%
#473670000000
0!
0%
#473675000000
1!
1%
#473680000000
0!
0%
#473685000000
1!
1%
#473690000000
0!
0%
#473695000000
1!
1%
#473700000000
0!
0%
#473705000000
1!
1%
#473710000000
0!
0%
#473715000000
1!
1%
#473720000000
0!
0%
#473725000000
1!
1%
#473730000000
0!
0%
#473735000000
1!
1%
#473740000000
0!
0%
#473745000000
1!
1%
#473750000000
0!
0%
#473755000000
1!
1%
#473760000000
0!
0%
#473765000000
1!
1%
#473770000000
0!
0%
#473775000000
1!
1%
#473780000000
0!
0%
#473785000000
1!
1%
#473790000000
0!
0%
#473795000000
1!
1%
#473800000000
0!
0%
#473805000000
1!
1%
#473810000000
0!
0%
#473815000000
1!
1%
#473820000000
0!
0%
#473825000000
1!
1%
#473830000000
0!
0%
#473835000000
1!
1%
#473840000000
0!
0%
#473845000000
1!
1%
#473850000000
0!
0%
#473855000000
1!
1%
#473860000000
0!
0%
#473865000000
1!
1%
#473870000000
0!
0%
#473875000000
1!
1%
#473880000000
0!
0%
#473885000000
1!
1%
#473890000000
0!
0%
#473895000000
1!
1%
#473900000000
0!
0%
#473905000000
1!
1%
#473910000000
0!
0%
#473915000000
1!
1%
#473920000000
0!
0%
#473925000000
1!
1%
#473930000000
0!
0%
#473935000000
1!
1%
#473940000000
0!
0%
#473945000000
1!
1%
#473950000000
0!
0%
#473955000000
1!
1%
#473960000000
0!
0%
#473965000000
1!
1%
#473970000000
0!
0%
#473975000000
1!
1%
#473980000000
0!
0%
#473985000000
1!
1%
#473990000000
0!
0%
#473995000000
1!
1%
#474000000000
0!
0%
#474005000000
1!
1%
#474010000000
0!
0%
#474015000000
1!
1%
#474020000000
0!
0%
#474025000000
1!
1%
#474030000000
0!
0%
#474035000000
1!
1%
#474040000000
0!
0%
#474045000000
1!
1%
#474050000000
0!
0%
#474055000000
1!
1%
#474060000000
0!
0%
#474065000000
1!
1%
#474070000000
0!
0%
#474075000000
1!
1%
#474080000000
0!
0%
#474085000000
1!
1%
#474090000000
0!
0%
#474095000000
1!
1%
#474100000000
0!
0%
#474105000000
1!
1%
#474110000000
0!
0%
#474115000000
1!
1%
#474120000000
0!
0%
#474125000000
1!
1%
#474130000000
0!
0%
#474135000000
1!
1%
#474140000000
0!
0%
#474145000000
1!
1%
#474150000000
0!
0%
#474155000000
1!
1%
#474160000000
0!
0%
#474165000000
1!
1%
#474170000000
0!
0%
#474175000000
1!
1%
#474180000000
0!
0%
#474185000000
1!
1%
#474190000000
0!
0%
#474195000000
1!
1%
#474200000000
0!
0%
#474205000000
1!
1%
#474210000000
0!
0%
#474215000000
1!
1%
#474220000000
0!
0%
#474225000000
1!
1%
#474230000000
0!
0%
#474235000000
1!
1%
#474240000000
0!
0%
#474245000000
1!
1%
#474250000000
0!
0%
#474255000000
1!
1%
#474260000000
0!
0%
#474265000000
1!
1%
#474270000000
0!
0%
#474275000000
1!
1%
#474280000000
0!
0%
#474285000000
1!
1%
#474290000000
0!
0%
#474295000000
1!
1%
#474300000000
0!
0%
#474305000000
1!
1%
#474310000000
0!
0%
#474315000000
1!
1%
#474320000000
0!
0%
#474325000000
1!
1%
#474330000000
0!
0%
#474335000000
1!
1%
#474340000000
0!
0%
#474345000000
1!
1%
#474350000000
0!
0%
#474355000000
1!
1%
#474360000000
0!
0%
#474365000000
1!
1%
#474370000000
0!
0%
#474375000000
1!
1%
#474380000000
0!
0%
#474385000000
1!
1%
#474390000000
0!
0%
#474395000000
1!
1%
#474400000000
0!
0%
#474405000000
1!
1%
#474410000000
0!
0%
#474415000000
1!
1%
#474420000000
0!
0%
#474425000000
1!
1%
#474430000000
0!
0%
#474435000000
1!
1%
#474440000000
0!
0%
#474445000000
1!
1%
#474450000000
0!
0%
#474455000000
1!
1%
#474460000000
0!
0%
#474465000000
1!
1%
#474470000000
0!
0%
#474475000000
1!
1%
#474480000000
0!
0%
#474485000000
1!
1%
#474490000000
0!
0%
#474495000000
1!
1%
#474500000000
0!
0%
#474505000000
1!
1%
#474510000000
0!
0%
#474515000000
1!
1%
#474520000000
0!
0%
#474525000000
1!
1%
#474530000000
0!
0%
#474535000000
1!
1%
#474540000000
0!
0%
#474545000000
1!
1%
#474550000000
0!
0%
#474555000000
1!
1%
#474560000000
0!
0%
#474565000000
1!
1%
#474570000000
0!
0%
#474575000000
1!
1%
#474580000000
0!
0%
#474585000000
1!
1%
#474590000000
0!
0%
#474595000000
1!
1%
#474600000000
0!
0%
#474605000000
1!
1%
#474610000000
0!
0%
#474615000000
1!
1%
#474620000000
0!
0%
#474625000000
1!
1%
#474630000000
0!
0%
#474635000000
1!
1%
#474640000000
0!
0%
#474645000000
1!
1%
#474650000000
0!
0%
#474655000000
1!
1%
#474660000000
0!
0%
#474665000000
1!
1%
#474670000000
0!
0%
#474675000000
1!
1%
#474680000000
0!
0%
#474685000000
1!
1%
#474690000000
0!
0%
#474695000000
1!
1%
#474700000000
0!
0%
#474705000000
1!
1%
#474710000000
0!
0%
#474715000000
1!
1%
#474720000000
0!
0%
#474725000000
1!
1%
#474730000000
0!
0%
#474735000000
1!
1%
#474740000000
0!
0%
#474745000000
1!
1%
#474750000000
0!
0%
#474755000000
1!
1%
#474760000000
0!
0%
#474765000000
1!
1%
#474770000000
0!
0%
#474775000000
1!
1%
#474780000000
0!
0%
#474785000000
1!
1%
#474790000000
0!
0%
#474795000000
1!
1%
#474800000000
0!
0%
#474805000000
1!
1%
#474810000000
0!
0%
#474815000000
1!
1%
#474820000000
0!
0%
#474825000000
1!
1%
#474830000000
0!
0%
#474835000000
1!
1%
#474840000000
0!
0%
#474845000000
1!
1%
#474850000000
0!
0%
#474855000000
1!
1%
#474860000000
0!
0%
#474865000000
1!
1%
#474870000000
0!
0%
#474875000000
1!
1%
#474880000000
0!
0%
#474885000000
1!
1%
#474890000000
0!
0%
#474895000000
1!
1%
#474900000000
0!
0%
#474905000000
1!
1%
#474910000000
0!
0%
#474915000000
1!
1%
#474920000000
0!
0%
#474925000000
1!
1%
#474930000000
0!
0%
#474935000000
1!
1%
#474940000000
0!
0%
#474945000000
1!
1%
#474950000000
0!
0%
#474955000000
1!
1%
#474960000000
0!
0%
#474965000000
1!
1%
#474970000000
0!
0%
#474975000000
1!
1%
#474980000000
0!
0%
#474985000000
1!
1%
#474990000000
0!
0%
#474995000000
1!
1%
#475000000000
0!
0%
#475005000000
1!
1%
#475010000000
0!
0%
#475015000000
1!
1%
#475020000000
0!
0%
#475025000000
1!
1%
#475030000000
0!
0%
#475035000000
1!
1%
#475040000000
0!
0%
#475045000000
1!
1%
#475050000000
0!
0%
#475055000000
1!
1%
#475060000000
0!
0%
#475065000000
1!
1%
#475070000000
0!
0%
#475075000000
1!
1%
#475080000000
0!
0%
#475085000000
1!
1%
#475090000000
0!
0%
#475095000000
1!
1%
#475100000000
0!
0%
#475105000000
1!
1%
#475110000000
0!
0%
#475115000000
1!
1%
#475120000000
0!
0%
#475125000000
1!
1%
#475130000000
0!
0%
#475135000000
1!
1%
#475140000000
0!
0%
#475145000000
1!
1%
#475150000000
0!
0%
#475155000000
1!
1%
#475160000000
0!
0%
#475165000000
1!
1%
#475170000000
0!
0%
#475175000000
1!
1%
#475180000000
0!
0%
#475185000000
1!
1%
#475190000000
0!
0%
#475195000000
1!
1%
#475200000000
0!
0%
#475205000000
1!
1%
#475210000000
0!
0%
#475215000000
1!
1%
#475220000000
0!
0%
#475225000000
1!
1%
#475230000000
0!
0%
#475235000000
1!
1%
#475240000000
0!
0%
#475245000000
1!
1%
#475250000000
0!
0%
#475255000000
1!
1%
#475260000000
0!
0%
#475265000000
1!
1%
#475270000000
0!
0%
#475275000000
1!
1%
#475280000000
0!
0%
#475285000000
1!
1%
#475290000000
0!
0%
#475295000000
1!
1%
#475300000000
0!
0%
#475305000000
1!
1%
#475310000000
0!
0%
#475315000000
1!
1%
#475320000000
0!
0%
#475325000000
1!
1%
#475330000000
0!
0%
#475335000000
1!
1%
#475340000000
0!
0%
#475345000000
1!
1%
#475350000000
0!
0%
#475355000000
1!
1%
#475360000000
0!
0%
#475365000000
1!
1%
#475370000000
0!
0%
#475375000000
1!
1%
#475380000000
0!
0%
#475385000000
1!
1%
#475390000000
0!
0%
#475395000000
1!
1%
#475400000000
0!
0%
#475405000000
1!
1%
#475410000000
0!
0%
#475415000000
1!
1%
#475420000000
0!
0%
#475425000000
1!
1%
#475430000000
0!
0%
#475435000000
1!
1%
#475440000000
0!
0%
#475445000000
1!
1%
#475450000000
0!
0%
#475455000000
1!
1%
#475460000000
0!
0%
#475465000000
1!
1%
#475470000000
0!
0%
#475475000000
1!
1%
#475480000000
0!
0%
#475485000000
1!
1%
#475490000000
0!
0%
#475495000000
1!
1%
#475500000000
0!
0%
#475505000000
1!
1%
#475510000000
0!
0%
#475515000000
1!
1%
#475520000000
0!
0%
#475525000000
1!
1%
#475530000000
0!
0%
#475535000000
1!
1%
#475540000000
0!
0%
#475545000000
1!
1%
#475550000000
0!
0%
#475555000000
1!
1%
#475560000000
0!
0%
#475565000000
1!
1%
#475570000000
0!
0%
#475575000000
1!
1%
#475580000000
0!
0%
#475585000000
1!
1%
#475590000000
0!
0%
#475595000000
1!
1%
#475600000000
0!
0%
#475605000000
1!
1%
#475610000000
0!
0%
#475615000000
1!
1%
#475620000000
0!
0%
#475625000000
1!
1%
#475630000000
0!
0%
#475635000000
1!
1%
#475640000000
0!
0%
#475645000000
1!
1%
#475650000000
0!
0%
#475655000000
1!
1%
#475660000000
0!
0%
#475665000000
1!
1%
#475670000000
0!
0%
#475675000000
1!
1%
#475680000000
0!
0%
#475685000000
1!
1%
#475690000000
0!
0%
#475695000000
1!
1%
#475700000000
0!
0%
#475705000000
1!
1%
#475710000000
0!
0%
#475715000000
1!
1%
#475720000000
0!
0%
#475725000000
1!
1%
#475730000000
0!
0%
#475735000000
1!
1%
#475740000000
0!
0%
#475745000000
1!
1%
#475750000000
0!
0%
#475755000000
1!
1%
#475760000000
0!
0%
#475765000000
1!
1%
#475770000000
0!
0%
#475775000000
1!
1%
#475780000000
0!
0%
#475785000000
1!
1%
#475790000000
0!
0%
#475795000000
1!
1%
#475800000000
0!
0%
#475805000000
1!
1%
#475810000000
0!
0%
#475815000000
1!
1%
#475820000000
0!
0%
#475825000000
1!
1%
#475830000000
0!
0%
#475835000000
1!
1%
#475840000000
0!
0%
#475845000000
1!
1%
#475850000000
0!
0%
#475855000000
1!
1%
#475860000000
0!
0%
#475865000000
1!
1%
#475870000000
0!
0%
#475875000000
1!
1%
#475880000000
0!
0%
#475885000000
1!
1%
#475890000000
0!
0%
#475895000000
1!
1%
#475900000000
0!
0%
#475905000000
1!
1%
#475910000000
0!
0%
#475915000000
1!
1%
#475920000000
0!
0%
#475925000000
1!
1%
#475930000000
0!
0%
#475935000000
1!
1%
#475940000000
0!
0%
#475945000000
1!
1%
#475950000000
0!
0%
#475955000000
1!
1%
#475960000000
0!
0%
#475965000000
1!
1%
#475970000000
0!
0%
#475975000000
1!
1%
#475980000000
0!
0%
#475985000000
1!
1%
#475990000000
0!
0%
#475995000000
1!
1%
#476000000000
0!
0%
#476005000000
1!
1%
#476010000000
0!
0%
#476015000000
1!
1%
#476020000000
0!
0%
#476025000000
1!
1%
#476030000000
0!
0%
#476035000000
1!
1%
#476040000000
0!
0%
#476045000000
1!
1%
#476050000000
0!
0%
#476055000000
1!
1%
#476060000000
0!
0%
#476065000000
1!
1%
#476070000000
0!
0%
#476075000000
1!
1%
#476080000000
0!
0%
#476085000000
1!
1%
#476090000000
0!
0%
#476095000000
1!
1%
#476100000000
0!
0%
#476105000000
1!
1%
#476110000000
0!
0%
#476115000000
1!
1%
#476120000000
0!
0%
#476125000000
1!
1%
#476130000000
0!
0%
#476135000000
1!
1%
#476140000000
0!
0%
#476145000000
1!
1%
#476150000000
0!
0%
#476155000000
1!
1%
#476160000000
0!
0%
#476165000000
1!
1%
#476170000000
0!
0%
#476175000000
1!
1%
#476180000000
0!
0%
#476185000000
1!
1%
#476190000000
0!
0%
#476195000000
1!
1%
#476200000000
0!
0%
#476205000000
1!
1%
#476210000000
0!
0%
#476215000000
1!
1%
#476220000000
0!
0%
#476225000000
1!
1%
#476230000000
0!
0%
#476235000000
1!
1%
#476240000000
0!
0%
#476245000000
1!
1%
#476250000000
0!
0%
#476255000000
1!
1%
#476260000000
0!
0%
#476265000000
1!
1%
#476270000000
0!
0%
#476275000000
1!
1%
#476280000000
0!
0%
#476285000000
1!
1%
#476290000000
0!
0%
#476295000000
1!
1%
#476300000000
0!
0%
#476305000000
1!
1%
#476310000000
0!
0%
#476315000000
1!
1%
#476320000000
0!
0%
#476325000000
1!
1%
#476330000000
0!
0%
#476335000000
1!
1%
#476340000000
0!
0%
#476345000000
1!
1%
#476350000000
0!
0%
#476355000000
1!
1%
#476360000000
0!
0%
#476365000000
1!
1%
#476370000000
0!
0%
#476375000000
1!
1%
#476380000000
0!
0%
#476385000000
1!
1%
#476390000000
0!
0%
#476395000000
1!
1%
#476400000000
0!
0%
#476405000000
1!
1%
#476410000000
0!
0%
#476415000000
1!
1%
#476420000000
0!
0%
#476425000000
1!
1%
#476430000000
0!
0%
#476435000000
1!
1%
#476440000000
0!
0%
#476445000000
1!
1%
#476450000000
0!
0%
#476455000000
1!
1%
#476460000000
0!
0%
#476465000000
1!
1%
#476470000000
0!
0%
#476475000000
1!
1%
#476480000000
0!
0%
#476485000000
1!
1%
#476490000000
0!
0%
#476495000000
1!
1%
#476500000000
0!
0%
#476505000000
1!
1%
#476510000000
0!
0%
#476515000000
1!
1%
#476520000000
0!
0%
#476525000000
1!
1%
#476530000000
0!
0%
#476535000000
1!
1%
#476540000000
0!
0%
#476545000000
1!
1%
#476550000000
0!
0%
#476555000000
1!
1%
#476560000000
0!
0%
#476565000000
1!
1%
#476570000000
0!
0%
#476575000000
1!
1%
#476580000000
0!
0%
#476585000000
1!
1%
#476590000000
0!
0%
#476595000000
1!
1%
#476600000000
0!
0%
#476605000000
1!
1%
#476610000000
0!
0%
#476615000000
1!
1%
#476620000000
0!
0%
#476625000000
1!
1%
#476630000000
0!
0%
#476635000000
1!
1%
#476640000000
0!
0%
#476645000000
1!
1%
#476650000000
0!
0%
#476655000000
1!
1%
#476660000000
0!
0%
#476665000000
1!
1%
#476670000000
0!
0%
#476675000000
1!
1%
#476680000000
0!
0%
#476685000000
1!
1%
#476690000000
0!
0%
#476695000000
1!
1%
#476700000000
0!
0%
#476705000000
1!
1%
#476710000000
0!
0%
#476715000000
1!
1%
#476720000000
0!
0%
#476725000000
1!
1%
#476730000000
0!
0%
#476735000000
1!
1%
#476740000000
0!
0%
#476745000000
1!
1%
#476750000000
0!
0%
#476755000000
1!
1%
#476760000000
0!
0%
#476765000000
1!
1%
#476770000000
0!
0%
#476775000000
1!
1%
#476780000000
0!
0%
#476785000000
1!
1%
#476790000000
0!
0%
#476795000000
1!
1%
#476800000000
0!
0%
#476805000000
1!
1%
#476810000000
0!
0%
#476815000000
1!
1%
#476820000000
0!
0%
#476825000000
1!
1%
#476830000000
0!
0%
#476835000000
1!
1%
#476840000000
0!
0%
#476845000000
1!
1%
#476850000000
0!
0%
#476855000000
1!
1%
#476860000000
0!
0%
#476865000000
1!
1%
#476870000000
0!
0%
#476875000000
1!
1%
#476880000000
0!
0%
#476885000000
1!
1%
#476890000000
0!
0%
#476895000000
1!
1%
#476900000000
0!
0%
#476905000000
1!
1%
#476910000000
0!
0%
#476915000000
1!
1%
#476920000000
0!
0%
#476925000000
1!
1%
#476930000000
0!
0%
#476935000000
1!
1%
#476940000000
0!
0%
#476945000000
1!
1%
#476950000000
0!
0%
#476955000000
1!
1%
#476960000000
0!
0%
#476965000000
1!
1%
#476970000000
0!
0%
#476975000000
1!
1%
#476980000000
0!
0%
#476985000000
1!
1%
#476990000000
0!
0%
#476995000000
1!
1%
#477000000000
0!
0%
#477005000000
1!
1%
#477010000000
0!
0%
#477015000000
1!
1%
#477020000000
0!
0%
#477025000000
1!
1%
#477030000000
0!
0%
#477035000000
1!
1%
#477040000000
0!
0%
#477045000000
1!
1%
#477050000000
0!
0%
#477055000000
1!
1%
#477060000000
0!
0%
#477065000000
1!
1%
#477070000000
0!
0%
#477075000000
1!
1%
#477080000000
0!
0%
#477085000000
1!
1%
#477090000000
0!
0%
#477095000000
1!
1%
#477100000000
0!
0%
#477105000000
1!
1%
#477110000000
0!
0%
#477115000000
1!
1%
#477120000000
0!
0%
#477125000000
1!
1%
#477130000000
0!
0%
#477135000000
1!
1%
#477140000000
0!
0%
#477145000000
1!
1%
#477150000000
0!
0%
#477155000000
1!
1%
#477160000000
0!
0%
#477165000000
1!
1%
#477170000000
0!
0%
#477175000000
1!
1%
#477180000000
0!
0%
#477185000000
1!
1%
#477190000000
0!
0%
#477195000000
1!
1%
#477200000000
0!
0%
#477205000000
1!
1%
#477210000000
0!
0%
#477215000000
1!
1%
#477220000000
0!
0%
#477225000000
1!
1%
#477230000000
0!
0%
#477235000000
1!
1%
#477240000000
0!
0%
#477245000000
1!
1%
#477250000000
0!
0%
#477255000000
1!
1%
#477260000000
0!
0%
#477265000000
1!
1%
#477270000000
0!
0%
#477275000000
1!
1%
#477280000000
0!
0%
#477285000000
1!
1%
#477290000000
0!
0%
#477295000000
1!
1%
#477300000000
0!
0%
#477305000000
1!
1%
#477310000000
0!
0%
#477315000000
1!
1%
#477320000000
0!
0%
#477325000000
1!
1%
#477330000000
0!
0%
#477335000000
1!
1%
#477340000000
0!
0%
#477345000000
1!
1%
#477350000000
0!
0%
#477355000000
1!
1%
#477360000000
0!
0%
#477365000000
1!
1%
#477370000000
0!
0%
#477375000000
1!
1%
#477380000000
0!
0%
#477385000000
1!
1%
#477390000000
0!
0%
#477395000000
1!
1%
#477400000000
0!
0%
#477405000000
1!
1%
#477410000000
0!
0%
#477415000000
1!
1%
#477420000000
0!
0%
#477425000000
1!
1%
#477430000000
0!
0%
#477435000000
1!
1%
#477440000000
0!
0%
#477445000000
1!
1%
#477450000000
0!
0%
#477455000000
1!
1%
#477460000000
0!
0%
#477465000000
1!
1%
#477470000000
0!
0%
#477475000000
1!
1%
#477480000000
0!
0%
#477485000000
1!
1%
#477490000000
0!
0%
#477495000000
1!
1%
#477500000000
0!
0%
#477505000000
1!
1%
#477510000000
0!
0%
#477515000000
1!
1%
#477520000000
0!
0%
#477525000000
1!
1%
#477530000000
0!
0%
#477535000000
1!
1%
#477540000000
0!
0%
#477545000000
1!
1%
#477550000000
0!
0%
#477555000000
1!
1%
#477560000000
0!
0%
#477565000000
1!
1%
#477570000000
0!
0%
#477575000000
1!
1%
#477580000000
0!
0%
#477585000000
1!
1%
#477590000000
0!
0%
#477595000000
1!
1%
#477600000000
0!
0%
#477605000000
1!
1%
#477610000000
0!
0%
#477615000000
1!
1%
#477620000000
0!
0%
#477625000000
1!
1%
#477630000000
0!
0%
#477635000000
1!
1%
#477640000000
0!
0%
#477645000000
1!
1%
#477650000000
0!
0%
#477655000000
1!
1%
#477660000000
0!
0%
#477665000000
1!
1%
#477670000000
0!
0%
#477675000000
1!
1%
#477680000000
0!
0%
#477685000000
1!
1%
#477690000000
0!
0%
#477695000000
1!
1%
#477700000000
0!
0%
#477705000000
1!
1%
#477710000000
0!
0%
#477715000000
1!
1%
#477720000000
0!
0%
#477725000000
1!
1%
#477730000000
0!
0%
#477735000000
1!
1%
#477740000000
0!
0%
#477745000000
1!
1%
#477750000000
0!
0%
#477755000000
1!
1%
#477760000000
0!
0%
#477765000000
1!
1%
#477770000000
0!
0%
#477775000000
1!
1%
#477780000000
0!
0%
#477785000000
1!
1%
#477790000000
0!
0%
#477795000000
1!
1%
#477800000000
0!
0%
#477805000000
1!
1%
#477810000000
0!
0%
#477815000000
1!
1%
#477820000000
0!
0%
#477825000000
1!
1%
#477830000000
0!
0%
#477835000000
1!
1%
#477840000000
0!
0%
#477845000000
1!
1%
#477850000000
0!
0%
#477855000000
1!
1%
#477860000000
0!
0%
#477865000000
1!
1%
#477870000000
0!
0%
#477875000000
1!
1%
#477880000000
0!
0%
#477885000000
1!
1%
#477890000000
0!
0%
#477895000000
1!
1%
#477900000000
0!
0%
#477905000000
1!
1%
#477910000000
0!
0%
#477915000000
1!
1%
#477920000000
0!
0%
#477925000000
1!
1%
#477930000000
0!
0%
#477935000000
1!
1%
#477940000000
0!
0%
#477945000000
1!
1%
#477950000000
0!
0%
#477955000000
1!
1%
#477960000000
0!
0%
#477965000000
1!
1%
#477970000000
0!
0%
#477975000000
1!
1%
#477980000000
0!
0%
#477985000000
1!
1%
#477990000000
0!
0%
#477995000000
1!
1%
#478000000000
0!
0%
#478005000000
1!
1%
#478010000000
0!
0%
#478015000000
1!
1%
#478020000000
0!
0%
#478025000000
1!
1%
#478030000000
0!
0%
#478035000000
1!
1%
#478040000000
0!
0%
#478045000000
1!
1%
#478050000000
0!
0%
#478055000000
1!
1%
#478060000000
0!
0%
#478065000000
1!
1%
#478070000000
0!
0%
#478075000000
1!
1%
#478080000000
0!
0%
#478085000000
1!
1%
#478090000000
0!
0%
#478095000000
1!
1%
#478100000000
0!
0%
#478105000000
1!
1%
#478110000000
0!
0%
#478115000000
1!
1%
#478120000000
0!
0%
#478125000000
1!
1%
#478130000000
0!
0%
#478135000000
1!
1%
#478140000000
0!
0%
#478145000000
1!
1%
#478150000000
0!
0%
#478155000000
1!
1%
#478160000000
0!
0%
#478165000000
1!
1%
#478170000000
0!
0%
#478175000000
1!
1%
#478180000000
0!
0%
#478185000000
1!
1%
#478190000000
0!
0%
#478195000000
1!
1%
#478200000000
0!
0%
#478205000000
1!
1%
#478210000000
0!
0%
#478215000000
1!
1%
#478220000000
0!
0%
#478225000000
1!
1%
#478230000000
0!
0%
#478235000000
1!
1%
#478240000000
0!
0%
#478245000000
1!
1%
#478250000000
0!
0%
#478255000000
1!
1%
#478260000000
0!
0%
#478265000000
1!
1%
#478270000000
0!
0%
#478275000000
1!
1%
#478280000000
0!
0%
#478285000000
1!
1%
#478290000000
0!
0%
#478295000000
1!
1%
#478300000000
0!
0%
#478305000000
1!
1%
#478310000000
0!
0%
#478315000000
1!
1%
#478320000000
0!
0%
#478325000000
1!
1%
#478330000000
0!
0%
#478335000000
1!
1%
#478340000000
0!
0%
#478345000000
1!
1%
#478350000000
0!
0%
#478355000000
1!
1%
#478360000000
0!
0%
#478365000000
1!
1%
#478370000000
0!
0%
#478375000000
1!
1%
#478380000000
0!
0%
#478385000000
1!
1%
#478390000000
0!
0%
#478395000000
1!
1%
#478400000000
0!
0%
#478405000000
1!
1%
#478410000000
0!
0%
#478415000000
1!
1%
#478420000000
0!
0%
#478425000000
1!
1%
#478430000000
0!
0%
#478435000000
1!
1%
#478440000000
0!
0%
#478445000000
1!
1%
#478450000000
0!
0%
#478455000000
1!
1%
#478460000000
0!
0%
#478465000000
1!
1%
#478470000000
0!
0%
#478475000000
1!
1%
#478480000000
0!
0%
#478485000000
1!
1%
#478490000000
0!
0%
#478495000000
1!
1%
#478500000000
0!
0%
#478505000000
1!
1%
#478510000000
0!
0%
#478515000000
1!
1%
#478520000000
0!
0%
#478525000000
1!
1%
#478530000000
0!
0%
#478535000000
1!
1%
#478540000000
0!
0%
#478545000000
1!
1%
#478550000000
0!
0%
#478555000000
1!
1%
#478560000000
0!
0%
#478565000000
1!
1%
#478570000000
0!
0%
#478575000000
1!
1%
#478580000000
0!
0%
#478585000000
1!
1%
#478590000000
0!
0%
#478595000000
1!
1%
#478600000000
0!
0%
#478605000000
1!
1%
#478610000000
0!
0%
#478615000000
1!
1%
#478620000000
0!
0%
#478625000000
1!
1%
#478630000000
0!
0%
#478635000000
1!
1%
#478640000000
0!
0%
#478645000000
1!
1%
#478650000000
0!
0%
#478655000000
1!
1%
#478660000000
0!
0%
#478665000000
1!
1%
#478670000000
0!
0%
#478675000000
1!
1%
#478680000000
0!
0%
#478685000000
1!
1%
#478690000000
0!
0%
#478695000000
1!
1%
#478700000000
0!
0%
#478705000000
1!
1%
#478710000000
0!
0%
#478715000000
1!
1%
#478720000000
0!
0%
#478725000000
1!
1%
#478730000000
0!
0%
#478735000000
1!
1%
#478740000000
0!
0%
#478745000000
1!
1%
#478750000000
0!
0%
#478755000000
1!
1%
#478760000000
0!
0%
#478765000000
1!
1%
#478770000000
0!
0%
#478775000000
1!
1%
#478780000000
0!
0%
#478785000000
1!
1%
#478790000000
0!
0%
#478795000000
1!
1%
#478800000000
0!
0%
#478805000000
1!
1%
#478810000000
0!
0%
#478815000000
1!
1%
#478820000000
0!
0%
#478825000000
1!
1%
#478830000000
0!
0%
#478835000000
1!
1%
#478840000000
0!
0%
#478845000000
1!
1%
#478850000000
0!
0%
#478855000000
1!
1%
#478860000000
0!
0%
#478865000000
1!
1%
#478870000000
0!
0%
#478875000000
1!
1%
#478880000000
0!
0%
#478885000000
1!
1%
#478890000000
0!
0%
#478895000000
1!
1%
#478900000000
0!
0%
#478905000000
1!
1%
#478910000000
0!
0%
#478915000000
1!
1%
#478920000000
0!
0%
#478925000000
1!
1%
#478930000000
0!
0%
#478935000000
1!
1%
#478940000000
0!
0%
#478945000000
1!
1%
#478950000000
0!
0%
#478955000000
1!
1%
#478960000000
0!
0%
#478965000000
1!
1%
#478970000000
0!
0%
#478975000000
1!
1%
#478980000000
0!
0%
#478985000000
1!
1%
#478990000000
0!
0%
#478995000000
1!
1%
#479000000000
0!
0%
#479005000000
1!
1%
#479010000000
0!
0%
#479015000000
1!
1%
#479020000000
0!
0%
#479025000000
1!
1%
#479030000000
0!
0%
#479035000000
1!
1%
#479040000000
0!
0%
#479045000000
1!
1%
#479050000000
0!
0%
#479055000000
1!
1%
#479060000000
0!
0%
#479065000000
1!
1%
#479070000000
0!
0%
#479075000000
1!
1%
#479080000000
0!
0%
#479085000000
1!
1%
#479090000000
0!
0%
#479095000000
1!
1%
#479100000000
0!
0%
#479105000000
1!
1%
#479110000000
0!
0%
#479115000000
1!
1%
#479120000000
0!
0%
#479125000000
1!
1%
#479130000000
0!
0%
#479135000000
1!
1%
#479140000000
0!
0%
#479145000000
1!
1%
#479150000000
0!
0%
#479155000000
1!
1%
#479160000000
0!
0%
#479165000000
1!
1%
#479170000000
0!
0%
#479175000000
1!
1%
#479180000000
0!
0%
#479185000000
1!
1%
#479190000000
0!
0%
#479195000000
1!
1%
#479200000000
0!
0%
#479205000000
1!
1%
#479210000000
0!
0%
#479215000000
1!
1%
#479220000000
0!
0%
#479225000000
1!
1%
#479230000000
0!
0%
#479235000000
1!
1%
#479240000000
0!
0%
#479245000000
1!
1%
#479250000000
0!
0%
#479255000000
1!
1%
#479260000000
0!
0%
#479265000000
1!
1%
#479270000000
0!
0%
#479275000000
1!
1%
#479280000000
0!
0%
#479285000000
1!
1%
#479290000000
0!
0%
#479295000000
1!
1%
#479300000000
0!
0%
#479305000000
1!
1%
#479310000000
0!
0%
#479315000000
1!
1%
#479320000000
0!
0%
#479325000000
1!
1%
#479330000000
0!
0%
#479335000000
1!
1%
#479340000000
0!
0%
#479345000000
1!
1%
#479350000000
0!
0%
#479355000000
1!
1%
#479360000000
0!
0%
#479365000000
1!
1%
#479370000000
0!
0%
#479375000000
1!
1%
#479380000000
0!
0%
#479385000000
1!
1%
#479390000000
0!
0%
#479395000000
1!
1%
#479400000000
0!
0%
#479405000000
1!
1%
#479410000000
0!
0%
#479415000000
1!
1%
#479420000000
0!
0%
#479425000000
1!
1%
#479430000000
0!
0%
#479435000000
1!
1%
#479440000000
0!
0%
#479445000000
1!
1%
#479450000000
0!
0%
#479455000000
1!
1%
#479460000000
0!
0%
#479465000000
1!
1%
#479470000000
0!
0%
#479475000000
1!
1%
#479480000000
0!
0%
#479485000000
1!
1%
#479490000000
0!
0%
#479495000000
1!
1%
#479500000000
0!
0%
#479505000000
1!
1%
#479510000000
0!
0%
#479515000000
1!
1%
#479520000000
0!
0%
#479525000000
1!
1%
#479530000000
0!
0%
#479535000000
1!
1%
#479540000000
0!
0%
#479545000000
1!
1%
#479550000000
0!
0%
#479555000000
1!
1%
#479560000000
0!
0%
#479565000000
1!
1%
#479570000000
0!
0%
#479575000000
1!
1%
#479580000000
0!
0%
#479585000000
1!
1%
#479590000000
0!
0%
#479595000000
1!
1%
#479600000000
0!
0%
#479605000000
1!
1%
#479610000000
0!
0%
#479615000000
1!
1%
#479620000000
0!
0%
#479625000000
1!
1%
#479630000000
0!
0%
#479635000000
1!
1%
#479640000000
0!
0%
#479645000000
1!
1%
#479650000000
0!
0%
#479655000000
1!
1%
#479660000000
0!
0%
#479665000000
1!
1%
#479670000000
0!
0%
#479675000000
1!
1%
#479680000000
0!
0%
#479685000000
1!
1%
#479690000000
0!
0%
#479695000000
1!
1%
#479700000000
0!
0%
#479705000000
1!
1%
#479710000000
0!
0%
#479715000000
1!
1%
#479720000000
0!
0%
#479725000000
1!
1%
#479730000000
0!
0%
#479735000000
1!
1%
#479740000000
0!
0%
#479745000000
1!
1%
#479750000000
0!
0%
#479755000000
1!
1%
#479760000000
0!
0%
#479765000000
1!
1%
#479770000000
0!
0%
#479775000000
1!
1%
#479780000000
0!
0%
#479785000000
1!
1%
#479790000000
0!
0%
#479795000000
1!
1%
#479800000000
0!
0%
#479805000000
1!
1%
#479810000000
0!
0%
#479815000000
1!
1%
#479820000000
0!
0%
#479825000000
1!
1%
#479830000000
0!
0%
#479835000000
1!
1%
#479840000000
0!
0%
#479845000000
1!
1%
#479850000000
0!
0%
#479855000000
1!
1%
#479860000000
0!
0%
#479865000000
1!
1%
#479870000000
0!
0%
#479875000000
1!
1%
#479880000000
0!
0%
#479885000000
1!
1%
#479890000000
0!
0%
#479895000000
1!
1%
#479900000000
0!
0%
#479905000000
1!
1%
#479910000000
0!
0%
#479915000000
1!
1%
#479920000000
0!
0%
#479925000000
1!
1%
#479930000000
0!
0%
#479935000000
1!
1%
#479940000000
0!
0%
#479945000000
1!
1%
#479950000000
0!
0%
#479955000000
1!
1%
#479960000000
0!
0%
#479965000000
1!
1%
#479970000000
0!
0%
#479975000000
1!
1%
#479980000000
0!
0%
#479985000000
1!
1%
#479990000000
0!
0%
#479995000000
1!
1%
#480000000000
0!
0%
#480005000000
1!
1%
#480010000000
0!
0%
#480015000000
1!
1%
#480020000000
0!
0%
#480025000000
1!
1%
#480030000000
0!
0%
#480035000000
1!
1%
#480040000000
0!
0%
#480045000000
1!
1%
#480050000000
0!
0%
#480055000000
1!
1%
#480060000000
0!
0%
#480065000000
1!
1%
#480070000000
0!
0%
#480075000000
1!
1%
#480080000000
0!
0%
#480085000000
1!
1%
#480090000000
0!
0%
#480095000000
1!
1%
#480100000000
0!
0%
#480105000000
1!
1%
#480110000000
0!
0%
#480115000000
1!
1%
#480120000000
0!
0%
#480125000000
1!
1%
#480130000000
0!
0%
#480135000000
1!
1%
#480140000000
0!
0%
#480145000000
1!
1%
#480150000000
0!
0%
#480155000000
1!
1%
#480160000000
0!
0%
#480165000000
1!
1%
#480170000000
0!
0%
#480175000000
1!
1%
#480180000000
0!
0%
#480185000000
1!
1%
#480190000000
0!
0%
#480195000000
1!
1%
#480200000000
0!
0%
#480205000000
1!
1%
#480210000000
0!
0%
#480215000000
1!
1%
#480220000000
0!
0%
#480225000000
1!
1%
#480230000000
0!
0%
#480235000000
1!
1%
#480240000000
0!
0%
#480245000000
1!
1%
#480250000000
0!
0%
#480255000000
1!
1%
#480260000000
0!
0%
#480265000000
1!
1%
#480270000000
0!
0%
#480275000000
1!
1%
#480280000000
0!
0%
#480285000000
1!
1%
#480290000000
0!
0%
#480295000000
1!
1%
#480300000000
0!
0%
#480305000000
1!
1%
#480310000000
0!
0%
#480315000000
1!
1%
#480320000000
0!
0%
#480325000000
1!
1%
#480330000000
0!
0%
#480335000000
1!
1%
#480340000000
0!
0%
#480345000000
1!
1%
#480350000000
0!
0%
#480355000000
1!
1%
#480360000000
0!
0%
#480365000000
1!
1%
#480370000000
0!
0%
#480375000000
1!
1%
#480380000000
0!
0%
#480385000000
1!
1%
#480390000000
0!
0%
#480395000000
1!
1%
#480400000000
0!
0%
#480405000000
1!
1%
#480410000000
0!
0%
#480415000000
1!
1%
#480420000000
0!
0%
#480425000000
1!
1%
#480430000000
0!
0%
#480435000000
1!
1%
#480440000000
0!
0%
#480445000000
1!
1%
#480450000000
0!
0%
#480455000000
1!
1%
#480460000000
0!
0%
#480465000000
1!
1%
#480470000000
0!
0%
#480475000000
1!
1%
#480480000000
0!
0%
#480485000000
1!
1%
#480490000000
0!
0%
#480495000000
1!
1%
#480500000000
0!
0%
#480505000000
1!
1%
#480510000000
0!
0%
#480515000000
1!
1%
#480520000000
0!
0%
#480525000000
1!
1%
#480530000000
0!
0%
#480535000000
1!
1%
#480540000000
0!
0%
#480545000000
1!
1%
#480550000000
0!
0%
#480555000000
1!
1%
#480560000000
0!
0%
#480565000000
1!
1%
#480570000000
0!
0%
#480575000000
1!
1%
#480580000000
0!
0%
#480585000000
1!
1%
#480590000000
0!
0%
#480595000000
1!
1%
#480600000000
0!
0%
#480605000000
1!
1%
#480610000000
0!
0%
#480615000000
1!
1%
#480620000000
0!
0%
#480625000000
1!
1%
#480630000000
0!
0%
#480635000000
1!
1%
#480640000000
0!
0%
#480645000000
1!
1%
#480650000000
0!
0%
#480655000000
1!
1%
#480660000000
0!
0%
#480665000000
1!
1%
#480670000000
0!
0%
#480675000000
1!
1%
#480680000000
0!
0%
#480685000000
1!
1%
#480690000000
0!
0%
#480695000000
1!
1%
#480700000000
0!
0%
#480705000000
1!
1%
#480710000000
0!
0%
#480715000000
1!
1%
#480720000000
0!
0%
#480725000000
1!
1%
#480730000000
0!
0%
#480735000000
1!
1%
#480740000000
0!
0%
#480745000000
1!
1%
#480750000000
0!
0%
#480755000000
1!
1%
#480760000000
0!
0%
#480765000000
1!
1%
#480770000000
0!
0%
#480775000000
1!
1%
#480780000000
0!
0%
#480785000000
1!
1%
#480790000000
0!
0%
#480795000000
1!
1%
#480800000000
0!
0%
#480805000000
1!
1%
#480810000000
0!
0%
#480815000000
1!
1%
#480820000000
0!
0%
#480825000000
1!
1%
#480830000000
0!
0%
#480835000000
1!
1%
#480840000000
0!
0%
#480845000000
1!
1%
#480850000000
0!
0%
#480855000000
1!
1%
#480860000000
0!
0%
#480865000000
1!
1%
#480870000000
0!
0%
#480875000000
1!
1%
#480880000000
0!
0%
#480885000000
1!
1%
#480890000000
0!
0%
#480895000000
1!
1%
#480900000000
0!
0%
#480905000000
1!
1%
#480910000000
0!
0%
#480915000000
1!
1%
#480920000000
0!
0%
#480925000000
1!
1%
#480930000000
0!
0%
#480935000000
1!
1%
#480940000000
0!
0%
#480945000000
1!
1%
#480950000000
0!
0%
#480955000000
1!
1%
#480960000000
0!
0%
#480965000000
1!
1%
#480970000000
0!
0%
#480975000000
1!
1%
#480980000000
0!
0%
#480985000000
1!
1%
#480990000000
0!
0%
#480995000000
1!
1%
#481000000000
0!
0%
#481005000000
1!
1%
#481010000000
0!
0%
#481015000000
1!
1%
#481020000000
0!
0%
#481025000000
1!
1%
#481030000000
0!
0%
#481035000000
1!
1%
#481040000000
0!
0%
#481045000000
1!
1%
#481050000000
0!
0%
#481055000000
1!
1%
#481060000000
0!
0%
#481065000000
1!
1%
#481070000000
0!
0%
#481075000000
1!
1%
#481080000000
0!
0%
#481085000000
1!
1%
#481090000000
0!
0%
#481095000000
1!
1%
#481100000000
0!
0%
#481105000000
1!
1%
#481110000000
0!
0%
#481115000000
1!
1%
#481120000000
0!
0%
#481125000000
1!
1%
#481130000000
0!
0%
#481135000000
1!
1%
#481140000000
0!
0%
#481145000000
1!
1%
#481150000000
0!
0%
#481155000000
1!
1%
#481160000000
0!
0%
#481165000000
1!
1%
#481170000000
0!
0%
#481175000000
1!
1%
#481180000000
0!
0%
#481185000000
1!
1%
#481190000000
0!
0%
#481195000000
1!
1%
#481200000000
0!
0%
#481205000000
1!
1%
#481210000000
0!
0%
#481215000000
1!
1%
#481220000000
0!
0%
#481225000000
1!
1%
#481230000000
0!
0%
#481235000000
1!
1%
#481240000000
0!
0%
#481245000000
1!
1%
#481250000000
0!
0%
#481255000000
1!
1%
#481260000000
0!
0%
#481265000000
1!
1%
#481270000000
0!
0%
#481275000000
1!
1%
#481280000000
0!
0%
#481285000000
1!
1%
#481290000000
0!
0%
#481295000000
1!
1%
#481300000000
0!
0%
#481305000000
1!
1%
#481310000000
0!
0%
#481315000000
1!
1%
#481320000000
0!
0%
#481325000000
1!
1%
#481330000000
0!
0%
#481335000000
1!
1%
#481340000000
0!
0%
#481345000000
1!
1%
#481350000000
0!
0%
#481355000000
1!
1%
#481360000000
0!
0%
#481365000000
1!
1%
#481370000000
0!
0%
#481375000000
1!
1%
#481380000000
0!
0%
#481385000000
1!
1%
#481390000000
0!
0%
#481395000000
1!
1%
#481400000000
0!
0%
#481405000000
1!
1%
#481410000000
0!
0%
#481415000000
1!
1%
#481420000000
0!
0%
#481425000000
1!
1%
#481430000000
0!
0%
#481435000000
1!
1%
#481440000000
0!
0%
#481445000000
1!
1%
#481450000000
0!
0%
#481455000000
1!
1%
#481460000000
0!
0%
#481465000000
1!
1%
#481470000000
0!
0%
#481475000000
1!
1%
#481480000000
0!
0%
#481485000000
1!
1%
#481490000000
0!
0%
#481495000000
1!
1%
#481500000000
0!
0%
#481505000000
1!
1%
#481510000000
0!
0%
#481515000000
1!
1%
#481520000000
0!
0%
#481525000000
1!
1%
#481530000000
0!
0%
#481535000000
1!
1%
#481540000000
0!
0%
#481545000000
1!
1%
#481550000000
0!
0%
#481555000000
1!
1%
#481560000000
0!
0%
#481565000000
1!
1%
#481570000000
0!
0%
#481575000000
1!
1%
#481580000000
0!
0%
#481585000000
1!
1%
#481590000000
0!
0%
#481595000000
1!
1%
#481600000000
0!
0%
#481605000000
1!
1%
#481610000000
0!
0%
#481615000000
1!
1%
#481620000000
0!
0%
#481625000000
1!
1%
#481630000000
0!
0%
#481635000000
1!
1%
#481640000000
0!
0%
#481645000000
1!
1%
#481650000000
0!
0%
#481655000000
1!
1%
#481660000000
0!
0%
#481665000000
1!
1%
#481670000000
0!
0%
#481675000000
1!
1%
#481680000000
0!
0%
#481685000000
1!
1%
#481690000000
0!
0%
#481695000000
1!
1%
#481700000000
0!
0%
#481705000000
1!
1%
#481710000000
0!
0%
#481715000000
1!
1%
#481720000000
0!
0%
#481725000000
1!
1%
#481730000000
0!
0%
#481735000000
1!
1%
#481740000000
0!
0%
#481745000000
1!
1%
#481750000000
0!
0%
#481755000000
1!
1%
#481760000000
0!
0%
#481765000000
1!
1%
#481770000000
0!
0%
#481775000000
1!
1%
#481780000000
0!
0%
#481785000000
1!
1%
#481790000000
0!
0%
#481795000000
1!
1%
#481800000000
0!
0%
#481805000000
1!
1%
#481810000000
0!
0%
#481815000000
1!
1%
#481820000000
0!
0%
#481825000000
1!
1%
#481830000000
0!
0%
#481835000000
1!
1%
#481840000000
0!
0%
#481845000000
1!
1%
#481850000000
0!
0%
#481855000000
1!
1%
#481860000000
0!
0%
#481865000000
1!
1%
#481870000000
0!
0%
#481875000000
1!
1%
#481880000000
0!
0%
#481885000000
1!
1%
#481890000000
0!
0%
#481895000000
1!
1%
#481900000000
0!
0%
#481905000000
1!
1%
#481910000000
0!
0%
#481915000000
1!
1%
#481920000000
0!
0%
#481925000000
1!
1%
#481930000000
0!
0%
#481935000000
1!
1%
#481940000000
0!
0%
#481945000000
1!
1%
#481950000000
0!
0%
#481955000000
1!
1%
#481960000000
0!
0%
#481965000000
1!
1%
#481970000000
0!
0%
#481975000000
1!
1%
#481980000000
0!
0%
#481985000000
1!
1%
#481990000000
0!
0%
#481995000000
1!
1%
#482000000000
0!
0%
#482005000000
1!
1%
#482010000000
0!
0%
#482015000000
1!
1%
#482020000000
0!
0%
#482025000000
1!
1%
#482030000000
0!
0%
#482035000000
1!
1%
#482040000000
0!
0%
#482045000000
1!
1%
#482050000000
0!
0%
#482055000000
1!
1%
#482060000000
0!
0%
#482065000000
1!
1%
#482070000000
0!
0%
#482075000000
1!
1%
#482080000000
0!
0%
#482085000000
1!
1%
#482090000000
0!
0%
#482095000000
1!
1%
#482100000000
0!
0%
#482105000000
1!
1%
#482110000000
0!
0%
#482115000000
1!
1%
#482120000000
0!
0%
#482125000000
1!
1%
#482130000000
0!
0%
#482135000000
1!
1%
#482140000000
0!
0%
#482145000000
1!
1%
#482150000000
0!
0%
#482155000000
1!
1%
#482160000000
0!
0%
#482165000000
1!
1%
#482170000000
0!
0%
#482175000000
1!
1%
#482180000000
0!
0%
#482185000000
1!
1%
#482190000000
0!
0%
#482195000000
1!
1%
#482200000000
0!
0%
#482205000000
1!
1%
#482210000000
0!
0%
#482215000000
1!
1%
#482220000000
0!
0%
#482225000000
1!
1%
#482230000000
0!
0%
#482235000000
1!
1%
#482240000000
0!
0%
#482245000000
1!
1%
#482250000000
0!
0%
#482255000000
1!
1%
#482260000000
0!
0%
#482265000000
1!
1%
#482270000000
0!
0%
#482275000000
1!
1%
#482280000000
0!
0%
#482285000000
1!
1%
#482290000000
0!
0%
#482295000000
1!
1%
#482300000000
0!
0%
#482305000000
1!
1%
#482310000000
0!
0%
#482315000000
1!
1%
#482320000000
0!
0%
#482325000000
1!
1%
#482330000000
0!
0%
#482335000000
1!
1%
#482340000000
0!
0%
#482345000000
1!
1%
#482350000000
0!
0%
#482355000000
1!
1%
#482360000000
0!
0%
#482365000000
1!
1%
#482370000000
0!
0%
#482375000000
1!
1%
#482380000000
0!
0%
#482385000000
1!
1%
#482390000000
0!
0%
#482395000000
1!
1%
#482400000000
0!
0%
#482405000000
1!
1%
#482410000000
0!
0%
#482415000000
1!
1%
#482420000000
0!
0%
#482425000000
1!
1%
#482430000000
0!
0%
#482435000000
1!
1%
#482440000000
0!
0%
#482445000000
1!
1%
#482450000000
0!
0%
#482455000000
1!
1%
#482460000000
0!
0%
#482465000000
1!
1%
#482470000000
0!
0%
#482475000000
1!
1%
#482480000000
0!
0%
#482485000000
1!
1%
#482490000000
0!
0%
#482495000000
1!
1%
#482500000000
0!
0%
#482505000000
1!
1%
#482510000000
0!
0%
#482515000000
1!
1%
#482520000000
0!
0%
#482525000000
1!
1%
#482530000000
0!
0%
#482535000000
1!
1%
#482540000000
0!
0%
#482545000000
1!
1%
#482550000000
0!
0%
#482555000000
1!
1%
#482560000000
0!
0%
#482565000000
1!
1%
#482570000000
0!
0%
#482575000000
1!
1%
#482580000000
0!
0%
#482585000000
1!
1%
#482590000000
0!
0%
#482595000000
1!
1%
#482600000000
0!
0%
#482605000000
1!
1%
#482610000000
0!
0%
#482615000000
1!
1%
#482620000000
0!
0%
#482625000000
1!
1%
#482630000000
0!
0%
#482635000000
1!
1%
#482640000000
0!
0%
#482645000000
1!
1%
#482650000000
0!
0%
#482655000000
1!
1%
#482660000000
0!
0%
#482665000000
1!
1%
#482670000000
0!
0%
#482675000000
1!
1%
#482680000000
0!
0%
#482685000000
1!
1%
#482690000000
0!
0%
#482695000000
1!
1%
#482700000000
0!
0%
#482705000000
1!
1%
#482710000000
0!
0%
#482715000000
1!
1%
#482720000000
0!
0%
#482725000000
1!
1%
#482730000000
0!
0%
#482735000000
1!
1%
#482740000000
0!
0%
#482745000000
1!
1%
#482750000000
0!
0%
#482755000000
1!
1%
#482760000000
0!
0%
#482765000000
1!
1%
#482770000000
0!
0%
#482775000000
1!
1%
#482780000000
0!
0%
#482785000000
1!
1%
#482790000000
0!
0%
#482795000000
1!
1%
#482800000000
0!
0%
#482805000000
1!
1%
#482810000000
0!
0%
#482815000000
1!
1%
#482820000000
0!
0%
#482825000000
1!
1%
#482830000000
0!
0%
#482835000000
1!
1%
#482840000000
0!
0%
#482845000000
1!
1%
#482850000000
0!
0%
#482855000000
1!
1%
#482860000000
0!
0%
#482865000000
1!
1%
#482870000000
0!
0%
#482875000000
1!
1%
#482880000000
0!
0%
#482885000000
1!
1%
#482890000000
0!
0%
#482895000000
1!
1%
#482900000000
0!
0%
#482905000000
1!
1%
#482910000000
0!
0%
#482915000000
1!
1%
#482920000000
0!
0%
#482925000000
1!
1%
#482930000000
0!
0%
#482935000000
1!
1%
#482940000000
0!
0%
#482945000000
1!
1%
#482950000000
0!
0%
#482955000000
1!
1%
#482960000000
0!
0%
#482965000000
1!
1%
#482970000000
0!
0%
#482975000000
1!
1%
#482980000000
0!
0%
#482985000000
1!
1%
#482990000000
0!
0%
#482995000000
1!
1%
#483000000000
0!
0%
#483005000000
1!
1%
#483010000000
0!
0%
#483015000000
1!
1%
#483020000000
0!
0%
#483025000000
1!
1%
#483030000000
0!
0%
#483035000000
1!
1%
#483040000000
0!
0%
#483045000000
1!
1%
#483050000000
0!
0%
#483055000000
1!
1%
#483060000000
0!
0%
#483065000000
1!
1%
#483070000000
0!
0%
#483075000000
1!
1%
#483080000000
0!
0%
#483085000000
1!
1%
#483090000000
0!
0%
#483095000000
1!
1%
#483100000000
0!
0%
#483105000000
1!
1%
#483110000000
0!
0%
#483115000000
1!
1%
#483120000000
0!
0%
#483125000000
1!
1%
#483130000000
0!
0%
#483135000000
1!
1%
#483140000000
0!
0%
#483145000000
1!
1%
#483150000000
0!
0%
#483155000000
1!
1%
#483160000000
0!
0%
#483165000000
1!
1%
#483170000000
0!
0%
#483175000000
1!
1%
#483180000000
0!
0%
#483185000000
1!
1%
#483190000000
0!
0%
#483195000000
1!
1%
#483200000000
0!
0%
#483205000000
1!
1%
#483210000000
0!
0%
#483215000000
1!
1%
#483220000000
0!
0%
#483225000000
1!
1%
#483230000000
0!
0%
#483235000000
1!
1%
#483240000000
0!
0%
#483245000000
1!
1%
#483250000000
0!
0%
#483255000000
1!
1%
#483260000000
0!
0%
#483265000000
1!
1%
#483270000000
0!
0%
#483275000000
1!
1%
#483280000000
0!
0%
#483285000000
1!
1%
#483290000000
0!
0%
#483295000000
1!
1%
#483300000000
0!
0%
#483305000000
1!
1%
#483310000000
0!
0%
#483315000000
1!
1%
#483320000000
0!
0%
#483325000000
1!
1%
#483330000000
0!
0%
#483335000000
1!
1%
#483340000000
0!
0%
#483345000000
1!
1%
#483350000000
0!
0%
#483355000000
1!
1%
#483360000000
0!
0%
#483365000000
1!
1%
#483370000000
0!
0%
#483375000000
1!
1%
#483380000000
0!
0%
#483385000000
1!
1%
#483390000000
0!
0%
#483395000000
1!
1%
#483400000000
0!
0%
#483405000000
1!
1%
#483410000000
0!
0%
#483415000000
1!
1%
#483420000000
0!
0%
#483425000000
1!
1%
#483430000000
0!
0%
#483435000000
1!
1%
#483440000000
0!
0%
#483445000000
1!
1%
#483450000000
0!
0%
#483455000000
1!
1%
#483460000000
0!
0%
#483465000000
1!
1%
#483470000000
0!
0%
#483475000000
1!
1%
#483480000000
0!
0%
#483485000000
1!
1%
#483490000000
0!
0%
#483495000000
1!
1%
#483500000000
0!
0%
#483505000000
1!
1%
#483510000000
0!
0%
#483515000000
1!
1%
#483520000000
0!
0%
#483525000000
1!
1%
#483530000000
0!
0%
#483535000000
1!
1%
#483540000000
0!
0%
#483545000000
1!
1%
#483550000000
0!
0%
#483555000000
1!
1%
#483560000000
0!
0%
#483565000000
1!
1%
#483570000000
0!
0%
#483575000000
1!
1%
#483580000000
0!
0%
#483585000000
1!
1%
#483590000000
0!
0%
#483595000000
1!
1%
#483600000000
0!
0%
#483605000000
1!
1%
#483610000000
0!
0%
#483615000000
1!
1%
#483620000000
0!
0%
#483625000000
1!
1%
#483630000000
0!
0%
#483635000000
1!
1%
#483640000000
0!
0%
#483645000000
1!
1%
#483650000000
0!
0%
#483655000000
1!
1%
#483660000000
0!
0%
#483665000000
1!
1%
#483670000000
0!
0%
#483675000000
1!
1%
#483680000000
0!
0%
#483685000000
1!
1%
#483690000000
0!
0%
#483695000000
1!
1%
#483700000000
0!
0%
#483705000000
1!
1%
#483710000000
0!
0%
#483715000000
1!
1%
#483720000000
0!
0%
#483725000000
1!
1%
#483730000000
0!
0%
#483735000000
1!
1%
#483740000000
0!
0%
#483745000000
1!
1%
#483750000000
0!
0%
#483755000000
1!
1%
#483760000000
0!
0%
#483765000000
1!
1%
#483770000000
0!
0%
#483775000000
1!
1%
#483780000000
0!
0%
#483785000000
1!
1%
#483790000000
0!
0%
#483795000000
1!
1%
#483800000000
0!
0%
#483805000000
1!
1%
#483810000000
0!
0%
#483815000000
1!
1%
#483820000000
0!
0%
#483825000000
1!
1%
#483830000000
0!
0%
#483835000000
1!
1%
#483840000000
0!
0%
#483845000000
1!
1%
#483850000000
0!
0%
#483855000000
1!
1%
#483860000000
0!
0%
#483865000000
1!
1%
#483870000000
0!
0%
#483875000000
1!
1%
#483880000000
0!
0%
#483885000000
1!
1%
#483890000000
0!
0%
#483895000000
1!
1%
#483900000000
0!
0%
#483905000000
1!
1%
#483910000000
0!
0%
#483915000000
1!
1%
#483920000000
0!
0%
#483925000000
1!
1%
#483930000000
0!
0%
#483935000000
1!
1%
#483940000000
0!
0%
#483945000000
1!
1%
#483950000000
0!
0%
#483955000000
1!
1%
#483960000000
0!
0%
#483965000000
1!
1%
#483970000000
0!
0%
#483975000000
1!
1%
#483980000000
0!
0%
#483985000000
1!
1%
#483990000000
0!
0%
#483995000000
1!
1%
#484000000000
0!
0%
#484005000000
1!
1%
#484010000000
0!
0%
#484015000000
1!
1%
#484020000000
0!
0%
#484025000000
1!
1%
#484030000000
0!
0%
#484035000000
1!
1%
#484040000000
0!
0%
#484045000000
1!
1%
#484050000000
0!
0%
#484055000000
1!
1%
#484060000000
0!
0%
#484065000000
1!
1%
#484070000000
0!
0%
#484075000000
1!
1%
#484080000000
0!
0%
#484085000000
1!
1%
#484090000000
0!
0%
#484095000000
1!
1%
#484100000000
0!
0%
#484105000000
1!
1%
#484110000000
0!
0%
#484115000000
1!
1%
#484120000000
0!
0%
#484125000000
1!
1%
#484130000000
0!
0%
#484135000000
1!
1%
#484140000000
0!
0%
#484145000000
1!
1%
#484150000000
0!
0%
#484155000000
1!
1%
#484160000000
0!
0%
#484165000000
1!
1%
#484170000000
0!
0%
#484175000000
1!
1%
#484180000000
0!
0%
#484185000000
1!
1%
#484190000000
0!
0%
#484195000000
1!
1%
#484200000000
0!
0%
#484205000000
1!
1%
#484210000000
0!
0%
#484215000000
1!
1%
#484220000000
0!
0%
#484225000000
1!
1%
#484230000000
0!
0%
#484235000000
1!
1%
#484240000000
0!
0%
#484245000000
1!
1%
#484250000000
0!
0%
#484255000000
1!
1%
#484260000000
0!
0%
#484265000000
1!
1%
#484270000000
0!
0%
#484275000000
1!
1%
#484280000000
0!
0%
#484285000000
1!
1%
#484290000000
0!
0%
#484295000000
1!
1%
#484300000000
0!
0%
#484305000000
1!
1%
#484310000000
0!
0%
#484315000000
1!
1%
#484320000000
0!
0%
#484325000000
1!
1%
#484330000000
0!
0%
#484335000000
1!
1%
#484340000000
0!
0%
#484345000000
1!
1%
#484350000000
0!
0%
#484355000000
1!
1%
#484360000000
0!
0%
#484365000000
1!
1%
#484370000000
0!
0%
#484375000000
1!
1%
#484380000000
0!
0%
#484385000000
1!
1%
#484390000000
0!
0%
#484395000000
1!
1%
#484400000000
0!
0%
#484405000000
1!
1%
#484410000000
0!
0%
#484415000000
1!
1%
#484420000000
0!
0%
#484425000000
1!
1%
#484430000000
0!
0%
#484435000000
1!
1%
#484440000000
0!
0%
#484445000000
1!
1%
#484450000000
0!
0%
#484455000000
1!
1%
#484460000000
0!
0%
#484465000000
1!
1%
#484470000000
0!
0%
#484475000000
1!
1%
#484480000000
0!
0%
#484485000000
1!
1%
#484490000000
0!
0%
#484495000000
1!
1%
#484500000000
0!
0%
#484505000000
1!
1%
#484510000000
0!
0%
#484515000000
1!
1%
#484520000000
0!
0%
#484525000000
1!
1%
#484530000000
0!
0%
#484535000000
1!
1%
#484540000000
0!
0%
#484545000000
1!
1%
#484550000000
0!
0%
#484555000000
1!
1%
#484560000000
0!
0%
#484565000000
1!
1%
#484570000000
0!
0%
#484575000000
1!
1%
#484580000000
0!
0%
#484585000000
1!
1%
#484590000000
0!
0%
#484595000000
1!
1%
#484600000000
0!
0%
#484605000000
1!
1%
#484610000000
0!
0%
#484615000000
1!
1%
#484620000000
0!
0%
#484625000000
1!
1%
#484630000000
0!
0%
#484635000000
1!
1%
#484640000000
0!
0%
#484645000000
1!
1%
#484650000000
0!
0%
#484655000000
1!
1%
#484660000000
0!
0%
#484665000000
1!
1%
#484670000000
0!
0%
#484675000000
1!
1%
#484680000000
0!
0%
#484685000000
1!
1%
#484690000000
0!
0%
#484695000000
1!
1%
#484700000000
0!
0%
#484705000000
1!
1%
#484710000000
0!
0%
#484715000000
1!
1%
#484720000000
0!
0%
#484725000000
1!
1%
#484730000000
0!
0%
#484735000000
1!
1%
#484740000000
0!
0%
#484745000000
1!
1%
#484750000000
0!
0%
#484755000000
1!
1%
#484760000000
0!
0%
#484765000000
1!
1%
#484770000000
0!
0%
#484775000000
1!
1%
#484780000000
0!
0%
#484785000000
1!
1%
#484790000000
0!
0%
#484795000000
1!
1%
#484800000000
0!
0%
#484805000000
1!
1%
#484810000000
0!
0%
#484815000000
1!
1%
#484820000000
0!
0%
#484825000000
1!
1%
#484830000000
0!
0%
#484835000000
1!
1%
#484840000000
0!
0%
#484845000000
1!
1%
#484850000000
0!
0%
#484855000000
1!
1%
#484860000000
0!
0%
#484865000000
1!
1%
#484870000000
0!
0%
#484875000000
1!
1%
#484880000000
0!
0%
#484885000000
1!
1%
#484890000000
0!
0%
#484895000000
1!
1%
#484900000000
0!
0%
#484905000000
1!
1%
#484910000000
0!
0%
#484915000000
1!
1%
#484920000000
0!
0%
#484925000000
1!
1%
#484930000000
0!
0%
#484935000000
1!
1%
#484940000000
0!
0%
#484945000000
1!
1%
#484950000000
0!
0%
#484955000000
1!
1%
#484960000000
0!
0%
#484965000000
1!
1%
#484970000000
0!
0%
#484975000000
1!
1%
#484980000000
0!
0%
#484985000000
1!
1%
#484990000000
0!
0%
#484995000000
1!
1%
#485000000000
0!
0%
#485005000000
1!
1%
#485010000000
0!
0%
#485015000000
1!
1%
#485020000000
0!
0%
#485025000000
1!
1%
#485030000000
0!
0%
#485035000000
1!
1%
#485040000000
0!
0%
#485045000000
1!
1%
#485050000000
0!
0%
#485055000000
1!
1%
#485060000000
0!
0%
#485065000000
1!
1%
#485070000000
0!
0%
#485075000000
1!
1%
#485080000000
0!
0%
#485085000000
1!
1%
#485090000000
0!
0%
#485095000000
1!
1%
#485100000000
0!
0%
#485105000000
1!
1%
#485110000000
0!
0%
#485115000000
1!
1%
#485120000000
0!
0%
#485125000000
1!
1%
#485130000000
0!
0%
#485135000000
1!
1%
#485140000000
0!
0%
#485145000000
1!
1%
#485150000000
0!
0%
#485155000000
1!
1%
#485160000000
0!
0%
#485165000000
1!
1%
#485170000000
0!
0%
#485175000000
1!
1%
#485180000000
0!
0%
#485185000000
1!
1%
#485190000000
0!
0%
#485195000000
1!
1%
#485200000000
0!
0%
#485205000000
1!
1%
#485210000000
0!
0%
#485215000000
1!
1%
#485220000000
0!
0%
#485225000000
1!
1%
#485230000000
0!
0%
#485235000000
1!
1%
#485240000000
0!
0%
#485245000000
1!
1%
#485250000000
0!
0%
#485255000000
1!
1%
#485260000000
0!
0%
#485265000000
1!
1%
#485270000000
0!
0%
#485275000000
1!
1%
#485280000000
0!
0%
#485285000000
1!
1%
#485290000000
0!
0%
#485295000000
1!
1%
#485300000000
0!
0%
#485305000000
1!
1%
#485310000000
0!
0%
#485315000000
1!
1%
#485320000000
0!
0%
#485325000000
1!
1%
#485330000000
0!
0%
#485335000000
1!
1%
#485340000000
0!
0%
#485345000000
1!
1%
#485350000000
0!
0%
#485355000000
1!
1%
#485360000000
0!
0%
#485365000000
1!
1%
#485370000000
0!
0%
#485375000000
1!
1%
#485380000000
0!
0%
#485385000000
1!
1%
#485390000000
0!
0%
#485395000000
1!
1%
#485400000000
0!
0%
#485405000000
1!
1%
#485410000000
0!
0%
#485415000000
1!
1%
#485420000000
0!
0%
#485425000000
1!
1%
#485430000000
0!
0%
#485435000000
1!
1%
#485440000000
0!
0%
#485445000000
1!
1%
#485450000000
0!
0%
#485455000000
1!
1%
#485460000000
0!
0%
#485465000000
1!
1%
#485470000000
0!
0%
#485475000000
1!
1%
#485480000000
0!
0%
#485485000000
1!
1%
#485490000000
0!
0%
#485495000000
1!
1%
#485500000000
0!
0%
#485505000000
1!
1%
#485510000000
0!
0%
#485515000000
1!
1%
#485520000000
0!
0%
#485525000000
1!
1%
#485530000000
0!
0%
#485535000000
1!
1%
#485540000000
0!
0%
#485545000000
1!
1%
#485550000000
0!
0%
#485555000000
1!
1%
#485560000000
0!
0%
#485565000000
1!
1%
#485570000000
0!
0%
#485575000000
1!
1%
#485580000000
0!
0%
#485585000000
1!
1%
#485590000000
0!
0%
#485595000000
1!
1%
#485600000000
0!
0%
#485605000000
1!
1%
#485610000000
0!
0%
#485615000000
1!
1%
#485620000000
0!
0%
#485625000000
1!
1%
#485630000000
0!
0%
#485635000000
1!
1%
#485640000000
0!
0%
#485645000000
1!
1%
#485650000000
0!
0%
#485655000000
1!
1%
#485660000000
0!
0%
#485665000000
1!
1%
#485670000000
0!
0%
#485675000000
1!
1%
#485680000000
0!
0%
#485685000000
1!
1%
#485690000000
0!
0%
#485695000000
1!
1%
#485700000000
0!
0%
#485705000000
1!
1%
#485710000000
0!
0%
#485715000000
1!
1%
#485720000000
0!
0%
#485725000000
1!
1%
#485730000000
0!
0%
#485735000000
1!
1%
#485740000000
0!
0%
#485745000000
1!
1%
#485750000000
0!
0%
#485755000000
1!
1%
#485760000000
0!
0%
#485765000000
1!
1%
#485770000000
0!
0%
#485775000000
1!
1%
#485780000000
0!
0%
#485785000000
1!
1%
#485790000000
0!
0%
#485795000000
1!
1%
#485800000000
0!
0%
#485805000000
1!
1%
#485810000000
0!
0%
#485815000000
1!
1%
#485820000000
0!
0%
#485825000000
1!
1%
#485830000000
0!
0%
#485835000000
1!
1%
#485840000000
0!
0%
#485845000000
1!
1%
#485850000000
0!
0%
#485855000000
1!
1%
#485860000000
0!
0%
#485865000000
1!
1%
#485870000000
0!
0%
#485875000000
1!
1%
#485880000000
0!
0%
#485885000000
1!
1%
#485890000000
0!
0%
#485895000000
1!
1%
#485900000000
0!
0%
#485905000000
1!
1%
#485910000000
0!
0%
#485915000000
1!
1%
#485920000000
0!
0%
#485925000000
1!
1%
#485930000000
0!
0%
#485935000000
1!
1%
#485940000000
0!
0%
#485945000000
1!
1%
#485950000000
0!
0%
#485955000000
1!
1%
#485960000000
0!
0%
#485965000000
1!
1%
#485970000000
0!
0%
#485975000000
1!
1%
#485980000000
0!
0%
#485985000000
1!
1%
#485990000000
0!
0%
#485995000000
1!
1%
#486000000000
0!
0%
#486005000000
1!
1%
#486010000000
0!
0%
#486015000000
1!
1%
#486020000000
0!
0%
#486025000000
1!
1%
#486030000000
0!
0%
#486035000000
1!
1%
#486040000000
0!
0%
#486045000000
1!
1%
#486050000000
0!
0%
#486055000000
1!
1%
#486060000000
0!
0%
#486065000000
1!
1%
#486070000000
0!
0%
#486075000000
1!
1%
#486080000000
0!
0%
#486085000000
1!
1%
#486090000000
0!
0%
#486095000000
1!
1%
#486100000000
0!
0%
#486105000000
1!
1%
#486110000000
0!
0%
#486115000000
1!
1%
#486120000000
0!
0%
#486125000000
1!
1%
#486130000000
0!
0%
#486135000000
1!
1%
#486140000000
0!
0%
#486145000000
1!
1%
#486150000000
0!
0%
#486155000000
1!
1%
#486160000000
0!
0%
#486165000000
1!
1%
#486170000000
0!
0%
#486175000000
1!
1%
#486180000000
0!
0%
#486185000000
1!
1%
#486190000000
0!
0%
#486195000000
1!
1%
#486200000000
0!
0%
#486205000000
1!
1%
#486210000000
0!
0%
#486215000000
1!
1%
#486220000000
0!
0%
#486225000000
1!
1%
#486230000000
0!
0%
#486235000000
1!
1%
#486240000000
0!
0%
#486245000000
1!
1%
#486250000000
0!
0%
#486255000000
1!
1%
#486260000000
0!
0%
#486265000000
1!
1%
#486270000000
0!
0%
#486275000000
1!
1%
#486280000000
0!
0%
#486285000000
1!
1%
#486290000000
0!
0%
#486295000000
1!
1%
#486300000000
0!
0%
#486305000000
1!
1%
#486310000000
0!
0%
#486315000000
1!
1%
#486320000000
0!
0%
#486325000000
1!
1%
#486330000000
0!
0%
#486335000000
1!
1%
#486340000000
0!
0%
#486345000000
1!
1%
#486350000000
0!
0%
#486355000000
1!
1%
#486360000000
0!
0%
#486365000000
1!
1%
#486370000000
0!
0%
#486375000000
1!
1%
#486380000000
0!
0%
#486385000000
1!
1%
#486390000000
0!
0%
#486395000000
1!
1%
#486400000000
0!
0%
#486405000000
1!
1%
#486410000000
0!
0%
#486415000000
1!
1%
#486420000000
0!
0%
#486425000000
1!
1%
#486430000000
0!
0%
#486435000000
1!
1%
#486440000000
0!
0%
#486445000000
1!
1%
#486450000000
0!
0%
#486455000000
1!
1%
#486460000000
0!
0%
#486465000000
1!
1%
#486470000000
0!
0%
#486475000000
1!
1%
#486480000000
0!
0%
#486485000000
1!
1%
#486490000000
0!
0%
#486495000000
1!
1%
#486500000000
0!
0%
#486505000000
1!
1%
#486510000000
0!
0%
#486515000000
1!
1%
#486520000000
0!
0%
#486525000000
1!
1%
#486530000000
0!
0%
#486535000000
1!
1%
#486540000000
0!
0%
#486545000000
1!
1%
#486550000000
0!
0%
#486555000000
1!
1%
#486560000000
0!
0%
#486565000000
1!
1%
#486570000000
0!
0%
#486575000000
1!
1%
#486580000000
0!
0%
#486585000000
1!
1%
#486590000000
0!
0%
#486595000000
1!
1%
#486600000000
0!
0%
#486605000000
1!
1%
#486610000000
0!
0%
#486615000000
1!
1%
#486620000000
0!
0%
#486625000000
1!
1%
#486630000000
0!
0%
#486635000000
1!
1%
#486640000000
0!
0%
#486645000000
1!
1%
#486650000000
0!
0%
#486655000000
1!
1%
#486660000000
0!
0%
#486665000000
1!
1%
#486670000000
0!
0%
#486675000000
1!
1%
#486680000000
0!
0%
#486685000000
1!
1%
#486690000000
0!
0%
#486695000000
1!
1%
#486700000000
0!
0%
#486705000000
1!
1%
#486710000000
0!
0%
#486715000000
1!
1%
#486720000000
0!
0%
#486725000000
1!
1%
#486730000000
0!
0%
#486735000000
1!
1%
#486740000000
0!
0%
#486745000000
1!
1%
#486750000000
0!
0%
#486755000000
1!
1%
#486760000000
0!
0%
#486765000000
1!
1%
#486770000000
0!
0%
#486775000000
1!
1%
#486780000000
0!
0%
#486785000000
1!
1%
#486790000000
0!
0%
#486795000000
1!
1%
#486800000000
0!
0%
#486805000000
1!
1%
#486810000000
0!
0%
#486815000000
1!
1%
#486820000000
0!
0%
#486825000000
1!
1%
#486830000000
0!
0%
#486835000000
1!
1%
#486840000000
0!
0%
#486845000000
1!
1%
#486850000000
0!
0%
#486855000000
1!
1%
#486860000000
0!
0%
#486865000000
1!
1%
#486870000000
0!
0%
#486875000000
1!
1%
#486880000000
0!
0%
#486885000000
1!
1%
#486890000000
0!
0%
#486895000000
1!
1%
#486900000000
0!
0%
#486905000000
1!
1%
#486910000000
0!
0%
#486915000000
1!
1%
#486920000000
0!
0%
#486925000000
1!
1%
#486930000000
0!
0%
#486935000000
1!
1%
#486940000000
0!
0%
#486945000000
1!
1%
#486950000000
0!
0%
#486955000000
1!
1%
#486960000000
0!
0%
#486965000000
1!
1%
#486970000000
0!
0%
#486975000000
1!
1%
#486980000000
0!
0%
#486985000000
1!
1%
#486990000000
0!
0%
#486995000000
1!
1%
#487000000000
0!
0%
#487005000000
1!
1%
#487010000000
0!
0%
#487015000000
1!
1%
#487020000000
0!
0%
#487025000000
1!
1%
#487030000000
0!
0%
#487035000000
1!
1%
#487040000000
0!
0%
#487045000000
1!
1%
#487050000000
0!
0%
#487055000000
1!
1%
#487060000000
0!
0%
#487065000000
1!
1%
#487070000000
0!
0%
#487075000000
1!
1%
#487080000000
0!
0%
#487085000000
1!
1%
#487090000000
0!
0%
#487095000000
1!
1%
#487100000000
0!
0%
#487105000000
1!
1%
#487110000000
0!
0%
#487115000000
1!
1%
#487120000000
0!
0%
#487125000000
1!
1%
#487130000000
0!
0%
#487135000000
1!
1%
#487140000000
0!
0%
#487145000000
1!
1%
#487150000000
0!
0%
#487155000000
1!
1%
#487160000000
0!
0%
#487165000000
1!
1%
#487170000000
0!
0%
#487175000000
1!
1%
#487180000000
0!
0%
#487185000000
1!
1%
#487190000000
0!
0%
#487195000000
1!
1%
#487200000000
0!
0%
#487205000000
1!
1%
#487210000000
0!
0%
#487215000000
1!
1%
#487220000000
0!
0%
#487225000000
1!
1%
#487230000000
0!
0%
#487235000000
1!
1%
#487240000000
0!
0%
#487245000000
1!
1%
#487250000000
0!
0%
#487255000000
1!
1%
#487260000000
0!
0%
#487265000000
1!
1%
#487270000000
0!
0%
#487275000000
1!
1%
#487280000000
0!
0%
#487285000000
1!
1%
#487290000000
0!
0%
#487295000000
1!
1%
#487300000000
0!
0%
#487305000000
1!
1%
#487310000000
0!
0%
#487315000000
1!
1%
#487320000000
0!
0%
#487325000000
1!
1%
#487330000000
0!
0%
#487335000000
1!
1%
#487340000000
0!
0%
#487345000000
1!
1%
#487350000000
0!
0%
#487355000000
1!
1%
#487360000000
0!
0%
#487365000000
1!
1%
#487370000000
0!
0%
#487375000000
1!
1%
#487380000000
0!
0%
#487385000000
1!
1%
#487390000000
0!
0%
#487395000000
1!
1%
#487400000000
0!
0%
#487405000000
1!
1%
#487410000000
0!
0%
#487415000000
1!
1%
#487420000000
0!
0%
#487425000000
1!
1%
#487430000000
0!
0%
#487435000000
1!
1%
#487440000000
0!
0%
#487445000000
1!
1%
#487450000000
0!
0%
#487455000000
1!
1%
#487460000000
0!
0%
#487465000000
1!
1%
#487470000000
0!
0%
#487475000000
1!
1%
#487480000000
0!
0%
#487485000000
1!
1%
#487490000000
0!
0%
#487495000000
1!
1%
#487500000000
0!
0%
#487505000000
1!
1%
#487510000000
0!
0%
#487515000000
1!
1%
#487520000000
0!
0%
#487525000000
1!
1%
#487530000000
0!
0%
#487535000000
1!
1%
#487540000000
0!
0%
#487545000000
1!
1%
#487550000000
0!
0%
#487555000000
1!
1%
#487560000000
0!
0%
#487565000000
1!
1%
#487570000000
0!
0%
#487575000000
1!
1%
#487580000000
0!
0%
#487585000000
1!
1%
#487590000000
0!
0%
#487595000000
1!
1%
#487600000000
0!
0%
#487605000000
1!
1%
#487610000000
0!
0%
#487615000000
1!
1%
#487620000000
0!
0%
#487625000000
1!
1%
#487630000000
0!
0%
#487635000000
1!
1%
#487640000000
0!
0%
#487645000000
1!
1%
#487650000000
0!
0%
#487655000000
1!
1%
#487660000000
0!
0%
#487665000000
1!
1%
#487670000000
0!
0%
#487675000000
1!
1%
#487680000000
0!
0%
#487685000000
1!
1%
#487690000000
0!
0%
#487695000000
1!
1%
#487700000000
0!
0%
#487705000000
1!
1%
#487710000000
0!
0%
#487715000000
1!
1%
#487720000000
0!
0%
#487725000000
1!
1%
#487730000000
0!
0%
#487735000000
1!
1%
#487740000000
0!
0%
#487745000000
1!
1%
#487750000000
0!
0%
#487755000000
1!
1%
#487760000000
0!
0%
#487765000000
1!
1%
#487770000000
0!
0%
#487775000000
1!
1%
#487780000000
0!
0%
#487785000000
1!
1%
#487790000000
0!
0%
#487795000000
1!
1%
#487800000000
0!
0%
#487805000000
1!
1%
#487810000000
0!
0%
#487815000000
1!
1%
#487820000000
0!
0%
#487825000000
1!
1%
#487830000000
0!
0%
#487835000000
1!
1%
#487840000000
0!
0%
#487845000000
1!
1%
#487850000000
0!
0%
#487855000000
1!
1%
#487860000000
0!
0%
#487865000000
1!
1%
#487870000000
0!
0%
#487875000000
1!
1%
#487880000000
0!
0%
#487885000000
1!
1%
#487890000000
0!
0%
#487895000000
1!
1%
#487900000000
0!
0%
#487905000000
1!
1%
#487910000000
0!
0%
#487915000000
1!
1%
#487920000000
0!
0%
#487925000000
1!
1%
#487930000000
0!
0%
#487935000000
1!
1%
#487940000000
0!
0%
#487945000000
1!
1%
#487950000000
0!
0%
#487955000000
1!
1%
#487960000000
0!
0%
#487965000000
1!
1%
#487970000000
0!
0%
#487975000000
1!
1%
#487980000000
0!
0%
#487985000000
1!
1%
#487990000000
0!
0%
#487995000000
1!
1%
#488000000000
0!
0%
#488005000000
1!
1%
#488010000000
0!
0%
#488015000000
1!
1%
#488020000000
0!
0%
#488025000000
1!
1%
#488030000000
0!
0%
#488035000000
1!
1%
#488040000000
0!
0%
#488045000000
1!
1%
#488050000000
0!
0%
#488055000000
1!
1%
#488060000000
0!
0%
#488065000000
1!
1%
#488070000000
0!
0%
#488075000000
1!
1%
#488080000000
0!
0%
#488085000000
1!
1%
#488090000000
0!
0%
#488095000000
1!
1%
#488100000000
0!
0%
#488105000000
1!
1%
#488110000000
0!
0%
#488115000000
1!
1%
#488120000000
0!
0%
#488125000000
1!
1%
#488130000000
0!
0%
#488135000000
1!
1%
#488140000000
0!
0%
#488145000000
1!
1%
#488150000000
0!
0%
#488155000000
1!
1%
#488160000000
0!
0%
#488165000000
1!
1%
#488170000000
0!
0%
#488175000000
1!
1%
#488180000000
0!
0%
#488185000000
1!
1%
#488190000000
0!
0%
#488195000000
1!
1%
#488200000000
0!
0%
#488205000000
1!
1%
#488210000000
0!
0%
#488215000000
1!
1%
#488220000000
0!
0%
#488225000000
1!
1%
#488230000000
0!
0%
#488235000000
1!
1%
#488240000000
0!
0%
#488245000000
1!
1%
#488250000000
0!
0%
#488255000000
1!
1%
#488260000000
0!
0%
#488265000000
1!
1%
#488270000000
0!
0%
#488275000000
1!
1%
#488280000000
0!
0%
#488285000000
1!
1%
#488290000000
0!
0%
#488295000000
1!
1%
#488300000000
0!
0%
#488305000000
1!
1%
#488310000000
0!
0%
#488315000000
1!
1%
#488320000000
0!
0%
#488325000000
1!
1%
#488330000000
0!
0%
#488335000000
1!
1%
#488340000000
0!
0%
#488345000000
1!
1%
#488350000000
0!
0%
#488355000000
1!
1%
#488360000000
0!
0%
#488365000000
1!
1%
#488370000000
0!
0%
#488375000000
1!
1%
#488380000000
0!
0%
#488385000000
1!
1%
#488390000000
0!
0%
#488395000000
1!
1%
#488400000000
0!
0%
#488405000000
1!
1%
#488410000000
0!
0%
#488415000000
1!
1%
#488420000000
0!
0%
#488425000000
1!
1%
#488430000000
0!
0%
#488435000000
1!
1%
#488440000000
0!
0%
#488445000000
1!
1%
#488450000000
0!
0%
#488455000000
1!
1%
#488460000000
0!
0%
#488465000000
1!
1%
#488470000000
0!
0%
#488475000000
1!
1%
#488480000000
0!
0%
#488485000000
1!
1%
#488490000000
0!
0%
#488495000000
1!
1%
#488500000000
0!
0%
#488505000000
1!
1%
#488510000000
0!
0%
#488515000000
1!
1%
#488520000000
0!
0%
#488525000000
1!
1%
#488530000000
0!
0%
#488535000000
1!
1%
#488540000000
0!
0%
#488545000000
1!
1%
#488550000000
0!
0%
#488555000000
1!
1%
#488560000000
0!
0%
#488565000000
1!
1%
#488570000000
0!
0%
#488575000000
1!
1%
#488580000000
0!
0%
#488585000000
1!
1%
#488590000000
0!
0%
#488595000000
1!
1%
#488600000000
0!
0%
#488605000000
1!
1%
#488610000000
0!
0%
#488615000000
1!
1%
#488620000000
0!
0%
#488625000000
1!
1%
#488630000000
0!
0%
#488635000000
1!
1%
#488640000000
0!
0%
#488645000000
1!
1%
#488650000000
0!
0%
#488655000000
1!
1%
#488660000000
0!
0%
#488665000000
1!
1%
#488670000000
0!
0%
#488675000000
1!
1%
#488680000000
0!
0%
#488685000000
1!
1%
#488690000000
0!
0%
#488695000000
1!
1%
#488700000000
0!
0%
#488705000000
1!
1%
#488710000000
0!
0%
#488715000000
1!
1%
#488720000000
0!
0%
#488725000000
1!
1%
#488730000000
0!
0%
#488735000000
1!
1%
#488740000000
0!
0%
#488745000000
1!
1%
#488750000000
0!
0%
#488755000000
1!
1%
#488760000000
0!
0%
#488765000000
1!
1%
#488770000000
0!
0%
#488775000000
1!
1%
#488780000000
0!
0%
#488785000000
1!
1%
#488790000000
0!
0%
#488795000000
1!
1%
#488800000000
0!
0%
#488805000000
1!
1%
#488810000000
0!
0%
#488815000000
1!
1%
#488820000000
0!
0%
#488825000000
1!
1%
#488830000000
0!
0%
#488835000000
1!
1%
#488840000000
0!
0%
#488845000000
1!
1%
#488850000000
0!
0%
#488855000000
1!
1%
#488860000000
0!
0%
#488865000000
1!
1%
#488870000000
0!
0%
#488875000000
1!
1%
#488880000000
0!
0%
#488885000000
1!
1%
#488890000000
0!
0%
#488895000000
1!
1%
#488900000000
0!
0%
#488905000000
1!
1%
#488910000000
0!
0%
#488915000000
1!
1%
#488920000000
0!
0%
#488925000000
1!
1%
#488930000000
0!
0%
#488935000000
1!
1%
#488940000000
0!
0%
#488945000000
1!
1%
#488950000000
0!
0%
#488955000000
1!
1%
#488960000000
0!
0%
#488965000000
1!
1%
#488970000000
0!
0%
#488975000000
1!
1%
#488980000000
0!
0%
#488985000000
1!
1%
#488990000000
0!
0%
#488995000000
1!
1%
#489000000000
0!
0%
#489005000000
1!
1%
#489010000000
0!
0%
#489015000000
1!
1%
#489020000000
0!
0%
#489025000000
1!
1%
#489030000000
0!
0%
#489035000000
1!
1%
#489040000000
0!
0%
#489045000000
1!
1%
#489050000000
0!
0%
#489055000000
1!
1%
#489060000000
0!
0%
#489065000000
1!
1%
#489070000000
0!
0%
#489075000000
1!
1%
#489080000000
0!
0%
#489085000000
1!
1%
#489090000000
0!
0%
#489095000000
1!
1%
#489100000000
0!
0%
#489105000000
1!
1%
#489110000000
0!
0%
#489115000000
1!
1%
#489120000000
0!
0%
#489125000000
1!
1%
#489130000000
0!
0%
#489135000000
1!
1%
#489140000000
0!
0%
#489145000000
1!
1%
#489150000000
0!
0%
#489155000000
1!
1%
#489160000000
0!
0%
#489165000000
1!
1%
#489170000000
0!
0%
#489175000000
1!
1%
#489180000000
0!
0%
#489185000000
1!
1%
#489190000000
0!
0%
#489195000000
1!
1%
#489200000000
0!
0%
#489205000000
1!
1%
#489210000000
0!
0%
#489215000000
1!
1%
#489220000000
0!
0%
#489225000000
1!
1%
#489230000000
0!
0%
#489235000000
1!
1%
#489240000000
0!
0%
#489245000000
1!
1%
#489250000000
0!
0%
#489255000000
1!
1%
#489260000000
0!
0%
#489265000000
1!
1%
#489270000000
0!
0%
#489275000000
1!
1%
#489280000000
0!
0%
#489285000000
1!
1%
#489290000000
0!
0%
#489295000000
1!
1%
#489300000000
0!
0%
#489305000000
1!
1%
#489310000000
0!
0%
#489315000000
1!
1%
#489320000000
0!
0%
#489325000000
1!
1%
#489330000000
0!
0%
#489335000000
1!
1%
#489340000000
0!
0%
#489345000000
1!
1%
#489350000000
0!
0%
#489355000000
1!
1%
#489360000000
0!
0%
#489365000000
1!
1%
#489370000000
0!
0%
#489375000000
1!
1%
#489380000000
0!
0%
#489385000000
1!
1%
#489390000000
0!
0%
#489395000000
1!
1%
#489400000000
0!
0%
#489405000000
1!
1%
#489410000000
0!
0%
#489415000000
1!
1%
#489420000000
0!
0%
#489425000000
1!
1%
#489430000000
0!
0%
#489435000000
1!
1%
#489440000000
0!
0%
#489445000000
1!
1%
#489450000000
0!
0%
#489455000000
1!
1%
#489460000000
0!
0%
#489465000000
1!
1%
#489470000000
0!
0%
#489475000000
1!
1%
#489480000000
0!
0%
#489485000000
1!
1%
#489490000000
0!
0%
#489495000000
1!
1%
#489500000000
0!
0%
#489505000000
1!
1%
#489510000000
0!
0%
#489515000000
1!
1%
#489520000000
0!
0%
#489525000000
1!
1%
#489530000000
0!
0%
#489535000000
1!
1%
#489540000000
0!
0%
#489545000000
1!
1%
#489550000000
0!
0%
#489555000000
1!
1%
#489560000000
0!
0%
#489565000000
1!
1%
#489570000000
0!
0%
#489575000000
1!
1%
#489580000000
0!
0%
#489585000000
1!
1%
#489590000000
0!
0%
#489595000000
1!
1%
#489600000000
0!
0%
#489605000000
1!
1%
#489610000000
0!
0%
#489615000000
1!
1%
#489620000000
0!
0%
#489625000000
1!
1%
#489630000000
0!
0%
#489635000000
1!
1%
#489640000000
0!
0%
#489645000000
1!
1%
#489650000000
0!
0%
#489655000000
1!
1%
#489660000000
0!
0%
#489665000000
1!
1%
#489670000000
0!
0%
#489675000000
1!
1%
#489680000000
0!
0%
#489685000000
1!
1%
#489690000000
0!
0%
#489695000000
1!
1%
#489700000000
0!
0%
#489705000000
1!
1%
#489710000000
0!
0%
#489715000000
1!
1%
#489720000000
0!
0%
#489725000000
1!
1%
#489730000000
0!
0%
#489735000000
1!
1%
#489740000000
0!
0%
#489745000000
1!
1%
#489750000000
0!
0%
#489755000000
1!
1%
#489760000000
0!
0%
#489765000000
1!
1%
#489770000000
0!
0%
#489775000000
1!
1%
#489780000000
0!
0%
#489785000000
1!
1%
#489790000000
0!
0%
#489795000000
1!
1%
#489800000000
0!
0%
#489805000000
1!
1%
#489810000000
0!
0%
#489815000000
1!
1%
#489820000000
0!
0%
#489825000000
1!
1%
#489830000000
0!
0%
#489835000000
1!
1%
#489840000000
0!
0%
#489845000000
1!
1%
#489850000000
0!
0%
#489855000000
1!
1%
#489860000000
0!
0%
#489865000000
1!
1%
#489870000000
0!
0%
#489875000000
1!
1%
#489880000000
0!
0%
#489885000000
1!
1%
#489890000000
0!
0%
#489895000000
1!
1%
#489900000000
0!
0%
#489905000000
1!
1%
#489910000000
0!
0%
#489915000000
1!
1%
#489920000000
0!
0%
#489925000000
1!
1%
#489930000000
0!
0%
#489935000000
1!
1%
#489940000000
0!
0%
#489945000000
1!
1%
#489950000000
0!
0%
#489955000000
1!
1%
#489960000000
0!
0%
#489965000000
1!
1%
#489970000000
0!
0%
#489975000000
1!
1%
#489980000000
0!
0%
#489985000000
1!
1%
#489990000000
0!
0%
#489995000000
1!
1%
#490000000000
0!
0%
#490005000000
1!
1%
#490010000000
0!
0%
#490015000000
1!
1%
#490020000000
0!
0%
#490025000000
1!
1%
#490030000000
0!
0%
#490035000000
1!
1%
#490040000000
0!
0%
#490045000000
1!
1%
#490050000000
0!
0%
#490055000000
1!
1%
#490060000000
0!
0%
#490065000000
1!
1%
#490070000000
0!
0%
#490075000000
1!
1%
#490080000000
0!
0%
#490085000000
1!
1%
#490090000000
0!
0%
#490095000000
1!
1%
#490100000000
0!
0%
#490105000000
1!
1%
#490110000000
0!
0%
#490115000000
1!
1%
#490120000000
0!
0%
#490125000000
1!
1%
#490130000000
0!
0%
#490135000000
1!
1%
#490140000000
0!
0%
#490145000000
1!
1%
#490150000000
0!
0%
#490155000000
1!
1%
#490160000000
0!
0%
#490165000000
1!
1%
#490170000000
0!
0%
#490175000000
1!
1%
#490180000000
0!
0%
#490185000000
1!
1%
#490190000000
0!
0%
#490195000000
1!
1%
#490200000000
0!
0%
#490205000000
1!
1%
#490210000000
0!
0%
#490215000000
1!
1%
#490220000000
0!
0%
#490225000000
1!
1%
#490230000000
0!
0%
#490235000000
1!
1%
#490240000000
0!
0%
#490245000000
1!
1%
#490250000000
0!
0%
#490255000000
1!
1%
#490260000000
0!
0%
#490265000000
1!
1%
#490270000000
0!
0%
#490275000000
1!
1%
#490280000000
0!
0%
#490285000000
1!
1%
#490290000000
0!
0%
#490295000000
1!
1%
#490300000000
0!
0%
#490305000000
1!
1%
#490310000000
0!
0%
#490315000000
1!
1%
#490320000000
0!
0%
#490325000000
1!
1%
#490330000000
0!
0%
#490335000000
1!
1%
#490340000000
0!
0%
#490345000000
1!
1%
#490350000000
0!
0%
#490355000000
1!
1%
#490360000000
0!
0%
#490365000000
1!
1%
#490370000000
0!
0%
#490375000000
1!
1%
#490380000000
0!
0%
#490385000000
1!
1%
#490390000000
0!
0%
#490395000000
1!
1%
#490400000000
0!
0%
#490405000000
1!
1%
#490410000000
0!
0%
#490415000000
1!
1%
#490420000000
0!
0%
#490425000000
1!
1%
#490430000000
0!
0%
#490435000000
1!
1%
#490440000000
0!
0%
#490445000000
1!
1%
#490450000000
0!
0%
#490455000000
1!
1%
#490460000000
0!
0%
#490465000000
1!
1%
#490470000000
0!
0%
#490475000000
1!
1%
#490480000000
0!
0%
#490485000000
1!
1%
#490490000000
0!
0%
#490495000000
1!
1%
#490500000000
0!
0%
#490505000000
1!
1%
#490510000000
0!
0%
#490515000000
1!
1%
#490520000000
0!
0%
#490525000000
1!
1%
#490530000000
0!
0%
#490535000000
1!
1%
#490540000000
0!
0%
#490545000000
1!
1%
#490550000000
0!
0%
#490555000000
1!
1%
#490560000000
0!
0%
#490565000000
1!
1%
#490570000000
0!
0%
#490575000000
1!
1%
#490580000000
0!
0%
#490585000000
1!
1%
#490590000000
0!
0%
#490595000000
1!
1%
#490600000000
0!
0%
#490605000000
1!
1%
#490610000000
0!
0%
#490615000000
1!
1%
#490620000000
0!
0%
#490625000000
1!
1%
#490630000000
0!
0%
#490635000000
1!
1%
#490640000000
0!
0%
#490645000000
1!
1%
#490650000000
0!
0%
#490655000000
1!
1%
#490660000000
0!
0%
#490665000000
1!
1%
#490670000000
0!
0%
#490675000000
1!
1%
#490680000000
0!
0%
#490685000000
1!
1%
#490690000000
0!
0%
#490695000000
1!
1%
#490700000000
0!
0%
#490705000000
1!
1%
#490710000000
0!
0%
#490715000000
1!
1%
#490720000000
0!
0%
#490725000000
1!
1%
#490730000000
0!
0%
#490735000000
1!
1%
#490740000000
0!
0%
#490745000000
1!
1%
#490750000000
0!
0%
#490755000000
1!
1%
#490760000000
0!
0%
#490765000000
1!
1%
#490770000000
0!
0%
#490775000000
1!
1%
#490780000000
0!
0%
#490785000000
1!
1%
#490790000000
0!
0%
#490795000000
1!
1%
#490800000000
0!
0%
#490805000000
1!
1%
#490810000000
0!
0%
#490815000000
1!
1%
#490820000000
0!
0%
#490825000000
1!
1%
#490830000000
0!
0%
#490835000000
1!
1%
#490840000000
0!
0%
#490845000000
1!
1%
#490850000000
0!
0%
#490855000000
1!
1%
#490860000000
0!
0%
#490865000000
1!
1%
#490870000000
0!
0%
#490875000000
1!
1%
#490880000000
0!
0%
#490885000000
1!
1%
#490890000000
0!
0%
#490895000000
1!
1%
#490900000000
0!
0%
#490905000000
1!
1%
#490910000000
0!
0%
#490915000000
1!
1%
#490920000000
0!
0%
#490925000000
1!
1%
#490930000000
0!
0%
#490935000000
1!
1%
#490940000000
0!
0%
#490945000000
1!
1%
#490950000000
0!
0%
#490955000000
1!
1%
#490960000000
0!
0%
#490965000000
1!
1%
#490970000000
0!
0%
#490975000000
1!
1%
#490980000000
0!
0%
#490985000000
1!
1%
#490990000000
0!
0%
#490995000000
1!
1%
#491000000000
0!
0%
#491005000000
1!
1%
#491010000000
0!
0%
#491015000000
1!
1%
#491020000000
0!
0%
#491025000000
1!
1%
#491030000000
0!
0%
#491035000000
1!
1%
#491040000000
0!
0%
#491045000000
1!
1%
#491050000000
0!
0%
#491055000000
1!
1%
#491060000000
0!
0%
#491065000000
1!
1%
#491070000000
0!
0%
#491075000000
1!
1%
#491080000000
0!
0%
#491085000000
1!
1%
#491090000000
0!
0%
#491095000000
1!
1%
#491100000000
0!
0%
#491105000000
1!
1%
#491110000000
0!
0%
#491115000000
1!
1%
#491120000000
0!
0%
#491125000000
1!
1%
#491130000000
0!
0%
#491135000000
1!
1%
#491140000000
0!
0%
#491145000000
1!
1%
#491150000000
0!
0%
#491155000000
1!
1%
#491160000000
0!
0%
#491165000000
1!
1%
#491170000000
0!
0%
#491175000000
1!
1%
#491180000000
0!
0%
#491185000000
1!
1%
#491190000000
0!
0%
#491195000000
1!
1%
#491200000000
0!
0%
#491205000000
1!
1%
#491210000000
0!
0%
#491215000000
1!
1%
#491220000000
0!
0%
#491225000000
1!
1%
#491230000000
0!
0%
#491235000000
1!
1%
#491240000000
0!
0%
#491245000000
1!
1%
#491250000000
0!
0%
#491255000000
1!
1%
#491260000000
0!
0%
#491265000000
1!
1%
#491270000000
0!
0%
#491275000000
1!
1%
#491280000000
0!
0%
#491285000000
1!
1%
#491290000000
0!
0%
#491295000000
1!
1%
#491300000000
0!
0%
#491305000000
1!
1%
#491310000000
0!
0%
#491315000000
1!
1%
#491320000000
0!
0%
#491325000000
1!
1%
#491330000000
0!
0%
#491335000000
1!
1%
#491340000000
0!
0%
#491345000000
1!
1%
#491350000000
0!
0%
#491355000000
1!
1%
#491360000000
0!
0%
#491365000000
1!
1%
#491370000000
0!
0%
#491375000000
1!
1%
#491380000000
0!
0%
#491385000000
1!
1%
#491390000000
0!
0%
#491395000000
1!
1%
#491400000000
0!
0%
#491405000000
1!
1%
#491410000000
0!
0%
#491415000000
1!
1%
#491420000000
0!
0%
#491425000000
1!
1%
#491430000000
0!
0%
#491435000000
1!
1%
#491440000000
0!
0%
#491445000000
1!
1%
#491450000000
0!
0%
#491455000000
1!
1%
#491460000000
0!
0%
#491465000000
1!
1%
#491470000000
0!
0%
#491475000000
1!
1%
#491480000000
0!
0%
#491485000000
1!
1%
#491490000000
0!
0%
#491495000000
1!
1%
#491500000000
0!
0%
#491505000000
1!
1%
#491510000000
0!
0%
#491515000000
1!
1%
#491520000000
0!
0%
#491525000000
1!
1%
#491530000000
0!
0%
#491535000000
1!
1%
#491540000000
0!
0%
#491545000000
1!
1%
#491550000000
0!
0%
#491555000000
1!
1%
#491560000000
0!
0%
#491565000000
1!
1%
#491570000000
0!
0%
#491575000000
1!
1%
#491580000000
0!
0%
#491585000000
1!
1%
#491590000000
0!
0%
#491595000000
1!
1%
#491600000000
0!
0%
#491605000000
1!
1%
#491610000000
0!
0%
#491615000000
1!
1%
#491620000000
0!
0%
#491625000000
1!
1%
#491630000000
0!
0%
#491635000000
1!
1%
#491640000000
0!
0%
#491645000000
1!
1%
#491650000000
0!
0%
#491655000000
1!
1%
#491660000000
0!
0%
#491665000000
1!
1%
#491670000000
0!
0%
#491675000000
1!
1%
#491680000000
0!
0%
#491685000000
1!
1%
#491690000000
0!
0%
#491695000000
1!
1%
#491700000000
0!
0%
#491705000000
1!
1%
#491710000000
0!
0%
#491715000000
1!
1%
#491720000000
0!
0%
#491725000000
1!
1%
#491730000000
0!
0%
#491735000000
1!
1%
#491740000000
0!
0%
#491745000000
1!
1%
#491750000000
0!
0%
#491755000000
1!
1%
#491760000000
0!
0%
#491765000000
1!
1%
#491770000000
0!
0%
#491775000000
1!
1%
#491780000000
0!
0%
#491785000000
1!
1%
#491790000000
0!
0%
#491795000000
1!
1%
#491800000000
0!
0%
#491805000000
1!
1%
#491810000000
0!
0%
#491815000000
1!
1%
#491820000000
0!
0%
#491825000000
1!
1%
#491830000000
0!
0%
#491835000000
1!
1%
#491840000000
0!
0%
#491845000000
1!
1%
#491850000000
0!
0%
#491855000000
1!
1%
#491860000000
0!
0%
#491865000000
1!
1%
#491870000000
0!
0%
#491875000000
1!
1%
#491880000000
0!
0%
#491885000000
1!
1%
#491890000000
0!
0%
#491895000000
1!
1%
#491900000000
0!
0%
#491905000000
1!
1%
#491910000000
0!
0%
#491915000000
1!
1%
#491920000000
0!
0%
#491925000000
1!
1%
#491930000000
0!
0%
#491935000000
1!
1%
#491940000000
0!
0%
#491945000000
1!
1%
#491950000000
0!
0%
#491955000000
1!
1%
#491960000000
0!
0%
#491965000000
1!
1%
#491970000000
0!
0%
#491975000000
1!
1%
#491980000000
0!
0%
#491985000000
1!
1%
#491990000000
0!
0%
#491995000000
1!
1%
#492000000000
0!
0%
#492005000000
1!
1%
#492010000000
0!
0%
#492015000000
1!
1%
#492020000000
0!
0%
#492025000000
1!
1%
#492030000000
0!
0%
#492035000000
1!
1%
#492040000000
0!
0%
#492045000000
1!
1%
#492050000000
0!
0%
#492055000000
1!
1%
#492060000000
0!
0%
#492065000000
1!
1%
#492070000000
0!
0%
#492075000000
1!
1%
#492080000000
0!
0%
#492085000000
1!
1%
#492090000000
0!
0%
#492095000000
1!
1%
#492100000000
0!
0%
#492105000000
1!
1%
#492110000000
0!
0%
#492115000000
1!
1%
#492120000000
0!
0%
#492125000000
1!
1%
#492130000000
0!
0%
#492135000000
1!
1%
#492140000000
0!
0%
#492145000000
1!
1%
#492150000000
0!
0%
#492155000000
1!
1%
#492160000000
0!
0%
#492165000000
1!
1%
#492170000000
0!
0%
#492175000000
1!
1%
#492180000000
0!
0%
#492185000000
1!
1%
#492190000000
0!
0%
#492195000000
1!
1%
#492200000000
0!
0%
#492205000000
1!
1%
#492210000000
0!
0%
#492215000000
1!
1%
#492220000000
0!
0%
#492225000000
1!
1%
#492230000000
0!
0%
#492235000000
1!
1%
#492240000000
0!
0%
#492245000000
1!
1%
#492250000000
0!
0%
#492255000000
1!
1%
#492260000000
0!
0%
#492265000000
1!
1%
#492270000000
0!
0%
#492275000000
1!
1%
#492280000000
0!
0%
#492285000000
1!
1%
#492290000000
0!
0%
#492295000000
1!
1%
#492300000000
0!
0%
#492305000000
1!
1%
#492310000000
0!
0%
#492315000000
1!
1%
#492320000000
0!
0%
#492325000000
1!
1%
#492330000000
0!
0%
#492335000000
1!
1%
#492340000000
0!
0%
#492345000000
1!
1%
#492350000000
0!
0%
#492355000000
1!
1%
#492360000000
0!
0%
#492365000000
1!
1%
#492370000000
0!
0%
#492375000000
1!
1%
#492380000000
0!
0%
#492385000000
1!
1%
#492390000000
0!
0%
#492395000000
1!
1%
#492400000000
0!
0%
#492405000000
1!
1%
#492410000000
0!
0%
#492415000000
1!
1%
#492420000000
0!
0%
#492425000000
1!
1%
#492430000000
0!
0%
#492435000000
1!
1%
#492440000000
0!
0%
#492445000000
1!
1%
#492450000000
0!
0%
#492455000000
1!
1%
#492460000000
0!
0%
#492465000000
1!
1%
#492470000000
0!
0%
#492475000000
1!
1%
#492480000000
0!
0%
#492485000000
1!
1%
#492490000000
0!
0%
#492495000000
1!
1%
#492500000000
0!
0%
#492505000000
1!
1%
#492510000000
0!
0%
#492515000000
1!
1%
#492520000000
0!
0%
#492525000000
1!
1%
#492530000000
0!
0%
#492535000000
1!
1%
#492540000000
0!
0%
#492545000000
1!
1%
#492550000000
0!
0%
#492555000000
1!
1%
#492560000000
0!
0%
#492565000000
1!
1%
#492570000000
0!
0%
#492575000000
1!
1%
#492580000000
0!
0%
#492585000000
1!
1%
#492590000000
0!
0%
#492595000000
1!
1%
#492600000000
0!
0%
#492605000000
1!
1%
#492610000000
0!
0%
#492615000000
1!
1%
#492620000000
0!
0%
#492625000000
1!
1%
#492630000000
0!
0%
#492635000000
1!
1%
#492640000000
0!
0%
#492645000000
1!
1%
#492650000000
0!
0%
#492655000000
1!
1%
#492660000000
0!
0%
#492665000000
1!
1%
#492670000000
0!
0%
#492675000000
1!
1%
#492680000000
0!
0%
#492685000000
1!
1%
#492690000000
0!
0%
#492695000000
1!
1%
#492700000000
0!
0%
#492705000000
1!
1%
#492710000000
0!
0%
#492715000000
1!
1%
#492720000000
0!
0%
#492725000000
1!
1%
#492730000000
0!
0%
#492735000000
1!
1%
#492740000000
0!
0%
#492745000000
1!
1%
#492750000000
0!
0%
#492755000000
1!
1%
#492760000000
0!
0%
#492765000000
1!
1%
#492770000000
0!
0%
#492775000000
1!
1%
#492780000000
0!
0%
#492785000000
1!
1%
#492790000000
0!
0%
#492795000000
1!
1%
#492800000000
0!
0%
#492805000000
1!
1%
#492810000000
0!
0%
#492815000000
1!
1%
#492820000000
0!
0%
#492825000000
1!
1%
#492830000000
0!
0%
#492835000000
1!
1%
#492840000000
0!
0%
#492845000000
1!
1%
#492850000000
0!
0%
#492855000000
1!
1%
#492860000000
0!
0%
#492865000000
1!
1%
#492870000000
0!
0%
#492875000000
1!
1%
#492880000000
0!
0%
#492885000000
1!
1%
#492890000000
0!
0%
#492895000000
1!
1%
#492900000000
0!
0%
#492905000000
1!
1%
#492910000000
0!
0%
#492915000000
1!
1%
#492920000000
0!
0%
#492925000000
1!
1%
#492930000000
0!
0%
#492935000000
1!
1%
#492940000000
0!
0%
#492945000000
1!
1%
#492950000000
0!
0%
#492955000000
1!
1%
#492960000000
0!
0%
#492965000000
1!
1%
#492970000000
0!
0%
#492975000000
1!
1%
#492980000000
0!
0%
#492985000000
1!
1%
#492990000000
0!
0%
#492995000000
1!
1%
#493000000000
0!
0%
#493005000000
1!
1%
#493010000000
0!
0%
#493015000000
1!
1%
#493020000000
0!
0%
#493025000000
1!
1%
#493030000000
0!
0%
#493035000000
1!
1%
#493040000000
0!
0%
#493045000000
1!
1%
#493050000000
0!
0%
#493055000000
1!
1%
#493060000000
0!
0%
#493065000000
1!
1%
#493070000000
0!
0%
#493075000000
1!
1%
#493080000000
0!
0%
#493085000000
1!
1%
#493090000000
0!
0%
#493095000000
1!
1%
#493100000000
0!
0%
#493105000000
1!
1%
#493110000000
0!
0%
#493115000000
1!
1%
#493120000000
0!
0%
#493125000000
1!
1%
#493130000000
0!
0%
#493135000000
1!
1%
#493140000000
0!
0%
#493145000000
1!
1%
#493150000000
0!
0%
#493155000000
1!
1%
#493160000000
0!
0%
#493165000000
1!
1%
#493170000000
0!
0%
#493175000000
1!
1%
#493180000000
0!
0%
#493185000000
1!
1%
#493190000000
0!
0%
#493195000000
1!
1%
#493200000000
0!
0%
#493205000000
1!
1%
#493210000000
0!
0%
#493215000000
1!
1%
#493220000000
0!
0%
#493225000000
1!
1%
#493230000000
0!
0%
#493235000000
1!
1%
#493240000000
0!
0%
#493245000000
1!
1%
#493250000000
0!
0%
#493255000000
1!
1%
#493260000000
0!
0%
#493265000000
1!
1%
#493270000000
0!
0%
#493275000000
1!
1%
#493280000000
0!
0%
#493285000000
1!
1%
#493290000000
0!
0%
#493295000000
1!
1%
#493300000000
0!
0%
#493305000000
1!
1%
#493310000000
0!
0%
#493315000000
1!
1%
#493320000000
0!
0%
#493325000000
1!
1%
#493330000000
0!
0%
#493335000000
1!
1%
#493340000000
0!
0%
#493345000000
1!
1%
#493350000000
0!
0%
#493355000000
1!
1%
#493360000000
0!
0%
#493365000000
1!
1%
#493370000000
0!
0%
#493375000000
1!
1%
#493380000000
0!
0%
#493385000000
1!
1%
#493390000000
0!
0%
#493395000000
1!
1%
#493400000000
0!
0%
#493405000000
1!
1%
#493410000000
0!
0%
#493415000000
1!
1%
#493420000000
0!
0%
#493425000000
1!
1%
#493430000000
0!
0%
#493435000000
1!
1%
#493440000000
0!
0%
#493445000000
1!
1%
#493450000000
0!
0%
#493455000000
1!
1%
#493460000000
0!
0%
#493465000000
1!
1%
#493470000000
0!
0%
#493475000000
1!
1%
#493480000000
0!
0%
#493485000000
1!
1%
#493490000000
0!
0%
#493495000000
1!
1%
#493500000000
0!
0%
#493505000000
1!
1%
#493510000000
0!
0%
#493515000000
1!
1%
#493520000000
0!
0%
#493525000000
1!
1%
#493530000000
0!
0%
#493535000000
1!
1%
#493540000000
0!
0%
#493545000000
1!
1%
#493550000000
0!
0%
#493555000000
1!
1%
#493560000000
0!
0%
#493565000000
1!
1%
#493570000000
0!
0%
#493575000000
1!
1%
#493580000000
0!
0%
#493585000000
1!
1%
#493590000000
0!
0%
#493595000000
1!
1%
#493600000000
0!
0%
#493605000000
1!
1%
#493610000000
0!
0%
#493615000000
1!
1%
#493620000000
0!
0%
#493625000000
1!
1%
#493630000000
0!
0%
#493635000000
1!
1%
#493640000000
0!
0%
#493645000000
1!
1%
#493650000000
0!
0%
#493655000000
1!
1%
#493660000000
0!
0%
#493665000000
1!
1%
#493670000000
0!
0%
#493675000000
1!
1%
#493680000000
0!
0%
#493685000000
1!
1%
#493690000000
0!
0%
#493695000000
1!
1%
#493700000000
0!
0%
#493705000000
1!
1%
#493710000000
0!
0%
#493715000000
1!
1%
#493720000000
0!
0%
#493725000000
1!
1%
#493730000000
0!
0%
#493735000000
1!
1%
#493740000000
0!
0%
#493745000000
1!
1%
#493750000000
0!
0%
#493755000000
1!
1%
#493760000000
0!
0%
#493765000000
1!
1%
#493770000000
0!
0%
#493775000000
1!
1%
#493780000000
0!
0%
#493785000000
1!
1%
#493790000000
0!
0%
#493795000000
1!
1%
#493800000000
0!
0%
#493805000000
1!
1%
#493810000000
0!
0%
#493815000000
1!
1%
#493820000000
0!
0%
#493825000000
1!
1%
#493830000000
0!
0%
#493835000000
1!
1%
#493840000000
0!
0%
#493845000000
1!
1%
#493850000000
0!
0%
#493855000000
1!
1%
#493860000000
0!
0%
#493865000000
1!
1%
#493870000000
0!
0%
#493875000000
1!
1%
#493880000000
0!
0%
#493885000000
1!
1%
#493890000000
0!
0%
#493895000000
1!
1%
#493900000000
0!
0%
#493905000000
1!
1%
#493910000000
0!
0%
#493915000000
1!
1%
#493920000000
0!
0%
#493925000000
1!
1%
#493930000000
0!
0%
#493935000000
1!
1%
#493940000000
0!
0%
#493945000000
1!
1%
#493950000000
0!
0%
#493955000000
1!
1%
#493960000000
0!
0%
#493965000000
1!
1%
#493970000000
0!
0%
#493975000000
1!
1%
#493980000000
0!
0%
#493985000000
1!
1%
#493990000000
0!
0%
#493995000000
1!
1%
#494000000000
0!
0%
#494005000000
1!
1%
#494010000000
0!
0%
#494015000000
1!
1%
#494020000000
0!
0%
#494025000000
1!
1%
#494030000000
0!
0%
#494035000000
1!
1%
#494040000000
0!
0%
#494045000000
1!
1%
#494050000000
0!
0%
#494055000000
1!
1%
#494060000000
0!
0%
#494065000000
1!
1%
#494070000000
0!
0%
#494075000000
1!
1%
#494080000000
0!
0%
#494085000000
1!
1%
#494090000000
0!
0%
#494095000000
1!
1%
#494100000000
0!
0%
#494105000000
1!
1%
#494110000000
0!
0%
#494115000000
1!
1%
#494120000000
0!
0%
#494125000000
1!
1%
#494130000000
0!
0%
#494135000000
1!
1%
#494140000000
0!
0%
#494145000000
1!
1%
#494150000000
0!
0%
#494155000000
1!
1%
#494160000000
0!
0%
#494165000000
1!
1%
#494170000000
0!
0%
#494175000000
1!
1%
#494180000000
0!
0%
#494185000000
1!
1%
#494190000000
0!
0%
#494195000000
1!
1%
#494200000000
0!
0%
#494205000000
1!
1%
#494210000000
0!
0%
#494215000000
1!
1%
#494220000000
0!
0%
#494225000000
1!
1%
#494230000000
0!
0%
#494235000000
1!
1%
#494240000000
0!
0%
#494245000000
1!
1%
#494250000000
0!
0%
#494255000000
1!
1%
#494260000000
0!
0%
#494265000000
1!
1%
#494270000000
0!
0%
#494275000000
1!
1%
#494280000000
0!
0%
#494285000000
1!
1%
#494290000000
0!
0%
#494295000000
1!
1%
#494300000000
0!
0%
#494305000000
1!
1%
#494310000000
0!
0%
#494315000000
1!
1%
#494320000000
0!
0%
#494325000000
1!
1%
#494330000000
0!
0%
#494335000000
1!
1%
#494340000000
0!
0%
#494345000000
1!
1%
#494350000000
0!
0%
#494355000000
1!
1%
#494360000000
0!
0%
#494365000000
1!
1%
#494370000000
0!
0%
#494375000000
1!
1%
#494380000000
0!
0%
#494385000000
1!
1%
#494390000000
0!
0%
#494395000000
1!
1%
#494400000000
0!
0%
#494405000000
1!
1%
#494410000000
0!
0%
#494415000000
1!
1%
#494420000000
0!
0%
#494425000000
1!
1%
#494430000000
0!
0%
#494435000000
1!
1%
#494440000000
0!
0%
#494445000000
1!
1%
#494450000000
0!
0%
#494455000000
1!
1%
#494460000000
0!
0%
#494465000000
1!
1%
#494470000000
0!
0%
#494475000000
1!
1%
#494480000000
0!
0%
#494485000000
1!
1%
#494490000000
0!
0%
#494495000000
1!
1%
#494500000000
0!
0%
#494505000000
1!
1%
#494510000000
0!
0%
#494515000000
1!
1%
#494520000000
0!
0%
#494525000000
1!
1%
#494530000000
0!
0%
#494535000000
1!
1%
#494540000000
0!
0%
#494545000000
1!
1%
#494550000000
0!
0%
#494555000000
1!
1%
#494560000000
0!
0%
#494565000000
1!
1%
#494570000000
0!
0%
#494575000000
1!
1%
#494580000000
0!
0%
#494585000000
1!
1%
#494590000000
0!
0%
#494595000000
1!
1%
#494600000000
0!
0%
#494605000000
1!
1%
#494610000000
0!
0%
#494615000000
1!
1%
#494620000000
0!
0%
#494625000000
1!
1%
#494630000000
0!
0%
#494635000000
1!
1%
#494640000000
0!
0%
#494645000000
1!
1%
#494650000000
0!
0%
#494655000000
1!
1%
#494660000000
0!
0%
#494665000000
1!
1%
#494670000000
0!
0%
#494675000000
1!
1%
#494680000000
0!
0%
#494685000000
1!
1%
#494690000000
0!
0%
#494695000000
1!
1%
#494700000000
0!
0%
#494705000000
1!
1%
#494710000000
0!
0%
#494715000000
1!
1%
#494720000000
0!
0%
#494725000000
1!
1%
#494730000000
0!
0%
#494735000000
1!
1%
#494740000000
0!
0%
#494745000000
1!
1%
#494750000000
0!
0%
#494755000000
1!
1%
#494760000000
0!
0%
#494765000000
1!
1%
#494770000000
0!
0%
#494775000000
1!
1%
#494780000000
0!
0%
#494785000000
1!
1%
#494790000000
0!
0%
#494795000000
1!
1%
#494800000000
0!
0%
#494805000000
1!
1%
#494810000000
0!
0%
#494815000000
1!
1%
#494820000000
0!
0%
#494825000000
1!
1%
#494830000000
0!
0%
#494835000000
1!
1%
#494840000000
0!
0%
#494845000000
1!
1%
#494850000000
0!
0%
#494855000000
1!
1%
#494860000000
0!
0%
#494865000000
1!
1%
#494870000000
0!
0%
#494875000000
1!
1%
#494880000000
0!
0%
#494885000000
1!
1%
#494890000000
0!
0%
#494895000000
1!
1%
#494900000000
0!
0%
#494905000000
1!
1%
#494910000000
0!
0%
#494915000000
1!
1%
#494920000000
0!
0%
#494925000000
1!
1%
#494930000000
0!
0%
#494935000000
1!
1%
#494940000000
0!
0%
#494945000000
1!
1%
#494950000000
0!
0%
#494955000000
1!
1%
#494960000000
0!
0%
#494965000000
1!
1%
#494970000000
0!
0%
#494975000000
1!
1%
#494980000000
0!
0%
#494985000000
1!
1%
#494990000000
0!
0%
#494995000000
1!
1%
#495000000000
0!
0%
#495005000000
1!
1%
#495010000000
0!
0%
#495015000000
1!
1%
#495020000000
0!
0%
#495025000000
1!
1%
#495030000000
0!
0%
#495035000000
1!
1%
#495040000000
0!
0%
#495045000000
1!
1%
#495050000000
0!
0%
#495055000000
1!
1%
#495060000000
0!
0%
#495065000000
1!
1%
#495070000000
0!
0%
#495075000000
1!
1%
#495080000000
0!
0%
#495085000000
1!
1%
#495090000000
0!
0%
#495095000000
1!
1%
#495100000000
0!
0%
#495105000000
1!
1%
#495110000000
0!
0%
#495115000000
1!
1%
#495120000000
0!
0%
#495125000000
1!
1%
#495130000000
0!
0%
#495135000000
1!
1%
#495140000000
0!
0%
#495145000000
1!
1%
#495150000000
0!
0%
#495155000000
1!
1%
#495160000000
0!
0%
#495165000000
1!
1%
#495170000000
0!
0%
#495175000000
1!
1%
#495180000000
0!
0%
#495185000000
1!
1%
#495190000000
0!
0%
#495195000000
1!
1%
#495200000000
0!
0%
#495205000000
1!
1%
#495210000000
0!
0%
#495215000000
1!
1%
#495220000000
0!
0%
#495225000000
1!
1%
#495230000000
0!
0%
#495235000000
1!
1%
#495240000000
0!
0%
#495245000000
1!
1%
#495250000000
0!
0%
#495255000000
1!
1%
#495260000000
0!
0%
#495265000000
1!
1%
#495270000000
0!
0%
#495275000000
1!
1%
#495280000000
0!
0%
#495285000000
1!
1%
#495290000000
0!
0%
#495295000000
1!
1%
#495300000000
0!
0%
#495305000000
1!
1%
#495310000000
0!
0%
#495315000000
1!
1%
#495320000000
0!
0%
#495325000000
1!
1%
#495330000000
0!
0%
#495335000000
1!
1%
#495340000000
0!
0%
#495345000000
1!
1%
#495350000000
0!
0%
#495355000000
1!
1%
#495360000000
0!
0%
#495365000000
1!
1%
#495370000000
0!
0%
#495375000000
1!
1%
#495380000000
0!
0%
#495385000000
1!
1%
#495390000000
0!
0%
#495395000000
1!
1%
#495400000000
0!
0%
#495405000000
1!
1%
#495410000000
0!
0%
#495415000000
1!
1%
#495420000000
0!
0%
#495425000000
1!
1%
#495430000000
0!
0%
#495435000000
1!
1%
#495440000000
0!
0%
#495445000000
1!
1%
#495450000000
0!
0%
#495455000000
1!
1%
#495460000000
0!
0%
#495465000000
1!
1%
#495470000000
0!
0%
#495475000000
1!
1%
#495480000000
0!
0%
#495485000000
1!
1%
#495490000000
0!
0%
#495495000000
1!
1%
#495500000000
0!
0%
#495505000000
1!
1%
#495510000000
0!
0%
#495515000000
1!
1%
#495520000000
0!
0%
#495525000000
1!
1%
#495530000000
0!
0%
#495535000000
1!
1%
#495540000000
0!
0%
#495545000000
1!
1%
#495550000000
0!
0%
#495555000000
1!
1%
#495560000000
0!
0%
#495565000000
1!
1%
#495570000000
0!
0%
#495575000000
1!
1%
#495580000000
0!
0%
#495585000000
1!
1%
#495590000000
0!
0%
#495595000000
1!
1%
#495600000000
0!
0%
#495605000000
1!
1%
#495610000000
0!
0%
#495615000000
1!
1%
#495620000000
0!
0%
#495625000000
1!
1%
#495630000000
0!
0%
#495635000000
1!
1%
#495640000000
0!
0%
#495645000000
1!
1%
#495650000000
0!
0%
#495655000000
1!
1%
#495660000000
0!
0%
#495665000000
1!
1%
#495670000000
0!
0%
#495675000000
1!
1%
#495680000000
0!
0%
#495685000000
1!
1%
#495690000000
0!
0%
#495695000000
1!
1%
#495700000000
0!
0%
#495705000000
1!
1%
#495710000000
0!
0%
#495715000000
1!
1%
#495720000000
0!
0%
#495725000000
1!
1%
#495730000000
0!
0%
#495735000000
1!
1%
#495740000000
0!
0%
#495745000000
1!
1%
#495750000000
0!
0%
#495755000000
1!
1%
#495760000000
0!
0%
#495765000000
1!
1%
#495770000000
0!
0%
#495775000000
1!
1%
#495780000000
0!
0%
#495785000000
1!
1%
#495790000000
0!
0%
#495795000000
1!
1%
#495800000000
0!
0%
#495805000000
1!
1%
#495810000000
0!
0%
#495815000000
1!
1%
#495820000000
0!
0%
#495825000000
1!
1%
#495830000000
0!
0%
#495835000000
1!
1%
#495840000000
0!
0%
#495845000000
1!
1%
#495850000000
0!
0%
#495855000000
1!
1%
#495860000000
0!
0%
#495865000000
1!
1%
#495870000000
0!
0%
#495875000000
1!
1%
#495880000000
0!
0%
#495885000000
1!
1%
#495890000000
0!
0%
#495895000000
1!
1%
#495900000000
0!
0%
#495905000000
1!
1%
#495910000000
0!
0%
#495915000000
1!
1%
#495920000000
0!
0%
#495925000000
1!
1%
#495930000000
0!
0%
#495935000000
1!
1%
#495940000000
0!
0%
#495945000000
1!
1%
#495950000000
0!
0%
#495955000000
1!
1%
#495960000000
0!
0%
#495965000000
1!
1%
#495970000000
0!
0%
#495975000000
1!
1%
#495980000000
0!
0%
#495985000000
1!
1%
#495990000000
0!
0%
#495995000000
1!
1%
#496000000000
0!
0%
#496005000000
1!
1%
#496010000000
0!
0%
#496015000000
1!
1%
#496020000000
0!
0%
#496025000000
1!
1%
#496030000000
0!
0%
#496035000000
1!
1%
#496040000000
0!
0%
#496045000000
1!
1%
#496050000000
0!
0%
#496055000000
1!
1%
#496060000000
0!
0%
#496065000000
1!
1%
#496070000000
0!
0%
#496075000000
1!
1%
#496080000000
0!
0%
#496085000000
1!
1%
#496090000000
0!
0%
#496095000000
1!
1%
#496100000000
0!
0%
#496105000000
1!
1%
#496110000000
0!
0%
#496115000000
1!
1%
#496120000000
0!
0%
#496125000000
1!
1%
#496130000000
0!
0%
#496135000000
1!
1%
#496140000000
0!
0%
#496145000000
1!
1%
#496150000000
0!
0%
#496155000000
1!
1%
#496160000000
0!
0%
#496165000000
1!
1%
#496170000000
0!
0%
#496175000000
1!
1%
#496180000000
0!
0%
#496185000000
1!
1%
#496190000000
0!
0%
#496195000000
1!
1%
#496200000000
0!
0%
#496205000000
1!
1%
#496210000000
0!
0%
#496215000000
1!
1%
#496220000000
0!
0%
#496225000000
1!
1%
#496230000000
0!
0%
#496235000000
1!
1%
#496240000000
0!
0%
#496245000000
1!
1%
#496250000000
0!
0%
#496255000000
1!
1%
#496260000000
0!
0%
#496265000000
1!
1%
#496270000000
0!
0%
#496275000000
1!
1%
#496280000000
0!
0%
#496285000000
1!
1%
#496290000000
0!
0%
#496295000000
1!
1%
#496300000000
0!
0%
#496305000000
1!
1%
#496310000000
0!
0%
#496315000000
1!
1%
#496320000000
0!
0%
#496325000000
1!
1%
#496330000000
0!
0%
#496335000000
1!
1%
#496340000000
0!
0%
#496345000000
1!
1%
#496350000000
0!
0%
#496355000000
1!
1%
#496360000000
0!
0%
#496365000000
1!
1%
#496370000000
0!
0%
#496375000000
1!
1%
#496380000000
0!
0%
#496385000000
1!
1%
#496390000000
0!
0%
#496395000000
1!
1%
#496400000000
0!
0%
#496405000000
1!
1%
#496410000000
0!
0%
#496415000000
1!
1%
#496420000000
0!
0%
#496425000000
1!
1%
#496430000000
0!
0%
#496435000000
1!
1%
#496440000000
0!
0%
#496445000000
1!
1%
#496450000000
0!
0%
#496455000000
1!
1%
#496460000000
0!
0%
#496465000000
1!
1%
#496470000000
0!
0%
#496475000000
1!
1%
#496480000000
0!
0%
#496485000000
1!
1%
#496490000000
0!
0%
#496495000000
1!
1%
#496500000000
0!
0%
#496505000000
1!
1%
#496510000000
0!
0%
#496515000000
1!
1%
#496520000000
0!
0%
#496525000000
1!
1%
#496530000000
0!
0%
#496535000000
1!
1%
#496540000000
0!
0%
#496545000000
1!
1%
#496550000000
0!
0%
#496555000000
1!
1%
#496560000000
0!
0%
#496565000000
1!
1%
#496570000000
0!
0%
#496575000000
1!
1%
#496580000000
0!
0%
#496585000000
1!
1%
#496590000000
0!
0%
#496595000000
1!
1%
#496600000000
0!
0%
#496605000000
1!
1%
#496610000000
0!
0%
#496615000000
1!
1%
#496620000000
0!
0%
#496625000000
1!
1%
#496630000000
0!
0%
#496635000000
1!
1%
#496640000000
0!
0%
#496645000000
1!
1%
#496650000000
0!
0%
#496655000000
1!
1%
#496660000000
0!
0%
#496665000000
1!
1%
#496670000000
0!
0%
#496675000000
1!
1%
#496680000000
0!
0%
#496685000000
1!
1%
#496690000000
0!
0%
#496695000000
1!
1%
#496700000000
0!
0%
#496705000000
1!
1%
#496710000000
0!
0%
#496715000000
1!
1%
#496720000000
0!
0%
#496725000000
1!
1%
#496730000000
0!
0%
#496735000000
1!
1%
#496740000000
0!
0%
#496745000000
1!
1%
#496750000000
0!
0%
#496755000000
1!
1%
#496760000000
0!
0%
#496765000000
1!
1%
#496770000000
0!
0%
#496775000000
1!
1%
#496780000000
0!
0%
#496785000000
1!
1%
#496790000000
0!
0%
#496795000000
1!
1%
#496800000000
0!
0%
#496805000000
1!
1%
#496810000000
0!
0%
#496815000000
1!
1%
#496820000000
0!
0%
#496825000000
1!
1%
#496830000000
0!
0%
#496835000000
1!
1%
#496840000000
0!
0%
#496845000000
1!
1%
#496850000000
0!
0%
#496855000000
1!
1%
#496860000000
0!
0%
#496865000000
1!
1%
#496870000000
0!
0%
#496875000000
1!
1%
#496880000000
0!
0%
#496885000000
1!
1%
#496890000000
0!
0%
#496895000000
1!
1%
#496900000000
0!
0%
#496905000000
1!
1%
#496910000000
0!
0%
#496915000000
1!
1%
#496920000000
0!
0%
#496925000000
1!
1%
#496930000000
0!
0%
#496935000000
1!
1%
#496940000000
0!
0%
#496945000000
1!
1%
#496950000000
0!
0%
#496955000000
1!
1%
#496960000000
0!
0%
#496965000000
1!
1%
#496970000000
0!
0%
#496975000000
1!
1%
#496980000000
0!
0%
#496985000000
1!
1%
#496990000000
0!
0%
#496995000000
1!
1%
#497000000000
0!
0%
#497005000000
1!
1%
#497010000000
0!
0%
#497015000000
1!
1%
#497020000000
0!
0%
#497025000000
1!
1%
#497030000000
0!
0%
#497035000000
1!
1%
#497040000000
0!
0%
#497045000000
1!
1%
#497050000000
0!
0%
#497055000000
1!
1%
#497060000000
0!
0%
#497065000000
1!
1%
#497070000000
0!
0%
#497075000000
1!
1%
#497080000000
0!
0%
#497085000000
1!
1%
#497090000000
0!
0%
#497095000000
1!
1%
#497100000000
0!
0%
#497105000000
1!
1%
#497110000000
0!
0%
#497115000000
1!
1%
#497120000000
0!
0%
#497125000000
1!
1%
#497130000000
0!
0%
#497135000000
1!
1%
#497140000000
0!
0%
#497145000000
1!
1%
#497150000000
0!
0%
#497155000000
1!
1%
#497160000000
0!
0%
#497165000000
1!
1%
#497170000000
0!
0%
#497175000000
1!
1%
#497180000000
0!
0%
#497185000000
1!
1%
#497190000000
0!
0%
#497195000000
1!
1%
#497200000000
0!
0%
#497205000000
1!
1%
#497210000000
0!
0%
#497215000000
1!
1%
#497220000000
0!
0%
#497225000000
1!
1%
#497230000000
0!
0%
#497235000000
1!
1%
#497240000000
0!
0%
#497245000000
1!
1%
#497250000000
0!
0%
#497255000000
1!
1%
#497260000000
0!
0%
#497265000000
1!
1%
#497270000000
0!
0%
#497275000000
1!
1%
#497280000000
0!
0%
#497285000000
1!
1%
#497290000000
0!
0%
#497295000000
1!
1%
#497300000000
0!
0%
#497305000000
1!
1%
#497310000000
0!
0%
#497315000000
1!
1%
#497320000000
0!
0%
#497325000000
1!
1%
#497330000000
0!
0%
#497335000000
1!
1%
#497340000000
0!
0%
#497345000000
1!
1%
#497350000000
0!
0%
#497355000000
1!
1%
#497360000000
0!
0%
#497365000000
1!
1%
#497370000000
0!
0%
#497375000000
1!
1%
#497380000000
0!
0%
#497385000000
1!
1%
#497390000000
0!
0%
#497395000000
1!
1%
#497400000000
0!
0%
#497405000000
1!
1%
#497410000000
0!
0%
#497415000000
1!
1%
#497420000000
0!
0%
#497425000000
1!
1%
#497430000000
0!
0%
#497435000000
1!
1%
#497440000000
0!
0%
#497445000000
1!
1%
#497450000000
0!
0%
#497455000000
1!
1%
#497460000000
0!
0%
#497465000000
1!
1%
#497470000000
0!
0%
#497475000000
1!
1%
#497480000000
0!
0%
#497485000000
1!
1%
#497490000000
0!
0%
#497495000000
1!
1%
#497500000000
0!
0%
#497505000000
1!
1%
#497510000000
0!
0%
#497515000000
1!
1%
#497520000000
0!
0%
#497525000000
1!
1%
#497530000000
0!
0%
#497535000000
1!
1%
#497540000000
0!
0%
#497545000000
1!
1%
#497550000000
0!
0%
#497555000000
1!
1%
#497560000000
0!
0%
#497565000000
1!
1%
#497570000000
0!
0%
#497575000000
1!
1%
#497580000000
0!
0%
#497585000000
1!
1%
#497590000000
0!
0%
#497595000000
1!
1%
#497600000000
0!
0%
#497605000000
1!
1%
#497610000000
0!
0%
#497615000000
1!
1%
#497620000000
0!
0%
#497625000000
1!
1%
#497630000000
0!
0%
#497635000000
1!
1%
#497640000000
0!
0%
#497645000000
1!
1%
#497650000000
0!
0%
#497655000000
1!
1%
#497660000000
0!
0%
#497665000000
1!
1%
#497670000000
0!
0%
#497675000000
1!
1%
#497680000000
0!
0%
#497685000000
1!
1%
#497690000000
0!
0%
#497695000000
1!
1%
#497700000000
0!
0%
#497705000000
1!
1%
#497710000000
0!
0%
#497715000000
1!
1%
#497720000000
0!
0%
#497725000000
1!
1%
#497730000000
0!
0%
#497735000000
1!
1%
#497740000000
0!
0%
#497745000000
1!
1%
#497750000000
0!
0%
#497755000000
1!
1%
#497760000000
0!
0%
#497765000000
1!
1%
#497770000000
0!
0%
#497775000000
1!
1%
#497780000000
0!
0%
#497785000000
1!
1%
#497790000000
0!
0%
#497795000000
1!
1%
#497800000000
0!
0%
#497805000000
1!
1%
#497810000000
0!
0%
#497815000000
1!
1%
#497820000000
0!
0%
#497825000000
1!
1%
#497830000000
0!
0%
#497835000000
1!
1%
#497840000000
0!
0%
#497845000000
1!
1%
#497850000000
0!
0%
#497855000000
1!
1%
#497860000000
0!
0%
#497865000000
1!
1%
#497870000000
0!
0%
#497875000000
1!
1%
#497880000000
0!
0%
#497885000000
1!
1%
#497890000000
0!
0%
#497895000000
1!
1%
#497900000000
0!
0%
#497905000000
1!
1%
#497910000000
0!
0%
#497915000000
1!
1%
#497920000000
0!
0%
#497925000000
1!
1%
#497930000000
0!
0%
#497935000000
1!
1%
#497940000000
0!
0%
#497945000000
1!
1%
#497950000000
0!
0%
#497955000000
1!
1%
#497960000000
0!
0%
#497965000000
1!
1%
#497970000000
0!
0%
#497975000000
1!
1%
#497980000000
0!
0%
#497985000000
1!
1%
#497990000000
0!
0%
#497995000000
1!
1%
#498000000000
0!
0%
#498005000000
1!
1%
#498010000000
0!
0%
#498015000000
1!
1%
#498020000000
0!
0%
#498025000000
1!
1%
#498030000000
0!
0%
#498035000000
1!
1%
#498040000000
0!
0%
#498045000000
1!
1%
#498050000000
0!
0%
#498055000000
1!
1%
#498060000000
0!
0%
#498065000000
1!
1%
#498070000000
0!
0%
#498075000000
1!
1%
#498080000000
0!
0%
#498085000000
1!
1%
#498090000000
0!
0%
#498095000000
1!
1%
#498100000000
0!
0%
#498105000000
1!
1%
#498110000000
0!
0%
#498115000000
1!
1%
#498120000000
0!
0%
#498125000000
1!
1%
#498130000000
0!
0%
#498135000000
1!
1%
#498140000000
0!
0%
#498145000000
1!
1%
#498150000000
0!
0%
#498155000000
1!
1%
#498160000000
0!
0%
#498165000000
1!
1%
#498170000000
0!
0%
#498175000000
1!
1%
#498180000000
0!
0%
#498185000000
1!
1%
#498190000000
0!
0%
#498195000000
1!
1%
#498200000000
0!
0%
#498205000000
1!
1%
#498210000000
0!
0%
#498215000000
1!
1%
#498220000000
0!
0%
#498225000000
1!
1%
#498230000000
0!
0%
#498235000000
1!
1%
#498240000000
0!
0%
#498245000000
1!
1%
#498250000000
0!
0%
#498255000000
1!
1%
#498260000000
0!
0%
#498265000000
1!
1%
#498270000000
0!
0%
#498275000000
1!
1%
#498280000000
0!
0%
#498285000000
1!
1%
#498290000000
0!
0%
#498295000000
1!
1%
#498300000000
0!
0%
#498305000000
1!
1%
#498310000000
0!
0%
#498315000000
1!
1%
#498320000000
0!
0%
#498325000000
1!
1%
#498330000000
0!
0%
#498335000000
1!
1%
#498340000000
0!
0%
#498345000000
1!
1%
#498350000000
0!
0%
#498355000000
1!
1%
#498360000000
0!
0%
#498365000000
1!
1%
#498370000000
0!
0%
#498375000000
1!
1%
#498380000000
0!
0%
#498385000000
1!
1%
#498390000000
0!
0%
#498395000000
1!
1%
#498400000000
0!
0%
#498405000000
1!
1%
#498410000000
0!
0%
#498415000000
1!
1%
#498420000000
0!
0%
#498425000000
1!
1%
#498430000000
0!
0%
#498435000000
1!
1%
#498440000000
0!
0%
#498445000000
1!
1%
#498450000000
0!
0%
#498455000000
1!
1%
#498460000000
0!
0%
#498465000000
1!
1%
#498470000000
0!
0%
#498475000000
1!
1%
#498480000000
0!
0%
#498485000000
1!
1%
#498490000000
0!
0%
#498495000000
1!
1%
#498500000000
0!
0%
#498505000000
1!
1%
#498510000000
0!
0%
#498515000000
1!
1%
#498520000000
0!
0%
#498525000000
1!
1%
#498530000000
0!
0%
#498535000000
1!
1%
#498540000000
0!
0%
#498545000000
1!
1%
#498550000000
0!
0%
#498555000000
1!
1%
#498560000000
0!
0%
#498565000000
1!
1%
#498570000000
0!
0%
#498575000000
1!
1%
#498580000000
0!
0%
#498585000000
1!
1%
#498590000000
0!
0%
#498595000000
1!
1%
#498600000000
0!
0%
#498605000000
1!
1%
#498610000000
0!
0%
#498615000000
1!
1%
#498620000000
0!
0%
#498625000000
1!
1%
#498630000000
0!
0%
#498635000000
1!
1%
#498640000000
0!
0%
#498645000000
1!
1%
#498650000000
0!
0%
#498655000000
1!
1%
#498660000000
0!
0%
#498665000000
1!
1%
#498670000000
0!
0%
#498675000000
1!
1%
#498680000000
0!
0%
#498685000000
1!
1%
#498690000000
0!
0%
#498695000000
1!
1%
#498700000000
0!
0%
#498705000000
1!
1%
#498710000000
0!
0%
#498715000000
1!
1%
#498720000000
0!
0%
#498725000000
1!
1%
#498730000000
0!
0%
#498735000000
1!
1%
#498740000000
0!
0%
#498745000000
1!
1%
#498750000000
0!
0%
#498755000000
1!
1%
#498760000000
0!
0%
#498765000000
1!
1%
#498770000000
0!
0%
#498775000000
1!
1%
#498780000000
0!
0%
#498785000000
1!
1%
#498790000000
0!
0%
#498795000000
1!
1%
#498800000000
0!
0%
#498805000000
1!
1%
#498810000000
0!
0%
#498815000000
1!
1%
#498820000000
0!
0%
#498825000000
1!
1%
#498830000000
0!
0%
#498835000000
1!
1%
#498840000000
0!
0%
#498845000000
1!
1%
#498850000000
0!
0%
#498855000000
1!
1%
#498860000000
0!
0%
#498865000000
1!
1%
#498870000000
0!
0%
#498875000000
1!
1%
#498880000000
0!
0%
#498885000000
1!
1%
#498890000000
0!
0%
#498895000000
1!
1%
#498900000000
0!
0%
#498905000000
1!
1%
#498910000000
0!
0%
#498915000000
1!
1%
#498920000000
0!
0%
#498925000000
1!
1%
#498930000000
0!
0%
#498935000000
1!
1%
#498940000000
0!
0%
#498945000000
1!
1%
#498950000000
0!
0%
#498955000000
1!
1%
#498960000000
0!
0%
#498965000000
1!
1%
#498970000000
0!
0%
#498975000000
1!
1%
#498980000000
0!
0%
#498985000000
1!
1%
#498990000000
0!
0%
#498995000000
1!
1%
#499000000000
0!
0%
#499005000000
1!
1%
#499010000000
0!
0%
#499015000000
1!
1%
#499020000000
0!
0%
#499025000000
1!
1%
#499030000000
0!
0%
#499035000000
1!
1%
#499040000000
0!
0%
#499045000000
1!
1%
#499050000000
0!
0%
#499055000000
1!
1%
#499060000000
0!
0%
#499065000000
1!
1%
#499070000000
0!
0%
#499075000000
1!
1%
#499080000000
0!
0%
#499085000000
1!
1%
#499090000000
0!
0%
#499095000000
1!
1%
#499100000000
0!
0%
#499105000000
1!
1%
#499110000000
0!
0%
#499115000000
1!
1%
#499120000000
0!
0%
#499125000000
1!
1%
#499130000000
0!
0%
#499135000000
1!
1%
#499140000000
0!
0%
#499145000000
1!
1%
#499150000000
0!
0%
#499155000000
1!
1%
#499160000000
0!
0%
#499165000000
1!
1%
#499170000000
0!
0%
#499175000000
1!
1%
#499180000000
0!
0%
#499185000000
1!
1%
#499190000000
0!
0%
#499195000000
1!
1%
#499200000000
0!
0%
#499205000000
1!
1%
#499210000000
0!
0%
#499215000000
1!
1%
#499220000000
0!
0%
#499225000000
1!
1%
#499230000000
0!
0%
#499235000000
1!
1%
#499240000000
0!
0%
#499245000000
1!
1%
#499250000000
0!
0%
#499255000000
1!
1%
#499260000000
0!
0%
#499265000000
1!
1%
#499270000000
0!
0%
#499275000000
1!
1%
#499280000000
0!
0%
#499285000000
1!
1%
#499290000000
0!
0%
#499295000000
1!
1%
#499300000000
0!
0%
#499305000000
1!
1%
#499310000000
0!
0%
#499315000000
1!
1%
#499320000000
0!
0%
#499325000000
1!
1%
#499330000000
0!
0%
#499335000000
1!
1%
#499340000000
0!
0%
#499345000000
1!
1%
#499350000000
0!
0%
#499355000000
1!
1%
#499360000000
0!
0%
#499365000000
1!
1%
#499370000000
0!
0%
#499375000000
1!
1%
#499380000000
0!
0%
#499385000000
1!
1%
#499390000000
0!
0%
#499395000000
1!
1%
#499400000000
0!
0%
#499405000000
1!
1%
#499410000000
0!
0%
#499415000000
1!
1%
#499420000000
0!
0%
#499425000000
1!
1%
#499430000000
0!
0%
#499435000000
1!
1%
#499440000000
0!
0%
#499445000000
1!
1%
#499450000000
0!
0%
#499455000000
1!
1%
#499460000000
0!
0%
#499465000000
1!
1%
#499470000000
0!
0%
#499475000000
1!
1%
#499480000000
0!
0%
#499485000000
1!
1%
#499490000000
0!
0%
#499495000000
1!
1%
#499500000000
0!
0%
#499505000000
1!
1%
#499510000000
0!
0%
#499515000000
1!
1%
#499520000000
0!
0%
#499525000000
1!
1%
#499530000000
0!
0%
#499535000000
1!
1%
#499540000000
0!
0%
#499545000000
1!
1%
#499550000000
0!
0%
#499555000000
1!
1%
#499560000000
0!
0%
#499565000000
1!
1%
#499570000000
0!
0%
#499575000000
1!
1%
#499580000000
0!
0%
#499585000000
1!
1%
#499590000000
0!
0%
#499595000000
1!
1%
#499600000000
0!
0%
#499605000000
1!
1%
#499610000000
0!
0%
#499615000000
1!
1%
#499620000000
0!
0%
#499625000000
1!
1%
#499630000000
0!
0%
#499635000000
1!
1%
#499640000000
0!
0%
#499645000000
1!
1%
#499650000000
0!
0%
#499655000000
1!
1%
#499660000000
0!
0%
#499665000000
1!
1%
#499670000000
0!
0%
#499675000000
1!
1%
#499680000000
0!
0%
#499685000000
1!
1%
#499690000000
0!
0%
#499695000000
1!
1%
#499700000000
0!
0%
#499705000000
1!
1%
#499710000000
0!
0%
#499715000000
1!
1%
#499720000000
0!
0%
#499725000000
1!
1%
#499730000000
0!
0%
#499735000000
1!
1%
#499740000000
0!
0%
#499745000000
1!
1%
#499750000000
0!
0%
#499755000000
1!
1%
#499760000000
0!
0%
#499765000000
1!
1%
#499770000000
0!
0%
#499775000000
1!
1%
#499780000000
0!
0%
#499785000000
1!
1%
#499790000000
0!
0%
#499795000000
1!
1%
#499800000000
0!
0%
#499805000000
1!
1%
#499810000000
0!
0%
#499815000000
1!
1%
#499820000000
0!
0%
#499825000000
1!
1%
#499830000000
0!
0%
#499835000000
1!
1%
#499840000000
0!
0%
#499845000000
1!
1%
#499850000000
0!
0%
#499855000000
1!
1%
#499860000000
0!
0%
#499865000000
1!
1%
#499870000000
0!
0%
#499875000000
1!
1%
#499880000000
0!
0%
#499885000000
1!
1%
#499890000000
0!
0%
#499895000000
1!
1%
#499900000000
0!
0%
#499905000000
1!
1%
#499910000000
0!
0%
#499915000000
1!
1%
#499920000000
0!
0%
#499925000000
1!
1%
#499930000000
0!
0%
#499935000000
1!
1%
#499940000000
0!
0%
#499945000000
1!
1%
#499950000000
0!
0%
#499955000000
1!
1%
#499960000000
0!
0%
#499965000000
1!
1%
#499970000000
0!
0%
#499975000000
1!
1%
#499980000000
0!
0%
#499985000000
1!
1%
#499990000000
0!
0%
#499995000000
1!
1%
#500000000000
0!
0%
#500005000000
1!
1%
#500010000000
0!
0%
#500015000000
1!
1%
#500020000000
0!
0%
#500025000000
1!
1%
#500030000000
0!
0%
#500035000000
1!
1%
#500040000000
0!
0%
#500045000000
1!
1%
#500050000000
0!
0%
#500055000000
1!
1%
#500060000000
0!
0%
#500065000000
1!
1%
#500070000000
0!
0%
#500075000000
1!
1%
#500080000000
0!
0%
#500085000000
1!
1%
#500090000000
0!
0%
#500095000000
1!
1%
#500100000000
0!
0%
#500105000000
1!
1%
#500110000000
0!
0%
#500115000000
1!
1%
#500120000000
0!
0%
#500125000000
1!
1%
#500130000000
0!
0%
#500135000000
1!
1%
#500140000000
0!
0%
#500145000000
1!
1%
#500150000000
0!
0%
#500155000000
1!
1%
#500160000000
0!
0%
#500165000000
1!
1%
#500170000000
0!
0%
#500175000000
1!
1%
#500180000000
0!
0%
#500185000000
1!
1%
#500190000000
0!
0%
#500195000000
1!
1%
#500200000000
0!
0%
#500205000000
1!
1%
#500210000000
0!
0%
#500215000000
1!
1%
#500220000000
0!
0%
#500225000000
1!
1%
#500230000000
0!
0%
#500235000000
1!
1%
#500240000000
0!
0%
#500245000000
1!
1%
#500250000000
0!
0%
#500255000000
1!
1%
#500260000000
0!
0%
#500265000000
1!
1%
#500270000000
0!
0%
#500275000000
1!
1%
#500280000000
0!
0%
#500285000000
1!
1%
#500290000000
0!
0%
#500295000000
1!
1%
#500300000000
0!
0%
#500305000000
1!
1%
#500310000000
0!
0%
#500315000000
1!
1%
#500320000000
0!
0%
#500325000000
1!
1%
#500330000000
0!
0%
#500335000000
1!
1%
#500340000000
0!
0%
#500345000000
1!
1%
#500350000000
0!
0%
#500355000000
1!
1%
#500360000000
0!
0%
#500365000000
1!
1%
#500370000000
0!
0%
#500375000000
1!
1%
#500380000000
0!
0%
#500385000000
1!
1%
#500390000000
0!
0%
#500395000000
1!
1%
#500400000000
0!
0%
#500405000000
1!
1%
#500410000000
0!
0%
#500415000000
1!
1%
#500420000000
0!
0%
#500425000000
1!
1%
#500430000000
0!
0%
#500435000000
1!
1%
#500440000000
0!
0%
#500445000000
1!
1%
#500450000000
0!
0%
#500455000000
1!
1%
#500460000000
0!
0%
#500465000000
1!
1%
#500470000000
0!
0%
#500475000000
1!
1%
#500480000000
0!
0%
#500485000000
1!
1%
#500490000000
0!
0%
#500495000000
1!
1%
#500500000000
0!
0%
#500505000000
1!
1%
#500510000000
0!
0%
#500515000000
1!
1%
#500520000000
0!
0%
#500525000000
1!
1%
#500530000000
0!
0%
#500535000000
1!
1%
#500540000000
0!
0%
#500545000000
1!
1%
#500550000000
0!
0%
#500555000000
1!
1%
#500560000000
0!
0%
#500565000000
1!
1%
#500570000000
0!
0%
#500575000000
1!
1%
#500580000000
0!
0%
#500585000000
1!
1%
#500590000000
0!
0%
#500595000000
1!
1%
#500600000000
0!
0%
#500605000000
1!
1%
#500610000000
0!
0%
#500615000000
1!
1%
#500620000000
0!
0%
#500625000000
1!
1%
#500630000000
0!
0%
#500635000000
1!
1%
#500640000000
0!
0%
#500645000000
1!
1%
#500650000000
0!
0%
#500655000000
1!
1%
#500660000000
0!
0%
#500665000000
1!
1%
#500670000000
0!
0%
#500675000000
1!
1%
#500680000000
0!
0%
#500685000000
1!
1%
#500690000000
0!
0%
#500695000000
1!
1%
#500700000000
0!
0%
#500705000000
1!
1%
#500710000000
0!
0%
#500715000000
1!
1%
#500720000000
0!
0%
#500725000000
1!
1%
#500730000000
0!
0%
#500735000000
1!
1%
#500740000000
0!
0%
#500745000000
1!
1%
#500750000000
0!
0%
#500755000000
1!
1%
#500760000000
0!
0%
#500765000000
1!
1%
#500770000000
0!
0%
#500775000000
1!
1%
#500780000000
0!
0%
#500785000000
1!
1%
#500790000000
0!
0%
#500795000000
1!
1%
#500800000000
0!
0%
#500805000000
1!
1%
#500810000000
0!
0%
#500815000000
1!
1%
#500820000000
0!
0%
#500825000000
1!
1%
#500830000000
0!
0%
#500835000000
1!
1%
#500840000000
0!
0%
#500845000000
1!
1%
#500850000000
0!
0%
#500855000000
1!
1%
#500860000000
0!
0%
#500865000000
1!
1%
#500870000000
0!
0%
#500875000000
1!
1%
#500880000000
0!
0%
#500885000000
1!
1%
#500890000000
0!
0%
#500895000000
1!
1%
#500900000000
0!
0%
#500905000000
1!
1%
#500910000000
0!
0%
#500915000000
1!
1%
#500920000000
0!
0%
#500925000000
1!
1%
#500930000000
0!
0%
#500935000000
1!
1%
#500940000000
0!
0%
#500945000000
1!
1%
#500950000000
0!
0%
#500955000000
1!
1%
#500960000000
0!
0%
#500965000000
1!
1%
#500970000000
0!
0%
#500975000000
1!
1%
#500980000000
0!
0%
#500985000000
1!
1%
#500990000000
0!
0%
#500995000000
1!
1%
#501000000000
0!
0%
#501005000000
1!
1%
#501010000000
0!
0%
#501015000000
1!
1%
#501020000000
0!
0%
#501025000000
1!
1%
#501030000000
0!
0%
#501035000000
1!
1%
#501040000000
0!
0%
#501045000000
1!
1%
#501050000000
0!
0%
#501055000000
1!
1%
#501060000000
0!
0%
#501065000000
1!
1%
#501070000000
0!
0%
#501075000000
1!
1%
#501080000000
0!
0%
#501085000000
1!
1%
#501090000000
0!
0%
#501095000000
1!
1%
#501100000000
0!
0%
#501105000000
1!
1%
#501110000000
0!
0%
#501115000000
1!
1%
#501120000000
0!
0%
#501125000000
1!
1%
#501130000000
0!
0%
#501135000000
1!
1%
#501140000000
0!
0%
#501145000000
1!
1%
#501150000000
0!
0%
#501155000000
1!
1%
#501160000000
0!
0%
#501165000000
1!
1%
#501170000000
0!
0%
#501175000000
1!
1%
#501180000000
0!
0%
#501185000000
1!
1%
#501190000000
0!
0%
#501195000000
1!
1%
#501200000000
0!
0%
#501205000000
1!
1%
#501210000000
0!
0%
#501215000000
1!
1%
#501220000000
0!
0%
#501225000000
1!
1%
#501230000000
0!
0%
#501235000000
1!
1%
#501240000000
0!
0%
#501245000000
1!
1%
#501250000000
0!
0%
#501255000000
1!
1%
#501260000000
0!
0%
#501265000000
1!
1%
#501270000000
0!
0%
#501275000000
1!
1%
#501280000000
0!
0%
#501285000000
1!
1%
#501290000000
0!
0%
#501295000000
1!
1%
#501300000000
0!
0%
#501305000000
1!
1%
#501310000000
0!
0%
#501315000000
1!
1%
#501320000000
0!
0%
#501325000000
1!
1%
#501330000000
0!
0%
#501335000000
1!
1%
#501340000000
0!
0%
#501345000000
1!
1%
#501350000000
0!
0%
#501355000000
1!
1%
#501360000000
0!
0%
#501365000000
1!
1%
#501370000000
0!
0%
#501375000000
1!
1%
#501380000000
0!
0%
#501385000000
1!
1%
#501390000000
0!
0%
#501395000000
1!
1%
#501400000000
0!
0%
#501405000000
1!
1%
#501410000000
0!
0%
#501415000000
1!
1%
#501420000000
0!
0%
#501425000000
1!
1%
#501430000000
0!
0%
#501435000000
1!
1%
#501440000000
0!
0%
#501445000000
1!
1%
#501450000000
0!
0%
#501455000000
1!
1%
#501460000000
0!
0%
#501465000000
1!
1%
#501470000000
0!
0%
#501475000000
1!
1%
#501480000000
0!
0%
#501485000000
1!
1%
#501490000000
0!
0%
#501495000000
1!
1%
#501500000000
0!
0%
#501505000000
1!
1%
#501510000000
0!
0%
#501515000000
1!
1%
#501520000000
0!
0%
#501525000000
1!
1%
#501530000000
0!
0%
#501535000000
1!
1%
#501540000000
0!
0%
#501545000000
1!
1%
#501550000000
0!
0%
#501555000000
1!
1%
#501560000000
0!
0%
#501565000000
1!
1%
#501570000000
0!
0%
#501575000000
1!
1%
#501580000000
0!
0%
#501585000000
1!
1%
#501590000000
0!
0%
#501595000000
1!
1%
#501600000000
0!
0%
#501605000000
1!
1%
#501610000000
0!
0%
#501615000000
1!
1%
#501620000000
0!
0%
#501625000000
1!
1%
#501630000000
0!
0%
#501635000000
1!
1%
#501640000000
0!
0%
#501645000000
1!
1%
#501650000000
0!
0%
#501655000000
1!
1%
#501660000000
0!
0%
#501665000000
1!
1%
#501670000000
0!
0%
#501675000000
1!
1%
#501680000000
0!
0%
#501685000000
1!
1%
#501690000000
0!
0%
#501695000000
1!
1%
#501700000000
0!
0%
#501705000000
1!
1%
#501710000000
0!
0%
#501715000000
1!
1%
#501720000000
0!
0%
#501725000000
1!
1%
#501730000000
0!
0%
#501735000000
1!
1%
#501740000000
0!
0%
#501745000000
1!
1%
#501750000000
0!
0%
#501755000000
1!
1%
#501760000000
0!
0%
#501765000000
1!
1%
#501770000000
0!
0%
#501775000000
1!
1%
#501780000000
0!
0%
#501785000000
1!
1%
#501790000000
0!
0%
#501795000000
1!
1%
#501800000000
0!
0%
#501805000000
1!
1%
#501810000000
0!
0%
#501815000000
1!
1%
#501820000000
0!
0%
#501825000000
1!
1%
#501830000000
0!
0%
#501835000000
1!
1%
#501840000000
0!
0%
#501845000000
1!
1%
#501850000000
0!
0%
#501855000000
1!
1%
#501860000000
0!
0%
#501865000000
1!
1%
#501870000000
0!
0%
#501875000000
1!
1%
#501880000000
0!
0%
#501885000000
1!
1%
#501890000000
0!
0%
#501895000000
1!
1%
#501900000000
0!
0%
#501905000000
1!
1%
#501910000000
0!
0%
#501915000000
1!
1%
#501920000000
0!
0%
#501925000000
1!
1%
#501930000000
0!
0%
#501935000000
1!
1%
#501940000000
0!
0%
#501945000000
1!
1%
#501950000000
0!
0%
#501955000000
1!
1%
#501960000000
0!
0%
#501965000000
1!
1%
#501970000000
0!
0%
#501975000000
1!
1%
#501980000000
0!
0%
#501985000000
1!
1%
#501990000000
0!
0%
#501995000000
1!
1%
#502000000000
0!
0%
#502005000000
1!
1%
#502010000000
0!
0%
#502015000000
1!
1%
#502020000000
0!
0%
#502025000000
1!
1%
#502030000000
0!
0%
#502035000000
1!
1%
#502040000000
0!
0%
#502045000000
1!
1%
#502050000000
0!
0%
#502055000000
1!
1%
#502060000000
0!
0%
#502065000000
1!
1%
#502070000000
0!
0%
#502075000000
1!
1%
#502080000000
0!
0%
#502085000000
1!
1%
#502090000000
0!
0%
#502095000000
1!
1%
#502100000000
0!
0%
#502105000000
1!
1%
#502110000000
0!
0%
#502115000000
1!
1%
#502120000000
0!
0%
#502125000000
1!
1%
#502130000000
0!
0%
#502135000000
1!
1%
#502140000000
0!
0%
#502145000000
1!
1%
#502150000000
0!
0%
#502155000000
1!
1%
#502160000000
0!
0%
#502165000000
1!
1%
#502170000000
0!
0%
#502175000000
1!
1%
#502180000000
0!
0%
#502185000000
1!
1%
#502190000000
0!
0%
#502195000000
1!
1%
#502200000000
0!
0%
#502205000000
1!
1%
#502210000000
0!
0%
#502215000000
1!
1%
#502220000000
0!
0%
#502225000000
1!
1%
#502230000000
0!
0%
#502235000000
1!
1%
#502240000000
0!
0%
#502245000000
1!
1%
#502250000000
0!
0%
#502255000000
1!
1%
#502260000000
0!
0%
#502265000000
1!
1%
#502270000000
0!
0%
#502275000000
1!
1%
#502280000000
0!
0%
#502285000000
1!
1%
#502290000000
0!
0%
#502295000000
1!
1%
#502300000000
0!
0%
#502305000000
1!
1%
#502310000000
0!
0%
#502315000000
1!
1%
#502320000000
0!
0%
#502325000000
1!
1%
#502330000000
0!
0%
#502335000000
1!
1%
#502340000000
0!
0%
#502345000000
1!
1%
#502350000000
0!
0%
#502355000000
1!
1%
#502360000000
0!
0%
#502365000000
1!
1%
#502370000000
0!
0%
#502375000000
1!
1%
#502380000000
0!
0%
#502385000000
1!
1%
#502390000000
0!
0%
#502395000000
1!
1%
#502400000000
0!
0%
#502405000000
1!
1%
#502410000000
0!
0%
#502415000000
1!
1%
#502420000000
0!
0%
#502425000000
1!
1%
#502430000000
0!
0%
#502435000000
1!
1%
#502440000000
0!
0%
#502445000000
1!
1%
#502450000000
0!
0%
#502455000000
1!
1%
#502460000000
0!
0%
#502465000000
1!
1%
#502470000000
0!
0%
#502475000000
1!
1%
#502480000000
0!
0%
#502485000000
1!
1%
#502490000000
0!
0%
#502495000000
1!
1%
#502500000000
0!
0%
#502505000000
1!
1%
#502510000000
0!
0%
#502515000000
1!
1%
#502520000000
0!
0%
#502525000000
1!
1%
#502530000000
0!
0%
#502535000000
1!
1%
#502540000000
0!
0%
#502545000000
1!
1%
#502550000000
0!
0%
#502555000000
1!
1%
#502560000000
0!
0%
#502565000000
1!
1%
#502570000000
0!
0%
#502575000000
1!
1%
#502580000000
0!
0%
#502585000000
1!
1%
#502590000000
0!
0%
#502595000000
1!
1%
#502600000000
0!
0%
#502605000000
1!
1%
#502610000000
0!
0%
#502615000000
1!
1%
#502620000000
0!
0%
#502625000000
1!
1%
#502630000000
0!
0%
#502635000000
1!
1%
#502640000000
0!
0%
#502645000000
1!
1%
#502650000000
0!
0%
#502655000000
1!
1%
#502660000000
0!
0%
#502665000000
1!
1%
#502670000000
0!
0%
#502675000000
1!
1%
#502680000000
0!
0%
#502685000000
1!
1%
#502690000000
0!
0%
#502695000000
1!
1%
#502700000000
0!
0%
#502705000000
1!
1%
#502710000000
0!
0%
#502715000000
1!
1%
#502720000000
0!
0%
#502725000000
1!
1%
#502730000000
0!
0%
#502735000000
1!
1%
#502740000000
0!
0%
#502745000000
1!
1%
#502750000000
0!
0%
#502755000000
1!
1%
#502760000000
0!
0%
#502765000000
1!
1%
#502770000000
0!
0%
#502775000000
1!
1%
#502780000000
0!
0%
#502785000000
1!
1%
#502790000000
0!
0%
#502795000000
1!
1%
#502800000000
0!
0%
#502805000000
1!
1%
#502810000000
0!
0%
#502815000000
1!
1%
#502820000000
0!
0%
#502825000000
1!
1%
#502830000000
0!
0%
#502835000000
1!
1%
#502840000000
0!
0%
#502845000000
1!
1%
#502850000000
0!
0%
#502855000000
1!
1%
#502860000000
0!
0%
#502865000000
1!
1%
#502870000000
0!
0%
#502875000000
1!
1%
#502880000000
0!
0%
#502885000000
1!
1%
#502890000000
0!
0%
#502895000000
1!
1%
#502900000000
0!
0%
#502905000000
1!
1%
#502910000000
0!
0%
#502915000000
1!
1%
#502920000000
0!
0%
#502925000000
1!
1%
#502930000000
0!
0%
#502935000000
1!
1%
#502940000000
0!
0%
#502945000000
1!
1%
#502950000000
0!
0%
#502955000000
1!
1%
#502960000000
0!
0%
#502965000000
1!
1%
#502970000000
0!
0%
#502975000000
1!
1%
#502980000000
0!
0%
#502985000000
1!
1%
#502990000000
0!
0%
#502995000000
1!
1%
#503000000000
0!
0%
#503005000000
1!
1%
#503010000000
0!
0%
#503015000000
1!
1%
#503020000000
0!
0%
#503025000000
1!
1%
#503030000000
0!
0%
#503035000000
1!
1%
#503040000000
0!
0%
#503045000000
1!
1%
#503050000000
0!
0%
#503055000000
1!
1%
#503060000000
0!
0%
#503065000000
1!
1%
#503070000000
0!
0%
#503075000000
1!
1%
#503080000000
0!
0%
#503085000000
1!
1%
#503090000000
0!
0%
#503095000000
1!
1%
#503100000000
0!
0%
#503105000000
1!
1%
#503110000000
0!
0%
#503115000000
1!
1%
#503120000000
0!
0%
#503125000000
1!
1%
#503130000000
0!
0%
#503135000000
1!
1%
#503140000000
0!
0%
#503145000000
1!
1%
#503150000000
0!
0%
#503155000000
1!
1%
#503160000000
0!
0%
#503165000000
1!
1%
#503170000000
0!
0%
#503175000000
1!
1%
#503180000000
0!
0%
#503185000000
1!
1%
#503190000000
0!
0%
#503195000000
1!
1%
#503200000000
0!
0%
#503205000000
1!
1%
#503210000000
0!
0%
#503215000000
1!
1%
#503220000000
0!
0%
#503225000000
1!
1%
#503230000000
0!
0%
#503235000000
1!
1%
#503240000000
0!
0%
#503245000000
1!
1%
#503250000000
0!
0%
#503255000000
1!
1%
#503260000000
0!
0%
#503265000000
1!
1%
#503270000000
0!
0%
#503275000000
1!
1%
#503280000000
0!
0%
#503285000000
1!
1%
#503290000000
0!
0%
#503295000000
1!
1%
#503300000000
0!
0%
#503305000000
1!
1%
#503310000000
0!
0%
#503315000000
1!
1%
#503320000000
0!
0%
#503325000000
1!
1%
#503330000000
0!
0%
#503335000000
1!
1%
#503340000000
0!
0%
#503345000000
1!
1%
#503350000000
0!
0%
#503355000000
1!
1%
#503360000000
0!
0%
#503365000000
1!
1%
#503370000000
0!
0%
#503375000000
1!
1%
#503380000000
0!
0%
#503385000000
1!
1%
#503390000000
0!
0%
#503395000000
1!
1%
#503400000000
0!
0%
#503405000000
1!
1%
#503410000000
0!
0%
#503415000000
1!
1%
#503420000000
0!
0%
#503425000000
1!
1%
#503430000000
0!
0%
#503435000000
1!
1%
#503440000000
0!
0%
#503445000000
1!
1%
#503450000000
0!
0%
#503455000000
1!
1%
#503460000000
0!
0%
#503465000000
1!
1%
#503470000000
0!
0%
#503475000000
1!
1%
#503480000000
0!
0%
#503485000000
1!
1%
#503490000000
0!
0%
#503495000000
1!
1%
#503500000000
0!
0%
#503505000000
1!
1%
#503510000000
0!
0%
#503515000000
1!
1%
#503520000000
0!
0%
#503525000000
1!
1%
#503530000000
0!
0%
#503535000000
1!
1%
#503540000000
0!
0%
#503545000000
1!
1%
#503550000000
0!
0%
#503555000000
1!
1%
#503560000000
0!
0%
#503565000000
1!
1%
#503570000000
0!
0%
#503575000000
1!
1%
#503580000000
0!
0%
#503585000000
1!
1%
#503590000000
0!
0%
#503595000000
1!
1%
#503600000000
0!
0%
#503605000000
1!
1%
#503610000000
0!
0%
#503615000000
1!
1%
#503620000000
0!
0%
#503625000000
1!
1%
#503630000000
0!
0%
#503635000000
1!
1%
#503640000000
0!
0%
#503645000000
1!
1%
#503650000000
0!
0%
#503655000000
1!
1%
#503660000000
0!
0%
#503665000000
1!
1%
#503670000000
0!
0%
#503675000000
1!
1%
#503680000000
0!
0%
#503685000000
1!
1%
#503690000000
0!
0%
#503695000000
1!
1%
#503700000000
0!
0%
#503705000000
1!
1%
#503710000000
0!
0%
#503715000000
1!
1%
#503720000000
0!
0%
#503725000000
1!
1%
#503730000000
0!
0%
#503735000000
1!
1%
#503740000000
0!
0%
#503745000000
1!
1%
#503750000000
0!
0%
#503755000000
1!
1%
#503760000000
0!
0%
#503765000000
1!
1%
#503770000000
0!
0%
#503775000000
1!
1%
#503780000000
0!
0%
#503785000000
1!
1%
#503790000000
0!
0%
#503795000000
1!
1%
#503800000000
0!
0%
#503805000000
1!
1%
#503810000000
0!
0%
#503815000000
1!
1%
#503820000000
0!
0%
#503825000000
1!
1%
#503830000000
0!
0%
#503835000000
1!
1%
#503840000000
0!
0%
#503845000000
1!
1%
#503850000000
0!
0%
#503855000000
1!
1%
#503860000000
0!
0%
#503865000000
1!
1%
#503870000000
0!
0%
#503875000000
1!
1%
#503880000000
0!
0%
#503885000000
1!
1%
#503890000000
0!
0%
#503895000000
1!
1%
#503900000000
0!
0%
#503905000000
1!
1%
#503910000000
0!
0%
#503915000000
1!
1%
#503920000000
0!
0%
#503925000000
1!
1%
#503930000000
0!
0%
#503935000000
1!
1%
#503940000000
0!
0%
#503945000000
1!
1%
#503950000000
0!
0%
#503955000000
1!
1%
#503960000000
0!
0%
#503965000000
1!
1%
#503970000000
0!
0%
#503975000000
1!
1%
#503980000000
0!
0%
#503985000000
1!
1%
#503990000000
0!
0%
#503995000000
1!
1%
#504000000000
0!
0%
#504005000000
1!
1%
#504010000000
0!
0%
#504015000000
1!
1%
#504020000000
0!
0%
#504025000000
1!
1%
#504030000000
0!
0%
#504035000000
1!
1%
#504040000000
0!
0%
#504045000000
1!
1%
#504050000000
0!
0%
#504055000000
1!
1%
#504060000000
0!
0%
#504065000000
1!
1%
#504070000000
0!
0%
#504075000000
1!
1%
#504080000000
0!
0%
#504085000000
1!
1%
#504090000000
0!
0%
#504095000000
1!
1%
#504100000000
0!
0%
#504105000000
1!
1%
#504110000000
0!
0%
#504115000000
1!
1%
#504120000000
0!
0%
#504125000000
1!
1%
#504130000000
0!
0%
#504135000000
1!
1%
#504140000000
0!
0%
#504145000000
1!
1%
#504150000000
0!
0%
#504155000000
1!
1%
#504160000000
0!
0%
#504165000000
1!
1%
#504170000000
0!
0%
#504175000000
1!
1%
#504180000000
0!
0%
#504185000000
1!
1%
#504190000000
0!
0%
#504195000000
1!
1%
#504200000000
0!
0%
#504205000000
1!
1%
#504210000000
0!
0%
#504215000000
1!
1%
#504220000000
0!
0%
#504225000000
1!
1%
#504230000000
0!
0%
#504235000000
1!
1%
#504240000000
0!
0%
#504245000000
1!
1%
#504250000000
0!
0%
#504255000000
1!
1%
#504260000000
0!
0%
#504265000000
1!
1%
#504270000000
0!
0%
#504275000000
1!
1%
#504280000000
0!
0%
#504285000000
1!
1%
#504290000000
0!
0%
#504295000000
1!
1%
#504300000000
0!
0%
#504305000000
1!
1%
#504310000000
0!
0%
#504315000000
1!
1%
#504320000000
0!
0%
#504325000000
1!
1%
#504330000000
0!
0%
#504335000000
1!
1%
#504340000000
0!
0%
#504345000000
1!
1%
#504350000000
0!
0%
#504355000000
1!
1%
#504360000000
0!
0%
#504365000000
1!
1%
#504370000000
0!
0%
#504375000000
1!
1%
#504380000000
0!
0%
#504385000000
1!
1%
#504390000000
0!
0%
#504395000000
1!
1%
#504400000000
0!
0%
#504405000000
1!
1%
#504410000000
0!
0%
#504415000000
1!
1%
#504420000000
0!
0%
#504425000000
1!
1%
#504430000000
0!
0%
#504435000000
1!
1%
#504440000000
0!
0%
#504445000000
1!
1%
#504450000000
0!
0%
#504455000000
1!
1%
#504460000000
0!
0%
#504465000000
1!
1%
#504470000000
0!
0%
#504475000000
1!
1%
#504480000000
0!
0%
#504485000000
1!
1%
#504490000000
0!
0%
#504495000000
1!
1%
#504500000000
0!
0%
#504505000000
1!
1%
#504510000000
0!
0%
#504515000000
1!
1%
#504520000000
0!
0%
#504525000000
1!
1%
#504530000000
0!
0%
#504535000000
1!
1%
#504540000000
0!
0%
#504545000000
1!
1%
#504550000000
0!
0%
#504555000000
1!
1%
#504560000000
0!
0%
#504565000000
1!
1%
#504570000000
0!
0%
#504575000000
1!
1%
#504580000000
0!
0%
#504585000000
1!
1%
#504590000000
0!
0%
#504595000000
1!
1%
#504600000000
0!
0%
#504605000000
1!
1%
#504610000000
0!
0%
#504615000000
1!
1%
#504620000000
0!
0%
#504625000000
1!
1%
#504630000000
0!
0%
#504635000000
1!
1%
#504640000000
0!
0%
#504645000000
1!
1%
#504650000000
0!
0%
#504655000000
1!
1%
#504660000000
0!
0%
#504665000000
1!
1%
#504670000000
0!
0%
#504675000000
1!
1%
#504680000000
0!
0%
#504685000000
1!
1%
#504690000000
0!
0%
#504695000000
1!
1%
#504700000000
0!
0%
#504705000000
1!
1%
#504710000000
0!
0%
#504715000000
1!
1%
#504720000000
0!
0%
#504725000000
1!
1%
#504730000000
0!
0%
#504735000000
1!
1%
#504740000000
0!
0%
#504745000000
1!
1%
#504750000000
0!
0%
#504755000000
1!
1%
#504760000000
0!
0%
#504765000000
1!
1%
#504770000000
0!
0%
#504775000000
1!
1%
#504780000000
0!
0%
#504785000000
1!
1%
#504790000000
0!
0%
#504795000000
1!
1%
#504800000000
0!
0%
#504805000000
1!
1%
#504810000000
0!
0%
#504815000000
1!
1%
#504820000000
0!
0%
#504825000000
1!
1%
#504830000000
0!
0%
#504835000000
1!
1%
#504840000000
0!
0%
#504845000000
1!
1%
#504850000000
0!
0%
#504855000000
1!
1%
#504860000000
0!
0%
#504865000000
1!
1%
#504870000000
0!
0%
#504875000000
1!
1%
#504880000000
0!
0%
#504885000000
1!
1%
#504890000000
0!
0%
#504895000000
1!
1%
#504900000000
0!
0%
#504905000000
1!
1%
#504910000000
0!
0%
#504915000000
1!
1%
#504920000000
0!
0%
#504925000000
1!
1%
#504930000000
0!
0%
#504935000000
1!
1%
#504940000000
0!
0%
#504945000000
1!
1%
#504950000000
0!
0%
#504955000000
1!
1%
#504960000000
0!
0%
#504965000000
1!
1%
#504970000000
0!
0%
#504975000000
1!
1%
#504980000000
0!
0%
#504985000000
1!
1%
#504990000000
0!
0%
#504995000000
1!
1%
#505000000000
0!
0%
#505005000000
1!
1%
#505010000000
0!
0%
#505015000000
1!
1%
#505020000000
0!
0%
#505025000000
1!
1%
#505030000000
0!
0%
#505035000000
1!
1%
#505040000000
0!
0%
#505045000000
1!
1%
#505050000000
0!
0%
#505055000000
1!
1%
#505060000000
0!
0%
#505065000000
1!
1%
#505070000000
0!
0%
#505075000000
1!
1%
#505080000000
0!
0%
#505085000000
1!
1%
#505090000000
0!
0%
#505095000000
1!
1%
#505100000000
0!
0%
#505105000000
1!
1%
#505110000000
0!
0%
#505115000000
1!
1%
#505120000000
0!
0%
#505125000000
1!
1%
#505130000000
0!
0%
#505135000000
1!
1%
#505140000000
0!
0%
#505145000000
1!
1%
#505150000000
0!
0%
#505155000000
1!
1%
#505160000000
0!
0%
#505165000000
1!
1%
#505170000000
0!
0%
#505175000000
1!
1%
#505180000000
0!
0%
#505185000000
1!
1%
#505190000000
0!
0%
#505195000000
1!
1%
#505200000000
0!
0%
#505205000000
1!
1%
#505210000000
0!
0%
#505215000000
1!
1%
#505220000000
0!
0%
#505225000000
1!
1%
#505230000000
0!
0%
#505235000000
1!
1%
#505240000000
0!
0%
#505245000000
1!
1%
#505250000000
0!
0%
#505255000000
1!
1%
#505260000000
0!
0%
#505265000000
1!
1%
#505270000000
0!
0%
#505275000000
1!
1%
#505280000000
0!
0%
#505285000000
1!
1%
#505290000000
0!
0%
#505295000000
1!
1%
#505300000000
0!
0%
#505305000000
1!
1%
#505310000000
0!
0%
#505315000000
1!
1%
#505320000000
0!
0%
#505325000000
1!
1%
#505330000000
0!
0%
#505335000000
1!
1%
#505340000000
0!
0%
#505345000000
1!
1%
#505350000000
0!
0%
#505355000000
1!
1%
#505360000000
0!
0%
#505365000000
1!
1%
#505370000000
0!
0%
#505375000000
1!
1%
#505380000000
0!
0%
#505385000000
1!
1%
#505390000000
0!
0%
#505395000000
1!
1%
#505400000000
0!
0%
#505405000000
1!
1%
#505410000000
0!
0%
#505415000000
1!
1%
#505420000000
0!
0%
#505425000000
1!
1%
#505430000000
0!
0%
#505435000000
1!
1%
#505440000000
0!
0%
#505445000000
1!
1%
#505450000000
0!
0%
#505455000000
1!
1%
#505460000000
0!
0%
#505465000000
1!
1%
#505470000000
0!
0%
#505475000000
1!
1%
#505480000000
0!
0%
#505485000000
1!
1%
#505490000000
0!
0%
#505495000000
1!
1%
#505500000000
0!
0%
#505505000000
1!
1%
#505510000000
0!
0%
#505515000000
1!
1%
#505520000000
0!
0%
#505525000000
1!
1%
#505530000000
0!
0%
#505535000000
1!
1%
#505540000000
0!
0%
#505545000000
1!
1%
#505550000000
0!
0%
#505555000000
1!
1%
#505560000000
0!
0%
#505565000000
1!
1%
#505570000000
0!
0%
#505575000000
1!
1%
#505580000000
0!
0%
#505585000000
1!
1%
#505590000000
0!
0%
#505595000000
1!
1%
#505600000000
0!
0%
#505605000000
1!
1%
#505610000000
0!
0%
#505615000000
1!
1%
#505620000000
0!
0%
#505625000000
1!
1%
#505630000000
0!
0%
#505635000000
1!
1%
#505640000000
0!
0%
#505645000000
1!
1%
#505650000000
0!
0%
#505655000000
1!
1%
#505660000000
0!
0%
#505665000000
1!
1%
#505670000000
0!
0%
#505675000000
1!
1%
#505680000000
0!
0%
#505685000000
1!
1%
#505690000000
0!
0%
#505695000000
1!
1%
#505700000000
0!
0%
#505705000000
1!
1%
#505710000000
0!
0%
#505715000000
1!
1%
#505720000000
0!
0%
#505725000000
1!
1%
#505730000000
0!
0%
#505735000000
1!
1%
#505740000000
0!
0%
#505745000000
1!
1%
#505750000000
0!
0%
#505755000000
1!
1%
#505760000000
0!
0%
#505765000000
1!
1%
#505770000000
0!
0%
#505775000000
1!
1%
#505780000000
0!
0%
#505785000000
1!
1%
#505790000000
0!
0%
#505795000000
1!
1%
#505800000000
0!
0%
#505805000000
1!
1%
#505810000000
0!
0%
#505815000000
1!
1%
#505820000000
0!
0%
#505825000000
1!
1%
#505830000000
0!
0%
#505835000000
1!
1%
#505840000000
0!
0%
#505845000000
1!
1%
#505850000000
0!
0%
#505855000000
1!
1%
#505860000000
0!
0%
#505865000000
1!
1%
#505870000000
0!
0%
#505875000000
1!
1%
#505880000000
0!
0%
#505885000000
1!
1%
#505890000000
0!
0%
#505895000000
1!
1%
#505900000000
0!
0%
#505905000000
1!
1%
#505910000000
0!
0%
#505915000000
1!
1%
#505920000000
0!
0%
#505925000000
1!
1%
#505930000000
0!
0%
#505935000000
1!
1%
#505940000000
0!
0%
#505945000000
1!
1%
#505950000000
0!
0%
#505955000000
1!
1%
#505960000000
0!
0%
#505965000000
1!
1%
#505970000000
0!
0%
#505975000000
1!
1%
#505980000000
0!
0%
#505985000000
1!
1%
#505990000000
0!
0%
#505995000000
1!
1%
#506000000000
0!
0%
#506005000000
1!
1%
#506010000000
0!
0%
#506015000000
1!
1%
#506020000000
0!
0%
#506025000000
1!
1%
#506030000000
0!
0%
#506035000000
1!
1%
#506040000000
0!
0%
#506045000000
1!
1%
#506050000000
0!
0%
#506055000000
1!
1%
#506060000000
0!
0%
#506065000000
1!
1%
#506070000000
0!
0%
#506075000000
1!
1%
#506080000000
0!
0%
#506085000000
1!
1%
#506090000000
0!
0%
#506095000000
1!
1%
#506100000000
0!
0%
#506105000000
1!
1%
#506110000000
0!
0%
#506115000000
1!
1%
#506120000000
0!
0%
#506125000000
1!
1%
#506130000000
0!
0%
#506135000000
1!
1%
#506140000000
0!
0%
#506145000000
1!
1%
#506150000000
0!
0%
#506155000000
1!
1%
#506160000000
0!
0%
#506165000000
1!
1%
#506170000000
0!
0%
#506175000000
1!
1%
#506180000000
0!
0%
#506185000000
1!
1%
#506190000000
0!
0%
#506195000000
1!
1%
#506200000000
0!
0%
#506205000000
1!
1%
#506210000000
0!
0%
#506215000000
1!
1%
#506220000000
0!
0%
#506225000000
1!
1%
#506230000000
0!
0%
#506235000000
1!
1%
#506240000000
0!
0%
#506245000000
1!
1%
#506250000000
0!
0%
#506255000000
1!
1%
#506260000000
0!
0%
#506265000000
1!
1%
#506270000000
0!
0%
#506275000000
1!
1%
#506280000000
0!
0%
#506285000000
1!
1%
#506290000000
0!
0%
#506295000000
1!
1%
#506300000000
0!
0%
#506305000000
1!
1%
#506310000000
0!
0%
#506315000000
1!
1%
#506320000000
0!
0%
#506325000000
1!
1%
#506330000000
0!
0%
#506335000000
1!
1%
#506340000000
0!
0%
#506345000000
1!
1%
#506350000000
0!
0%
#506355000000
1!
1%
#506360000000
0!
0%
#506365000000
1!
1%
#506370000000
0!
0%
#506375000000
1!
1%
#506380000000
0!
0%
#506385000000
1!
1%
#506390000000
0!
0%
#506395000000
1!
1%
#506400000000
0!
0%
#506405000000
1!
1%
#506410000000
0!
0%
#506415000000
1!
1%
#506420000000
0!
0%
#506425000000
1!
1%
#506430000000
0!
0%
#506435000000
1!
1%
#506440000000
0!
0%
#506445000000
1!
1%
#506450000000
0!
0%
#506455000000
1!
1%
#506460000000
0!
0%
#506465000000
1!
1%
#506470000000
0!
0%
#506475000000
1!
1%
#506480000000
0!
0%
#506485000000
1!
1%
#506490000000
0!
0%
#506495000000
1!
1%
#506500000000
0!
0%
#506505000000
1!
1%
#506510000000
0!
0%
#506515000000
1!
1%
#506520000000
0!
0%
#506525000000
1!
1%
#506530000000
0!
0%
#506535000000
1!
1%
#506540000000
0!
0%
#506545000000
1!
1%
#506550000000
0!
0%
#506555000000
1!
1%
#506560000000
0!
0%
#506565000000
1!
1%
#506570000000
0!
0%
#506575000000
1!
1%
#506580000000
0!
0%
#506585000000
1!
1%
#506590000000
0!
0%
#506595000000
1!
1%
#506600000000
0!
0%
#506605000000
1!
1%
#506610000000
0!
0%
#506615000000
1!
1%
#506620000000
0!
0%
#506625000000
1!
1%
#506630000000
0!
0%
#506635000000
1!
1%
#506640000000
0!
0%
#506645000000
1!
1%
#506650000000
0!
0%
#506655000000
1!
1%
#506660000000
0!
0%
#506665000000
1!
1%
#506670000000
0!
0%
#506675000000
1!
1%
#506680000000
0!
0%
#506685000000
1!
1%
#506690000000
0!
0%
#506695000000
1!
1%
#506700000000
0!
0%
#506705000000
1!
1%
#506710000000
0!
0%
#506715000000
1!
1%
#506720000000
0!
0%
#506725000000
1!
1%
#506730000000
0!
0%
#506735000000
1!
1%
#506740000000
0!
0%
#506745000000
1!
1%
#506750000000
0!
0%
#506755000000
1!
1%
#506760000000
0!
0%
#506765000000
1!
1%
#506770000000
0!
0%
#506775000000
1!
1%
#506780000000
0!
0%
#506785000000
1!
1%
#506790000000
0!
0%
#506795000000
1!
1%
#506800000000
0!
0%
#506805000000
1!
1%
#506810000000
0!
0%
#506815000000
1!
1%
#506820000000
0!
0%
#506825000000
1!
1%
#506830000000
0!
0%
#506835000000
1!
1%
#506840000000
0!
0%
#506845000000
1!
1%
#506850000000
0!
0%
#506855000000
1!
1%
#506860000000
0!
0%
#506865000000
1!
1%
#506870000000
0!
0%
#506875000000
1!
1%
#506880000000
0!
0%
#506885000000
1!
1%
#506890000000
0!
0%
#506895000000
1!
1%
#506900000000
0!
0%
#506905000000
1!
1%
#506910000000
0!
0%
#506915000000
1!
1%
#506920000000
0!
0%
#506925000000
1!
1%
#506930000000
0!
0%
#506935000000
1!
1%
#506940000000
0!
0%
#506945000000
1!
1%
#506950000000
0!
0%
#506955000000
1!
1%
#506960000000
0!
0%
#506965000000
1!
1%
#506970000000
0!
0%
#506975000000
1!
1%
#506980000000
0!
0%
#506985000000
1!
1%
#506990000000
0!
0%
#506995000000
1!
1%
#507000000000
0!
0%
#507005000000
1!
1%
#507010000000
0!
0%
#507015000000
1!
1%
#507020000000
0!
0%
#507025000000
1!
1%
#507030000000
0!
0%
#507035000000
1!
1%
#507040000000
0!
0%
#507045000000
1!
1%
#507050000000
0!
0%
#507055000000
1!
1%
#507060000000
0!
0%
#507065000000
1!
1%
#507070000000
0!
0%
#507075000000
1!
1%
#507080000000
0!
0%
#507085000000
1!
1%
#507090000000
0!
0%
#507095000000
1!
1%
#507100000000
0!
0%
#507105000000
1!
1%
#507110000000
0!
0%
#507115000000
1!
1%
#507120000000
0!
0%
#507125000000
1!
1%
#507130000000
0!
0%
#507135000000
1!
1%
#507140000000
0!
0%
#507145000000
1!
1%
#507150000000
0!
0%
#507155000000
1!
1%
#507160000000
0!
0%
#507165000000
1!
1%
#507170000000
0!
0%
#507175000000
1!
1%
#507180000000
0!
0%
#507185000000
1!
1%
#507190000000
0!
0%
#507195000000
1!
1%
#507200000000
0!
0%
#507205000000
1!
1%
#507210000000
0!
0%
#507215000000
1!
1%
#507220000000
0!
0%
#507225000000
1!
1%
#507230000000
0!
0%
#507235000000
1!
1%
#507240000000
0!
0%
#507245000000
1!
1%
#507250000000
0!
0%
#507255000000
1!
1%
#507260000000
0!
0%
#507265000000
1!
1%
#507270000000
0!
0%
#507275000000
1!
1%
#507280000000
0!
0%
#507285000000
1!
1%
#507290000000
0!
0%
#507295000000
1!
1%
#507300000000
0!
0%
#507305000000
1!
1%
#507310000000
0!
0%
#507315000000
1!
1%
#507320000000
0!
0%
#507325000000
1!
1%
#507330000000
0!
0%
#507335000000
1!
1%
#507340000000
0!
0%
#507345000000
1!
1%
#507350000000
0!
0%
#507355000000
1!
1%
#507360000000
0!
0%
#507365000000
1!
1%
#507370000000
0!
0%
#507375000000
1!
1%
#507380000000
0!
0%
#507385000000
1!
1%
#507390000000
0!
0%
#507395000000
1!
1%
#507400000000
0!
0%
#507405000000
1!
1%
#507410000000
0!
0%
#507415000000
1!
1%
#507420000000
0!
0%
#507425000000
1!
1%
#507430000000
0!
0%
#507435000000
1!
1%
#507440000000
0!
0%
#507445000000
1!
1%
#507450000000
0!
0%
#507455000000
1!
1%
#507460000000
0!
0%
#507465000000
1!
1%
#507470000000
0!
0%
#507475000000
1!
1%
#507480000000
0!
0%
#507485000000
1!
1%
#507490000000
0!
0%
#507495000000
1!
1%
#507500000000
0!
0%
#507505000000
1!
1%
#507510000000
0!
0%
#507515000000
1!
1%
#507520000000
0!
0%
#507525000000
1!
1%
#507530000000
0!
0%
#507535000000
1!
1%
#507540000000
0!
0%
#507545000000
1!
1%
#507550000000
0!
0%
#507555000000
1!
1%
#507560000000
0!
0%
#507565000000
1!
1%
#507570000000
0!
0%
#507575000000
1!
1%
#507580000000
0!
0%
#507585000000
1!
1%
#507590000000
0!
0%
#507595000000
1!
1%
#507600000000
0!
0%
#507605000000
1!
1%
#507610000000
0!
0%
#507615000000
1!
1%
#507620000000
0!
0%
#507625000000
1!
1%
#507630000000
0!
0%
#507635000000
1!
1%
#507640000000
0!
0%
#507645000000
1!
1%
#507650000000
0!
0%
#507655000000
1!
1%
#507660000000
0!
0%
#507665000000
1!
1%
#507670000000
0!
0%
#507675000000
1!
1%
#507680000000
0!
0%
#507685000000
1!
1%
#507690000000
0!
0%
#507695000000
1!
1%
#507700000000
0!
0%
#507705000000
1!
1%
#507710000000
0!
0%
#507715000000
1!
1%
#507720000000
0!
0%
#507725000000
1!
1%
#507730000000
0!
0%
#507735000000
1!
1%
#507740000000
0!
0%
#507745000000
1!
1%
#507750000000
0!
0%
#507755000000
1!
1%
#507760000000
0!
0%
#507765000000
1!
1%
#507770000000
0!
0%
#507775000000
1!
1%
#507780000000
0!
0%
#507785000000
1!
1%
#507790000000
0!
0%
#507795000000
1!
1%
#507800000000
0!
0%
#507805000000
1!
1%
#507810000000
0!
0%
#507815000000
1!
1%
#507820000000
0!
0%
#507825000000
1!
1%
#507830000000
0!
0%
#507835000000
1!
1%
#507840000000
0!
0%
#507845000000
1!
1%
#507850000000
0!
0%
#507855000000
1!
1%
#507860000000
0!
0%
#507865000000
1!
1%
#507870000000
0!
0%
#507875000000
1!
1%
#507880000000
0!
0%
#507885000000
1!
1%
#507890000000
0!
0%
#507895000000
1!
1%
#507900000000
0!
0%
#507905000000
1!
1%
#507910000000
0!
0%
#507915000000
1!
1%
#507920000000
0!
0%
#507925000000
1!
1%
#507930000000
0!
0%
#507935000000
1!
1%
#507940000000
0!
0%
#507945000000
1!
1%
#507950000000
0!
0%
#507955000000
1!
1%
#507960000000
0!
0%
#507965000000
1!
1%
#507970000000
0!
0%
#507975000000
1!
1%
#507980000000
0!
0%
#507985000000
1!
1%
#507990000000
0!
0%
#507995000000
1!
1%
#508000000000
0!
0%
#508005000000
1!
1%
#508010000000
0!
0%
#508015000000
1!
1%
#508020000000
0!
0%
#508025000000
1!
1%
#508030000000
0!
0%
#508035000000
1!
1%
#508040000000
0!
0%
#508045000000
1!
1%
#508050000000
0!
0%
#508055000000
1!
1%
#508060000000
0!
0%
#508065000000
1!
1%
#508070000000
0!
0%
#508075000000
1!
1%
#508080000000
0!
0%
#508085000000
1!
1%
#508090000000
0!
0%
#508095000000
1!
1%
#508100000000
0!
0%
#508105000000
1!
1%
#508110000000
0!
0%
#508115000000
1!
1%
#508120000000
0!
0%
#508125000000
1!
1%
#508130000000
0!
0%
#508135000000
1!
1%
#508140000000
0!
0%
#508145000000
1!
1%
#508150000000
0!
0%
#508155000000
1!
1%
#508160000000
0!
0%
#508165000000
1!
1%
#508170000000
0!
0%
#508175000000
1!
1%
#508180000000
0!
0%
#508185000000
1!
1%
#508190000000
0!
0%
#508195000000
1!
1%
#508200000000
0!
0%
#508205000000
1!
1%
#508210000000
0!
0%
#508215000000
1!
1%
#508220000000
0!
0%
#508225000000
1!
1%
#508230000000
0!
0%
#508235000000
1!
1%
#508240000000
0!
0%
#508245000000
1!
1%
#508250000000
0!
0%
#508255000000
1!
1%
#508260000000
0!
0%
#508265000000
1!
1%
#508270000000
0!
0%
#508275000000
1!
1%
#508280000000
0!
0%
#508285000000
1!
1%
#508290000000
0!
0%
#508295000000
1!
1%
#508300000000
0!
0%
#508305000000
1!
1%
#508310000000
0!
0%
#508315000000
1!
1%
#508320000000
0!
0%
#508325000000
1!
1%
#508330000000
0!
0%
#508335000000
1!
1%
#508340000000
0!
0%
#508345000000
1!
1%
#508350000000
0!
0%
#508355000000
1!
1%
#508360000000
0!
0%
#508365000000
1!
1%
#508370000000
0!
0%
#508375000000
1!
1%
#508380000000
0!
0%
#508385000000
1!
1%
#508390000000
0!
0%
#508395000000
1!
1%
#508400000000
0!
0%
#508405000000
1!
1%
#508410000000
0!
0%
#508415000000
1!
1%
#508420000000
0!
0%
#508425000000
1!
1%
#508430000000
0!
0%
#508435000000
1!
1%
#508440000000
0!
0%
#508445000000
1!
1%
#508450000000
0!
0%
#508455000000
1!
1%
#508460000000
0!
0%
#508465000000
1!
1%
#508470000000
0!
0%
#508475000000
1!
1%
#508480000000
0!
0%
#508485000000
1!
1%
#508490000000
0!
0%
#508495000000
1!
1%
#508500000000
0!
0%
#508505000000
1!
1%
#508510000000
0!
0%
#508515000000
1!
1%
#508520000000
0!
0%
#508525000000
1!
1%
#508530000000
0!
0%
#508535000000
1!
1%
#508540000000
0!
0%
#508545000000
1!
1%
#508550000000
0!
0%
#508555000000
1!
1%
#508560000000
0!
0%
#508565000000
1!
1%
#508570000000
0!
0%
#508575000000
1!
1%
#508580000000
0!
0%
#508585000000
1!
1%
#508590000000
0!
0%
#508595000000
1!
1%
#508600000000
0!
0%
#508605000000
1!
1%
#508610000000
0!
0%
#508615000000
1!
1%
#508620000000
0!
0%
#508625000000
1!
1%
#508630000000
0!
0%
#508635000000
1!
1%
#508640000000
0!
0%
#508645000000
1!
1%
#508650000000
0!
0%
#508655000000
1!
1%
#508660000000
0!
0%
#508665000000
1!
1%
#508670000000
0!
0%
#508675000000
1!
1%
#508680000000
0!
0%
#508685000000
1!
1%
#508690000000
0!
0%
#508695000000
1!
1%
#508700000000
0!
0%
#508705000000
1!
1%
#508710000000
0!
0%
#508715000000
1!
1%
#508720000000
0!
0%
#508725000000
1!
1%
#508730000000
0!
0%
#508735000000
1!
1%
#508740000000
0!
0%
#508745000000
1!
1%
#508750000000
0!
0%
#508755000000
1!
1%
#508760000000
0!
0%
#508765000000
1!
1%
#508770000000
0!
0%
#508775000000
1!
1%
#508780000000
0!
0%
#508785000000
1!
1%
#508790000000
0!
0%
#508795000000
1!
1%
#508800000000
0!
0%
#508805000000
1!
1%
#508810000000
0!
0%
#508815000000
1!
1%
#508820000000
0!
0%
#508825000000
1!
1%
#508830000000
0!
0%
#508835000000
1!
1%
#508840000000
0!
0%
#508845000000
1!
1%
#508850000000
0!
0%
#508855000000
1!
1%
#508860000000
0!
0%
#508865000000
1!
1%
#508870000000
0!
0%
#508875000000
1!
1%
#508880000000
0!
0%
#508885000000
1!
1%
#508890000000
0!
0%
#508895000000
1!
1%
#508900000000
0!
0%
#508905000000
1!
1%
#508910000000
0!
0%
#508915000000
1!
1%
#508920000000
0!
0%
#508925000000
1!
1%
#508930000000
0!
0%
#508935000000
1!
1%
#508940000000
0!
0%
#508945000000
1!
1%
#508950000000
0!
0%
#508955000000
1!
1%
#508960000000
0!
0%
#508965000000
1!
1%
#508970000000
0!
0%
#508975000000
1!
1%
#508980000000
0!
0%
#508985000000
1!
1%
#508990000000
0!
0%
#508995000000
1!
1%
#509000000000
0!
0%
#509005000000
1!
1%
#509010000000
0!
0%
#509015000000
1!
1%
#509020000000
0!
0%
#509025000000
1!
1%
#509030000000
0!
0%
#509035000000
1!
1%
#509040000000
0!
0%
#509045000000
1!
1%
#509050000000
0!
0%
#509055000000
1!
1%
#509060000000
0!
0%
#509065000000
1!
1%
#509070000000
0!
0%
#509075000000
1!
1%
#509080000000
0!
0%
#509085000000
1!
1%
#509090000000
0!
0%
#509095000000
1!
1%
#509100000000
0!
0%
#509105000000
1!
1%
#509110000000
0!
0%
#509115000000
1!
1%
#509120000000
0!
0%
#509125000000
1!
1%
#509130000000
0!
0%
#509135000000
1!
1%
#509140000000
0!
0%
#509145000000
1!
1%
#509150000000
0!
0%
#509155000000
1!
1%
#509160000000
0!
0%
#509165000000
1!
1%
#509170000000
0!
0%
#509175000000
1!
1%
#509180000000
0!
0%
#509185000000
1!
1%
#509190000000
0!
0%
#509195000000
1!
1%
#509200000000
0!
0%
#509205000000
1!
1%
#509210000000
0!
0%
#509215000000
1!
1%
#509220000000
0!
0%
#509225000000
1!
1%
#509230000000
0!
0%
#509235000000
1!
1%
#509240000000
0!
0%
#509245000000
1!
1%
#509250000000
0!
0%
#509255000000
1!
1%
#509260000000
0!
0%
#509265000000
1!
1%
#509270000000
0!
0%
#509275000000
1!
1%
#509280000000
0!
0%
#509285000000
1!
1%
#509290000000
0!
0%
#509295000000
1!
1%
#509300000000
0!
0%
#509305000000
1!
1%
#509310000000
0!
0%
#509315000000
1!
1%
#509320000000
0!
0%
#509325000000
1!
1%
#509330000000
0!
0%
#509335000000
1!
1%
#509340000000
0!
0%
#509345000000
1!
1%
#509350000000
0!
0%
#509355000000
1!
1%
#509360000000
0!
0%
#509365000000
1!
1%
#509370000000
0!
0%
#509375000000
1!
1%
#509380000000
0!
0%
#509385000000
1!
1%
#509390000000
0!
0%
#509395000000
1!
1%
#509400000000
0!
0%
#509405000000
1!
1%
#509410000000
0!
0%
#509415000000
1!
1%
#509420000000
0!
0%
#509425000000
1!
1%
#509430000000
0!
0%
#509435000000
1!
1%
#509440000000
0!
0%
#509445000000
1!
1%
#509450000000
0!
0%
#509455000000
1!
1%
#509460000000
0!
0%
#509465000000
1!
1%
#509470000000
0!
0%
#509475000000
1!
1%
#509480000000
0!
0%
#509485000000
1!
1%
#509490000000
0!
0%
#509495000000
1!
1%
#509500000000
0!
0%
#509505000000
1!
1%
#509510000000
0!
0%
#509515000000
1!
1%
#509520000000
0!
0%
#509525000000
1!
1%
#509530000000
0!
0%
#509535000000
1!
1%
#509540000000
0!
0%
#509545000000
1!
1%
#509550000000
0!
0%
#509555000000
1!
1%
#509560000000
0!
0%
#509565000000
1!
1%
#509570000000
0!
0%
#509575000000
1!
1%
#509580000000
0!
0%
#509585000000
1!
1%
#509590000000
0!
0%
#509595000000
1!
1%
#509600000000
0!
0%
#509605000000
1!
1%
#509610000000
0!
0%
#509615000000
1!
1%
#509620000000
0!
0%
#509625000000
1!
1%
#509630000000
0!
0%
#509635000000
1!
1%
#509640000000
0!
0%
#509645000000
1!
1%
#509650000000
0!
0%
#509655000000
1!
1%
#509660000000
0!
0%
#509665000000
1!
1%
#509670000000
0!
0%
#509675000000
1!
1%
#509680000000
0!
0%
#509685000000
1!
1%
#509690000000
0!
0%
#509695000000
1!
1%
#509700000000
0!
0%
#509705000000
1!
1%
#509710000000
0!
0%
#509715000000
1!
1%
#509720000000
0!
0%
#509725000000
1!
1%
#509730000000
0!
0%
#509735000000
1!
1%
#509740000000
0!
0%
#509745000000
1!
1%
#509750000000
0!
0%
#509755000000
1!
1%
#509760000000
0!
0%
#509765000000
1!
1%
#509770000000
0!
0%
#509775000000
1!
1%
#509780000000
0!
0%
#509785000000
1!
1%
#509790000000
0!
0%
#509795000000
1!
1%
#509800000000
0!
0%
#509805000000
1!
1%
#509810000000
0!
0%
#509815000000
1!
1%
#509820000000
0!
0%
#509825000000
1!
1%
#509830000000
0!
0%
#509835000000
1!
1%
#509840000000
0!
0%
#509845000000
1!
1%
#509850000000
0!
0%
#509855000000
1!
1%
#509860000000
0!
0%
#509865000000
1!
1%
#509870000000
0!
0%
#509875000000
1!
1%
#509880000000
0!
0%
#509885000000
1!
1%
#509890000000
0!
0%
#509895000000
1!
1%
#509900000000
0!
0%
#509905000000
1!
1%
#509910000000
0!
0%
#509915000000
1!
1%
#509920000000
0!
0%
#509925000000
1!
1%
#509930000000
0!
0%
#509935000000
1!
1%
#509940000000
0!
0%
#509945000000
1!
1%
#509950000000
0!
0%
#509955000000
1!
1%
#509960000000
0!
0%
#509965000000
1!
1%
#509970000000
0!
0%
#509975000000
1!
1%
#509980000000
0!
0%
#509985000000
1!
1%
#509990000000
0!
0%
#509995000000
1!
1%
#510000000000
0!
0%
#510005000000
1!
1%
#510010000000
0!
0%
#510015000000
1!
1%
#510020000000
0!
0%
#510025000000
1!
1%
#510030000000
0!
0%
#510035000000
1!
1%
#510040000000
0!
0%
#510045000000
1!
1%
#510050000000
0!
0%
#510055000000
1!
1%
#510060000000
0!
0%
#510065000000
1!
1%
#510070000000
0!
0%
#510075000000
1!
1%
#510080000000
0!
0%
#510085000000
1!
1%
#510090000000
0!
0%
#510095000000
1!
1%
#510100000000
0!
0%
#510105000000
1!
1%
#510110000000
0!
0%
#510115000000
1!
1%
#510120000000
0!
0%
#510125000000
1!
1%
#510130000000
0!
0%
#510135000000
1!
1%
#510140000000
0!
0%
#510145000000
1!
1%
#510150000000
0!
0%
#510155000000
1!
1%
#510160000000
0!
0%
#510165000000
1!
1%
#510170000000
0!
0%
#510175000000
1!
1%
#510180000000
0!
0%
#510185000000
1!
1%
#510190000000
0!
0%
#510195000000
1!
1%
#510200000000
0!
0%
#510205000000
1!
1%
#510210000000
0!
0%
#510215000000
1!
1%
#510220000000
0!
0%
#510225000000
1!
1%
#510230000000
0!
0%
#510235000000
1!
1%
#510240000000
0!
0%
#510245000000
1!
1%
#510250000000
0!
0%
#510255000000
1!
1%
#510260000000
0!
0%
#510265000000
1!
1%
#510270000000
0!
0%
#510275000000
1!
1%
#510280000000
0!
0%
#510285000000
1!
1%
#510290000000
0!
0%
#510295000000
1!
1%
#510300000000
0!
0%
#510305000000
1!
1%
#510310000000
0!
0%
#510315000000
1!
1%
#510320000000
0!
0%
#510325000000
1!
1%
#510330000000
0!
0%
#510335000000
1!
1%
#510340000000
0!
0%
#510345000000
1!
1%
#510350000000
0!
0%
#510355000000
1!
1%
#510360000000
0!
0%
#510365000000
1!
1%
#510370000000
0!
0%
#510375000000
1!
1%
#510380000000
0!
0%
#510385000000
1!
1%
#510390000000
0!
0%
#510395000000
1!
1%
#510400000000
0!
0%
#510405000000
1!
1%
#510410000000
0!
0%
#510415000000
1!
1%
#510420000000
0!
0%
#510425000000
1!
1%
#510430000000
0!
0%
#510435000000
1!
1%
#510440000000
0!
0%
#510445000000
1!
1%
#510450000000
0!
0%
#510455000000
1!
1%
#510460000000
0!
0%
#510465000000
1!
1%
#510470000000
0!
0%
#510475000000
1!
1%
#510480000000
0!
0%
#510485000000
1!
1%
#510490000000
0!
0%
#510495000000
1!
1%
#510500000000
0!
0%
#510505000000
1!
1%
#510510000000
0!
0%
#510515000000
1!
1%
#510520000000
0!
0%
#510525000000
1!
1%
#510530000000
0!
0%
#510535000000
1!
1%
#510540000000
0!
0%
#510545000000
1!
1%
#510550000000
0!
0%
#510555000000
1!
1%
#510560000000
0!
0%
#510565000000
1!
1%
#510570000000
0!
0%
#510575000000
1!
1%
#510580000000
0!
0%
#510585000000
1!
1%
#510590000000
0!
0%
#510595000000
1!
1%
#510600000000
0!
0%
#510605000000
1!
1%
#510610000000
0!
0%
#510615000000
1!
1%
#510620000000
0!
0%
#510625000000
1!
1%
#510630000000
0!
0%
#510635000000
1!
1%
#510640000000
0!
0%
#510645000000
1!
1%
#510650000000
0!
0%
#510655000000
1!
1%
#510660000000
0!
0%
#510665000000
1!
1%
#510670000000
0!
0%
#510675000000
1!
1%
#510680000000
0!
0%
#510685000000
1!
1%
#510690000000
0!
0%
#510695000000
1!
1%
#510700000000
0!
0%
#510705000000
1!
1%
#510710000000
0!
0%
#510715000000
1!
1%
#510720000000
0!
0%
#510725000000
1!
1%
#510730000000
0!
0%
#510735000000
1!
1%
#510740000000
0!
0%
#510745000000
1!
1%
#510750000000
0!
0%
#510755000000
1!
1%
#510760000000
0!
0%
#510765000000
1!
1%
#510770000000
0!
0%
#510775000000
1!
1%
#510780000000
0!
0%
#510785000000
1!
1%
#510790000000
0!
0%
#510795000000
1!
1%
#510800000000
0!
0%
#510805000000
1!
1%
#510810000000
0!
0%
#510815000000
1!
1%
#510820000000
0!
0%
#510825000000
1!
1%
#510830000000
0!
0%
#510835000000
1!
1%
#510840000000
0!
0%
#510845000000
1!
1%
#510850000000
0!
0%
#510855000000
1!
1%
#510860000000
0!
0%
#510865000000
1!
1%
#510870000000
0!
0%
#510875000000
1!
1%
#510880000000
0!
0%
#510885000000
1!
1%
#510890000000
0!
0%
#510895000000
1!
1%
#510900000000
0!
0%
#510905000000
1!
1%
#510910000000
0!
0%
#510915000000
1!
1%
#510920000000
0!
0%
#510925000000
1!
1%
#510930000000
0!
0%
#510935000000
1!
1%
#510940000000
0!
0%
#510945000000
1!
1%
#510950000000
0!
0%
#510955000000
1!
1%
#510960000000
0!
0%
#510965000000
1!
1%
#510970000000
0!
0%
#510975000000
1!
1%
#510980000000
0!
0%
#510985000000
1!
1%
#510990000000
0!
0%
#510995000000
1!
1%
#511000000000
0!
0%
#511005000000
1!
1%
#511010000000
0!
0%
#511015000000
1!
1%
#511020000000
0!
0%
#511025000000
1!
1%
#511030000000
0!
0%
#511035000000
1!
1%
#511040000000
0!
0%
#511045000000
1!
1%
#511050000000
0!
0%
#511055000000
1!
1%
#511060000000
0!
0%
#511065000000
1!
1%
#511070000000
0!
0%
#511075000000
1!
1%
#511080000000
0!
0%
#511085000000
1!
1%
#511090000000
0!
0%
#511095000000
1!
1%
#511100000000
0!
0%
#511105000000
1!
1%
#511110000000
0!
0%
#511115000000
1!
1%
#511120000000
0!
0%
#511125000000
1!
1%
#511130000000
0!
0%
#511135000000
1!
1%
#511140000000
0!
0%
#511145000000
1!
1%
#511150000000
0!
0%
#511155000000
1!
1%
#511160000000
0!
0%
#511165000000
1!
1%
#511170000000
0!
0%
#511175000000
1!
1%
#511180000000
0!
0%
#511185000000
1!
1%
#511190000000
0!
0%
#511195000000
1!
1%
#511200000000
0!
0%
#511205000000
1!
1%
#511210000000
0!
0%
#511215000000
1!
1%
#511220000000
0!
0%
#511225000000
1!
1%
#511230000000
0!
0%
#511235000000
1!
1%
#511240000000
0!
0%
#511245000000
1!
1%
#511250000000
0!
0%
#511255000000
1!
1%
#511260000000
0!
0%
#511265000000
1!
1%
#511270000000
0!
0%
#511275000000
1!
1%
#511280000000
0!
0%
#511285000000
1!
1%
#511290000000
0!
0%
#511295000000
1!
1%
#511300000000
0!
0%
#511305000000
1!
1%
#511310000000
0!
0%
#511315000000
1!
1%
#511320000000
0!
0%
#511325000000
1!
1%
#511330000000
0!
0%
#511335000000
1!
1%
#511340000000
0!
0%
#511345000000
1!
1%
#511350000000
0!
0%
#511355000000
1!
1%
#511360000000
0!
0%
#511365000000
1!
1%
#511370000000
0!
0%
#511375000000
1!
1%
#511380000000
0!
0%
#511385000000
1!
1%
#511390000000
0!
0%
#511395000000
1!
1%
#511400000000
0!
0%
#511405000000
1!
1%
#511410000000
0!
0%
#511415000000
1!
1%
#511420000000
0!
0%
#511425000000
1!
1%
#511430000000
0!
0%
#511435000000
1!
1%
#511440000000
0!
0%
#511445000000
1!
1%
#511450000000
0!
0%
#511455000000
1!
1%
#511460000000
0!
0%
#511465000000
1!
1%
#511470000000
0!
0%
#511475000000
1!
1%
#511480000000
0!
0%
#511485000000
1!
1%
#511490000000
0!
0%
#511495000000
1!
1%
#511500000000
0!
0%
#511505000000
1!
1%
#511510000000
0!
0%
#511515000000
1!
1%
#511520000000
0!
0%
#511525000000
1!
1%
#511530000000
0!
0%
#511535000000
1!
1%
#511540000000
0!
0%
#511545000000
1!
1%
#511550000000
0!
0%
#511555000000
1!
1%
#511560000000
0!
0%
#511565000000
1!
1%
#511570000000
0!
0%
#511575000000
1!
1%
#511580000000
0!
0%
#511585000000
1!
1%
#511590000000
0!
0%
#511595000000
1!
1%
#511600000000
0!
0%
#511605000000
1!
1%
#511610000000
0!
0%
#511615000000
1!
1%
#511620000000
0!
0%
#511625000000
1!
1%
#511630000000
0!
0%
#511635000000
1!
1%
#511640000000
0!
0%
#511645000000
1!
1%
#511650000000
0!
0%
#511655000000
1!
1%
#511660000000
0!
0%
#511665000000
1!
1%
#511670000000
0!
0%
#511675000000
1!
1%
#511680000000
0!
0%
#511685000000
1!
1%
#511690000000
0!
0%
#511695000000
1!
1%
#511700000000
0!
0%
#511705000000
1!
1%
#511710000000
0!
0%
#511715000000
1!
1%
#511720000000
0!
0%
#511725000000
1!
1%
#511730000000
0!
0%
#511735000000
1!
1%
#511740000000
0!
0%
#511745000000
1!
1%
#511750000000
0!
0%
#511755000000
1!
1%
#511760000000
0!
0%
#511765000000
1!
1%
#511770000000
0!
0%
#511775000000
1!
1%
#511780000000
0!
0%
#511785000000
1!
1%
#511790000000
0!
0%
#511795000000
1!
1%
#511800000000
0!
0%
#511805000000
1!
1%
#511810000000
0!
0%
#511815000000
1!
1%
#511820000000
0!
0%
#511825000000
1!
1%
#511830000000
0!
0%
#511835000000
1!
1%
#511840000000
0!
0%
#511845000000
1!
1%
#511850000000
0!
0%
#511855000000
1!
1%
#511860000000
0!
0%
#511865000000
1!
1%
#511870000000
0!
0%
#511875000000
1!
1%
#511880000000
0!
0%
#511885000000
1!
1%
#511890000000
0!
0%
#511895000000
1!
1%
#511900000000
0!
0%
#511905000000
1!
1%
#511910000000
0!
0%
#511915000000
1!
1%
#511920000000
0!
0%
#511925000000
1!
1%
#511930000000
0!
0%
#511935000000
1!
1%
#511940000000
0!
0%
#511945000000
1!
1%
#511950000000
0!
0%
#511955000000
1!
1%
#511960000000
0!
0%
#511965000000
1!
1%
#511970000000
0!
0%
#511975000000
1!
1%
#511980000000
0!
0%
#511985000000
1!
1%
#511990000000
0!
0%
#511995000000
1!
1%
#512000000000
0!
0%
#512005000000
1!
1%
#512010000000
0!
0%
#512015000000
1!
1%
#512020000000
0!
0%
#512025000000
1!
1%
#512030000000
0!
0%
#512035000000
1!
1%
#512040000000
0!
0%
#512045000000
1!
1%
#512050000000
0!
0%
#512055000000
1!
1%
#512060000000
0!
0%
#512065000000
1!
1%
#512070000000
0!
0%
#512075000000
1!
1%
#512080000000
0!
0%
#512085000000
1!
1%
#512090000000
0!
0%
#512095000000
1!
1%
#512100000000
0!
0%
#512105000000
1!
1%
#512110000000
0!
0%
#512115000000
1!
1%
#512120000000
0!
0%
#512125000000
1!
1%
#512130000000
0!
0%
#512135000000
1!
1%
#512140000000
0!
0%
#512145000000
1!
1%
#512150000000
0!
0%
#512155000000
1!
1%
#512160000000
0!
0%
#512165000000
1!
1%
#512170000000
0!
0%
#512175000000
1!
1%
#512180000000
0!
0%
#512185000000
1!
1%
#512190000000
0!
0%
#512195000000
1!
1%
#512200000000
0!
0%
#512205000000
1!
1%
#512210000000
0!
0%
#512215000000
1!
1%
#512220000000
0!
0%
#512225000000
1!
1%
#512230000000
0!
0%
#512235000000
1!
1%
#512240000000
0!
0%
#512245000000
1!
1%
#512250000000
0!
0%
#512255000000
1!
1%
#512260000000
0!
0%
#512265000000
1!
1%
#512270000000
0!
0%
#512275000000
1!
1%
#512280000000
0!
0%
#512285000000
1!
1%
#512290000000
0!
0%
#512295000000
1!
1%
#512300000000
0!
0%
#512305000000
1!
1%
#512310000000
0!
0%
#512315000000
1!
1%
#512320000000
0!
0%
#512325000000
1!
1%
#512330000000
0!
0%
#512335000000
1!
1%
#512340000000
0!
0%
#512345000000
1!
1%
#512350000000
0!
0%
#512355000000
1!
1%
#512360000000
0!
0%
#512365000000
1!
1%
#512370000000
0!
0%
#512375000000
1!
1%
#512380000000
0!
0%
#512385000000
1!
1%
#512390000000
0!
0%
#512395000000
1!
1%
#512400000000
0!
0%
#512405000000
1!
1%
#512410000000
0!
0%
#512415000000
1!
1%
#512420000000
0!
0%
#512425000000
1!
1%
#512430000000
0!
0%
#512435000000
1!
1%
#512440000000
0!
0%
#512445000000
1!
1%
#512450000000
0!
0%
#512455000000
1!
1%
#512460000000
0!
0%
#512465000000
1!
1%
#512470000000
0!
0%
#512475000000
1!
1%
#512480000000
0!
0%
#512485000000
1!
1%
#512490000000
0!
0%
#512495000000
1!
1%
#512500000000
0!
0%
#512505000000
1!
1%
#512510000000
0!
0%
#512515000000
1!
1%
#512520000000
0!
0%
#512525000000
1!
1%
#512530000000
0!
0%
#512535000000
1!
1%
#512540000000
0!
0%
#512545000000
1!
1%
#512550000000
0!
0%
#512555000000
1!
1%
#512560000000
0!
0%
#512565000000
1!
1%
#512570000000
0!
0%
#512575000000
1!
1%
#512580000000
0!
0%
#512585000000
1!
1%
#512590000000
0!
0%
#512595000000
1!
1%
#512600000000
0!
0%
#512605000000
1!
1%
#512610000000
0!
0%
#512615000000
1!
1%
#512620000000
0!
0%
#512625000000
1!
1%
#512630000000
0!
0%
#512635000000
1!
1%
#512640000000
0!
0%
#512645000000
1!
1%
#512650000000
0!
0%
#512655000000
1!
1%
#512660000000
0!
0%
#512665000000
1!
1%
#512670000000
0!
0%
#512675000000
1!
1%
#512680000000
0!
0%
#512685000000
1!
1%
#512690000000
0!
0%
#512695000000
1!
1%
#512700000000
0!
0%
#512705000000
1!
1%
#512710000000
0!
0%
#512715000000
1!
1%
#512720000000
0!
0%
#512725000000
1!
1%
#512730000000
0!
0%
#512735000000
1!
1%
#512740000000
0!
0%
#512745000000
1!
1%
#512750000000
0!
0%
#512755000000
1!
1%
#512760000000
0!
0%
#512765000000
1!
1%
#512770000000
0!
0%
#512775000000
1!
1%
#512780000000
0!
0%
#512785000000
1!
1%
#512790000000
0!
0%
#512795000000
1!
1%
#512800000000
0!
0%
#512805000000
1!
1%
#512810000000
0!
0%
#512815000000
1!
1%
#512820000000
0!
0%
#512825000000
1!
1%
#512830000000
0!
0%
#512835000000
1!
1%
#512840000000
0!
0%
#512845000000
1!
1%
#512850000000
0!
0%
#512855000000
1!
1%
#512860000000
0!
0%
#512865000000
1!
1%
#512870000000
0!
0%
#512875000000
1!
1%
#512880000000
0!
0%
#512885000000
1!
1%
#512890000000
0!
0%
#512895000000
1!
1%
#512900000000
0!
0%
#512905000000
1!
1%
#512910000000
0!
0%
#512915000000
1!
1%
#512920000000
0!
0%
#512925000000
1!
1%
#512930000000
0!
0%
#512935000000
1!
1%
#512940000000
0!
0%
#512945000000
1!
1%
#512950000000
0!
0%
#512955000000
1!
1%
#512960000000
0!
0%
#512965000000
1!
1%
#512970000000
0!
0%
#512975000000
1!
1%
#512980000000
0!
0%
#512985000000
1!
1%
#512990000000
0!
0%
#512995000000
1!
1%
#513000000000
0!
0%
#513005000000
1!
1%
#513010000000
0!
0%
#513015000000
1!
1%
#513020000000
0!
0%
#513025000000
1!
1%
#513030000000
0!
0%
#513035000000
1!
1%
#513040000000
0!
0%
#513045000000
1!
1%
#513050000000
0!
0%
#513055000000
1!
1%
#513060000000
0!
0%
#513065000000
1!
1%
#513070000000
0!
0%
#513075000000
1!
1%
#513080000000
0!
0%
#513085000000
1!
1%
#513090000000
0!
0%
#513095000000
1!
1%
#513100000000
0!
0%
#513105000000
1!
1%
#513110000000
0!
0%
#513115000000
1!
1%
#513120000000
0!
0%
#513125000000
1!
1%
#513130000000
0!
0%
#513135000000
1!
1%
#513140000000
0!
0%
#513145000000
1!
1%
#513150000000
0!
0%
#513155000000
1!
1%
#513160000000
0!
0%
#513165000000
1!
1%
#513170000000
0!
0%
#513175000000
1!
1%
#513180000000
0!
0%
#513185000000
1!
1%
#513190000000
0!
0%
#513195000000
1!
1%
#513200000000
0!
0%
#513205000000
1!
1%
#513210000000
0!
0%
#513215000000
1!
1%
#513220000000
0!
0%
#513225000000
1!
1%
#513230000000
0!
0%
#513235000000
1!
1%
#513240000000
0!
0%
#513245000000
1!
1%
#513250000000
0!
0%
#513255000000
1!
1%
#513260000000
0!
0%
#513265000000
1!
1%
#513270000000
0!
0%
#513275000000
1!
1%
#513280000000
0!
0%
#513285000000
1!
1%
#513290000000
0!
0%
#513295000000
1!
1%
#513300000000
0!
0%
#513305000000
1!
1%
#513310000000
0!
0%
#513315000000
1!
1%
#513320000000
0!
0%
#513325000000
1!
1%
#513330000000
0!
0%
#513335000000
1!
1%
#513340000000
0!
0%
#513345000000
1!
1%
#513350000000
0!
0%
#513355000000
1!
1%
#513360000000
0!
0%
#513365000000
1!
1%
#513370000000
0!
0%
#513375000000
1!
1%
#513380000000
0!
0%
#513385000000
1!
1%
#513390000000
0!
0%
#513395000000
1!
1%
#513400000000
0!
0%
#513405000000
1!
1%
#513410000000
0!
0%
#513415000000
1!
1%
#513420000000
0!
0%
#513425000000
1!
1%
#513430000000
0!
0%
#513435000000
1!
1%
#513440000000
0!
0%
#513445000000
1!
1%
#513450000000
0!
0%
#513455000000
1!
1%
#513460000000
0!
0%
#513465000000
1!
1%
#513470000000
0!
0%
#513475000000
1!
1%
#513480000000
0!
0%
#513485000000
1!
1%
#513490000000
0!
0%
#513495000000
1!
1%
#513500000000
0!
0%
#513505000000
1!
1%
#513510000000
0!
0%
#513515000000
1!
1%
#513520000000
0!
0%
#513525000000
1!
1%
#513530000000
0!
0%
#513535000000
1!
1%
#513540000000
0!
0%
#513545000000
1!
1%
#513550000000
0!
0%
#513555000000
1!
1%
#513560000000
0!
0%
#513565000000
1!
1%
#513570000000
0!
0%
#513575000000
1!
1%
#513580000000
0!
0%
#513585000000
1!
1%
#513590000000
0!
0%
#513595000000
1!
1%
#513600000000
0!
0%
#513605000000
1!
1%
#513610000000
0!
0%
#513615000000
1!
1%
#513620000000
0!
0%
#513625000000
1!
1%
#513630000000
0!
0%
#513635000000
1!
1%
#513640000000
0!
0%
#513645000000
1!
1%
#513650000000
0!
0%
#513655000000
1!
1%
#513660000000
0!
0%
#513665000000
1!
1%
#513670000000
0!
0%
#513675000000
1!
1%
#513680000000
0!
0%
#513685000000
1!
1%
#513690000000
0!
0%
#513695000000
1!
1%
#513700000000
0!
0%
#513705000000
1!
1%
#513710000000
0!
0%
#513715000000
1!
1%
#513720000000
0!
0%
#513725000000
1!
1%
#513730000000
0!
0%
#513735000000
1!
1%
#513740000000
0!
0%
#513745000000
1!
1%
#513750000000
0!
0%
#513755000000
1!
1%
#513760000000
0!
0%
#513765000000
1!
1%
#513770000000
0!
0%
#513775000000
1!
1%
#513780000000
0!
0%
#513785000000
1!
1%
#513790000000
0!
0%
#513795000000
1!
1%
#513800000000
0!
0%
#513805000000
1!
1%
#513810000000
0!
0%
#513815000000
1!
1%
#513820000000
0!
0%
#513825000000
1!
1%
#513830000000
0!
0%
#513835000000
1!
1%
#513840000000
0!
0%
#513845000000
1!
1%
#513850000000
0!
0%
#513855000000
1!
1%
#513860000000
0!
0%
#513865000000
1!
1%
#513870000000
0!
0%
#513875000000
1!
1%
#513880000000
0!
0%
#513885000000
1!
1%
#513890000000
0!
0%
#513895000000
1!
1%
#513900000000
0!
0%
#513905000000
1!
1%
#513910000000
0!
0%
#513915000000
1!
1%
#513920000000
0!
0%
#513925000000
1!
1%
#513930000000
0!
0%
#513935000000
1!
1%
#513940000000
0!
0%
#513945000000
1!
1%
#513950000000
0!
0%
#513955000000
1!
1%
#513960000000
0!
0%
#513965000000
1!
1%
#513970000000
0!
0%
#513975000000
1!
1%
#513980000000
0!
0%
#513985000000
1!
1%
#513990000000
0!
0%
#513995000000
1!
1%
#514000000000
0!
0%
#514005000000
1!
1%
#514010000000
0!
0%
#514015000000
1!
1%
#514020000000
0!
0%
#514025000000
1!
1%
#514030000000
0!
0%
#514035000000
1!
1%
#514040000000
0!
0%
#514045000000
1!
1%
#514050000000
0!
0%
#514055000000
1!
1%
#514060000000
0!
0%
#514065000000
1!
1%
#514070000000
0!
0%
#514075000000
1!
1%
#514080000000
0!
0%
#514085000000
1!
1%
#514090000000
0!
0%
#514095000000
1!
1%
#514100000000
0!
0%
#514105000000
1!
1%
#514110000000
0!
0%
#514115000000
1!
1%
#514120000000
0!
0%
#514125000000
1!
1%
#514130000000
0!
0%
#514135000000
1!
1%
#514140000000
0!
0%
#514145000000
1!
1%
#514150000000
0!
0%
#514155000000
1!
1%
#514160000000
0!
0%
#514165000000
1!
1%
#514170000000
0!
0%
#514175000000
1!
1%
#514180000000
0!
0%
#514185000000
1!
1%
#514190000000
0!
0%
#514195000000
1!
1%
#514200000000
0!
0%
#514205000000
1!
1%
#514210000000
0!
0%
#514215000000
1!
1%
#514220000000
0!
0%
#514225000000
1!
1%
#514230000000
0!
0%
#514235000000
1!
1%
#514240000000
0!
0%
#514245000000
1!
1%
#514250000000
0!
0%
#514255000000
1!
1%
#514260000000
0!
0%
#514265000000
1!
1%
#514270000000
0!
0%
#514275000000
1!
1%
#514280000000
0!
0%
#514285000000
1!
1%
#514290000000
0!
0%
#514295000000
1!
1%
#514300000000
0!
0%
#514305000000
1!
1%
#514310000000
0!
0%
#514315000000
1!
1%
#514320000000
0!
0%
#514325000000
1!
1%
#514330000000
0!
0%
#514335000000
1!
1%
#514340000000
0!
0%
#514345000000
1!
1%
#514350000000
0!
0%
#514355000000
1!
1%
#514360000000
0!
0%
#514365000000
1!
1%
#514370000000
0!
0%
#514375000000
1!
1%
#514380000000
0!
0%
#514385000000
1!
1%
#514390000000
0!
0%
#514395000000
1!
1%
#514400000000
0!
0%
#514405000000
1!
1%
#514410000000
0!
0%
#514415000000
1!
1%
#514420000000
0!
0%
#514425000000
1!
1%
#514430000000
0!
0%
#514435000000
1!
1%
#514440000000
0!
0%
#514445000000
1!
1%
#514450000000
0!
0%
#514455000000
1!
1%
#514460000000
0!
0%
#514465000000
1!
1%
#514470000000
0!
0%
#514475000000
1!
1%
#514480000000
0!
0%
#514485000000
1!
1%
#514490000000
0!
0%
#514495000000
1!
1%
#514500000000
0!
0%
#514505000000
1!
1%
#514510000000
0!
0%
#514515000000
1!
1%
#514520000000
0!
0%
#514525000000
1!
1%
#514530000000
0!
0%
#514535000000
1!
1%
#514540000000
0!
0%
#514545000000
1!
1%
#514550000000
0!
0%
#514555000000
1!
1%
#514560000000
0!
0%
#514565000000
1!
1%
#514570000000
0!
0%
#514575000000
1!
1%
#514580000000
0!
0%
#514585000000
1!
1%
#514590000000
0!
0%
#514595000000
1!
1%
#514600000000
0!
0%
#514605000000
1!
1%
#514610000000
0!
0%
#514615000000
1!
1%
#514620000000
0!
0%
#514625000000
1!
1%
#514630000000
0!
0%
#514635000000
1!
1%
#514640000000
0!
0%
#514645000000
1!
1%
#514650000000
0!
0%
#514655000000
1!
1%
#514660000000
0!
0%
#514665000000
1!
1%
#514670000000
0!
0%
#514675000000
1!
1%
#514680000000
0!
0%
#514685000000
1!
1%
#514690000000
0!
0%
#514695000000
1!
1%
#514700000000
0!
0%
#514705000000
1!
1%
#514710000000
0!
0%
#514715000000
1!
1%
#514720000000
0!
0%
#514725000000
1!
1%
#514730000000
0!
0%
#514735000000
1!
1%
#514740000000
0!
0%
#514745000000
1!
1%
#514750000000
0!
0%
#514755000000
1!
1%
#514760000000
0!
0%
#514765000000
1!
1%
#514770000000
0!
0%
#514775000000
1!
1%
#514780000000
0!
0%
#514785000000
1!
1%
#514790000000
0!
0%
#514795000000
1!
1%
#514800000000
0!
0%
#514805000000
1!
1%
#514810000000
0!
0%
#514815000000
1!
1%
#514820000000
0!
0%
#514825000000
1!
1%
#514830000000
0!
0%
#514835000000
1!
1%
#514840000000
0!
0%
#514845000000
1!
1%
#514850000000
0!
0%
#514855000000
1!
1%
#514860000000
0!
0%
#514865000000
1!
1%
#514870000000
0!
0%
#514875000000
1!
1%
#514880000000
0!
0%
#514885000000
1!
1%
#514890000000
0!
0%
#514895000000
1!
1%
#514900000000
0!
0%
#514905000000
1!
1%
#514910000000
0!
0%
#514915000000
1!
1%
#514920000000
0!
0%
#514925000000
1!
1%
#514930000000
0!
0%
#514935000000
1!
1%
#514940000000
0!
0%
#514945000000
1!
1%
#514950000000
0!
0%
#514955000000
1!
1%
#514960000000
0!
0%
#514965000000
1!
1%
#514970000000
0!
0%
#514975000000
1!
1%
#514980000000
0!
0%
#514985000000
1!
1%
#514990000000
0!
0%
#514995000000
1!
1%
#515000000000
0!
0%
#515005000000
1!
1%
#515010000000
0!
0%
#515015000000
1!
1%
#515020000000
0!
0%
#515025000000
1!
1%
#515030000000
0!
0%
#515035000000
1!
1%
#515040000000
0!
0%
#515045000000
1!
1%
#515050000000
0!
0%
#515055000000
1!
1%
#515060000000
0!
0%
#515065000000
1!
1%
#515070000000
0!
0%
#515075000000
1!
1%
#515080000000
0!
0%
#515085000000
1!
1%
#515090000000
0!
0%
#515095000000
1!
1%
#515100000000
0!
0%
#515105000000
1!
1%
#515110000000
0!
0%
#515115000000
1!
1%
#515120000000
0!
0%
#515125000000
1!
1%
#515130000000
0!
0%
#515135000000
1!
1%
#515140000000
0!
0%
#515145000000
1!
1%
#515150000000
0!
0%
#515155000000
1!
1%
#515160000000
0!
0%
#515165000000
1!
1%
#515170000000
0!
0%
#515175000000
1!
1%
#515180000000
0!
0%
#515185000000
1!
1%
#515190000000
0!
0%
#515195000000
1!
1%
#515200000000
0!
0%
#515205000000
1!
1%
#515210000000
0!
0%
#515215000000
1!
1%
#515220000000
0!
0%
#515225000000
1!
1%
#515230000000
0!
0%
#515235000000
1!
1%
#515240000000
0!
0%
#515245000000
1!
1%
#515250000000
0!
0%
#515255000000
1!
1%
#515260000000
0!
0%
#515265000000
1!
1%
#515270000000
0!
0%
#515275000000
1!
1%
#515280000000
0!
0%
#515285000000
1!
1%
#515290000000
0!
0%
#515295000000
1!
1%
#515300000000
0!
0%
#515305000000
1!
1%
#515310000000
0!
0%
#515315000000
1!
1%
#515320000000
0!
0%
#515325000000
1!
1%
#515330000000
0!
0%
#515335000000
1!
1%
#515340000000
0!
0%
#515345000000
1!
1%
#515350000000
0!
0%
#515355000000
1!
1%
#515360000000
0!
0%
#515365000000
1!
1%
#515370000000
0!
0%
#515375000000
1!
1%
#515380000000
0!
0%
#515385000000
1!
1%
#515390000000
0!
0%
#515395000000
1!
1%
#515400000000
0!
0%
#515405000000
1!
1%
#515410000000
0!
0%
#515415000000
1!
1%
#515420000000
0!
0%
#515425000000
1!
1%
#515430000000
0!
0%
#515435000000
1!
1%
#515440000000
0!
0%
#515445000000
1!
1%
#515450000000
0!
0%
#515455000000
1!
1%
#515460000000
0!
0%
#515465000000
1!
1%
#515470000000
0!
0%
#515475000000
1!
1%
#515480000000
0!
0%
#515485000000
1!
1%
#515490000000
0!
0%
#515495000000
1!
1%
#515500000000
0!
0%
#515505000000
1!
1%
#515510000000
0!
0%
#515515000000
1!
1%
#515520000000
0!
0%
#515525000000
1!
1%
#515530000000
0!
0%
#515535000000
1!
1%
#515540000000
0!
0%
#515545000000
1!
1%
#515550000000
0!
0%
#515555000000
1!
1%
#515560000000
0!
0%
#515565000000
1!
1%
#515570000000
0!
0%
#515575000000
1!
1%
#515580000000
0!
0%
#515585000000
1!
1%
#515590000000
0!
0%
#515595000000
1!
1%
#515600000000
0!
0%
#515605000000
1!
1%
#515610000000
0!
0%
#515615000000
1!
1%
#515620000000
0!
0%
#515625000000
1!
1%
#515630000000
0!
0%
#515635000000
1!
1%
#515640000000
0!
0%
#515645000000
1!
1%
#515650000000
0!
0%
#515655000000
1!
1%
#515660000000
0!
0%
#515665000000
1!
1%
#515670000000
0!
0%
#515675000000
1!
1%
#515680000000
0!
0%
#515685000000
1!
1%
#515690000000
0!
0%
#515695000000
1!
1%
#515700000000
0!
0%
#515705000000
1!
1%
#515710000000
0!
0%
#515715000000
1!
1%
#515720000000
0!
0%
#515725000000
1!
1%
#515730000000
0!
0%
#515735000000
1!
1%
#515740000000
0!
0%
#515745000000
1!
1%
#515750000000
0!
0%
#515755000000
1!
1%
#515760000000
0!
0%
#515765000000
1!
1%
#515770000000
0!
0%
#515775000000
1!
1%
#515780000000
0!
0%
#515785000000
1!
1%
#515790000000
0!
0%
#515795000000
1!
1%
#515800000000
0!
0%
#515805000000
1!
1%
#515810000000
0!
0%
#515815000000
1!
1%
#515820000000
0!
0%
#515825000000
1!
1%
#515830000000
0!
0%
#515835000000
1!
1%
#515840000000
0!
0%
#515845000000
1!
1%
#515850000000
0!
0%
#515855000000
1!
1%
#515860000000
0!
0%
#515865000000
1!
1%
#515870000000
0!
0%
#515875000000
1!
1%
#515880000000
0!
0%
#515885000000
1!
1%
#515890000000
0!
0%
#515895000000
1!
1%
#515900000000
0!
0%
#515905000000
1!
1%
#515910000000
0!
0%
#515915000000
1!
1%
#515920000000
0!
0%
#515925000000
1!
1%
#515930000000
0!
0%
#515935000000
1!
1%
#515940000000
0!
0%
#515945000000
1!
1%
#515950000000
0!
0%
#515955000000
1!
1%
#515960000000
0!
0%
#515965000000
1!
1%
#515970000000
0!
0%
#515975000000
1!
1%
#515980000000
0!
0%
#515985000000
1!
1%
#515990000000
0!
0%
#515995000000
1!
1%
#516000000000
0!
0%
#516005000000
1!
1%
#516010000000
0!
0%
#516015000000
1!
1%
#516020000000
0!
0%
#516025000000
1!
1%
#516030000000
0!
0%
#516035000000
1!
1%
#516040000000
0!
0%
#516045000000
1!
1%
#516050000000
0!
0%
#516055000000
1!
1%
#516060000000
0!
0%
#516065000000
1!
1%
#516070000000
0!
0%
#516075000000
1!
1%
#516080000000
0!
0%
#516085000000
1!
1%
#516090000000
0!
0%
#516095000000
1!
1%
#516100000000
0!
0%
#516105000000
1!
1%
#516110000000
0!
0%
#516115000000
1!
1%
#516120000000
0!
0%
#516125000000
1!
1%
#516130000000
0!
0%
#516135000000
1!
1%
#516140000000
0!
0%
#516145000000
1!
1%
#516150000000
0!
0%
#516155000000
1!
1%
#516160000000
0!
0%
#516165000000
1!
1%
#516170000000
0!
0%
#516175000000
1!
1%
#516180000000
0!
0%
#516185000000
1!
1%
#516190000000
0!
0%
#516195000000
1!
1%
#516200000000
0!
0%
#516205000000
1!
1%
#516210000000
0!
0%
#516215000000
1!
1%
#516220000000
0!
0%
#516225000000
1!
1%
#516230000000
0!
0%
#516235000000
1!
1%
#516240000000
0!
0%
#516245000000
1!
1%
#516250000000
0!
0%
#516255000000
1!
1%
#516260000000
0!
0%
#516265000000
1!
1%
#516270000000
0!
0%
#516275000000
1!
1%
#516280000000
0!
0%
#516285000000
1!
1%
#516290000000
0!
0%
#516295000000
1!
1%
#516300000000
0!
0%
#516305000000
1!
1%
#516310000000
0!
0%
#516315000000
1!
1%
#516320000000
0!
0%
#516325000000
1!
1%
#516330000000
0!
0%
#516335000000
1!
1%
#516340000000
0!
0%
#516345000000
1!
1%
#516350000000
0!
0%
#516355000000
1!
1%
#516360000000
0!
0%
#516365000000
1!
1%
#516370000000
0!
0%
#516375000000
1!
1%
#516380000000
0!
0%
#516385000000
1!
1%
#516390000000
0!
0%
#516395000000
1!
1%
#516400000000
0!
0%
#516405000000
1!
1%
#516410000000
0!
0%
#516415000000
1!
1%
#516420000000
0!
0%
#516425000000
1!
1%
#516430000000
0!
0%
#516435000000
1!
1%
#516440000000
0!
0%
#516445000000
1!
1%
#516450000000
0!
0%
#516455000000
1!
1%
#516460000000
0!
0%
#516465000000
1!
1%
#516470000000
0!
0%
#516475000000
1!
1%
#516480000000
0!
0%
#516485000000
1!
1%
#516490000000
0!
0%
#516495000000
1!
1%
#516500000000
0!
0%
#516505000000
1!
1%
#516510000000
0!
0%
#516515000000
1!
1%
#516520000000
0!
0%
#516525000000
1!
1%
#516530000000
0!
0%
#516535000000
1!
1%
#516540000000
0!
0%
#516545000000
1!
1%
#516550000000
0!
0%
#516555000000
1!
1%
#516560000000
0!
0%
#516565000000
1!
1%
#516570000000
0!
0%
#516575000000
1!
1%
#516580000000
0!
0%
#516585000000
1!
1%
#516590000000
0!
0%
#516595000000
1!
1%
#516600000000
0!
0%
#516605000000
1!
1%
#516610000000
0!
0%
#516615000000
1!
1%
#516620000000
0!
0%
#516625000000
1!
1%
#516630000000
0!
0%
#516635000000
1!
1%
#516640000000
0!
0%
#516645000000
1!
1%
#516650000000
0!
0%
#516655000000
1!
1%
#516660000000
0!
0%
#516665000000
1!
1%
#516670000000
0!
0%
#516675000000
1!
1%
#516680000000
0!
0%
#516685000000
1!
1%
#516690000000
0!
0%
#516695000000
1!
1%
#516700000000
0!
0%
#516705000000
1!
1%
#516710000000
0!
0%
#516715000000
1!
1%
#516720000000
0!
0%
#516725000000
1!
1%
#516730000000
0!
0%
#516735000000
1!
1%
#516740000000
0!
0%
#516745000000
1!
1%
#516750000000
0!
0%
#516755000000
1!
1%
#516760000000
0!
0%
#516765000000
1!
1%
#516770000000
0!
0%
#516775000000
1!
1%
#516780000000
0!
0%
#516785000000
1!
1%
#516790000000
0!
0%
#516795000000
1!
1%
#516800000000
0!
0%
#516805000000
1!
1%
#516810000000
0!
0%
#516815000000
1!
1%
#516820000000
0!
0%
#516825000000
1!
1%
#516830000000
0!
0%
#516835000000
1!
1%
#516840000000
0!
0%
#516845000000
1!
1%
#516850000000
0!
0%
#516855000000
1!
1%
#516860000000
0!
0%
#516865000000
1!
1%
#516870000000
0!
0%
#516875000000
1!
1%
#516880000000
0!
0%
#516885000000
1!
1%
#516890000000
0!
0%
#516895000000
1!
1%
#516900000000
0!
0%
#516905000000
1!
1%
#516910000000
0!
0%
#516915000000
1!
1%
#516920000000
0!
0%
#516925000000
1!
1%
#516930000000
0!
0%
#516935000000
1!
1%
#516940000000
0!
0%
#516945000000
1!
1%
#516950000000
0!
0%
#516955000000
1!
1%
#516960000000
0!
0%
#516965000000
1!
1%
#516970000000
0!
0%
#516975000000
1!
1%
#516980000000
0!
0%
#516985000000
1!
1%
#516990000000
0!
0%
#516995000000
1!
1%
#517000000000
0!
0%
#517005000000
1!
1%
#517010000000
0!
0%
#517015000000
1!
1%
#517020000000
0!
0%
#517025000000
1!
1%
#517030000000
0!
0%
#517035000000
1!
1%
#517040000000
0!
0%
#517045000000
1!
1%
#517050000000
0!
0%
#517055000000
1!
1%
#517060000000
0!
0%
#517065000000
1!
1%
#517070000000
0!
0%
#517075000000
1!
1%
#517080000000
0!
0%
#517085000000
1!
1%
#517090000000
0!
0%
#517095000000
1!
1%
#517100000000
0!
0%
#517105000000
1!
1%
#517110000000
0!
0%
#517115000000
1!
1%
#517120000000
0!
0%
#517125000000
1!
1%
#517130000000
0!
0%
#517135000000
1!
1%
#517140000000
0!
0%
#517145000000
1!
1%
#517150000000
0!
0%
#517155000000
1!
1%
#517160000000
0!
0%
#517165000000
1!
1%
#517170000000
0!
0%
#517175000000
1!
1%
#517180000000
0!
0%
#517185000000
1!
1%
#517190000000
0!
0%
#517195000000
1!
1%
#517200000000
0!
0%
#517205000000
1!
1%
#517210000000
0!
0%
#517215000000
1!
1%
#517220000000
0!
0%
#517225000000
1!
1%
#517230000000
0!
0%
#517235000000
1!
1%
#517240000000
0!
0%
#517245000000
1!
1%
#517250000000
0!
0%
#517255000000
1!
1%
#517260000000
0!
0%
#517265000000
1!
1%
#517270000000
0!
0%
#517275000000
1!
1%
#517280000000
0!
0%
#517285000000
1!
1%
#517290000000
0!
0%
#517295000000
1!
1%
#517300000000
0!
0%
#517305000000
1!
1%
#517310000000
0!
0%
#517315000000
1!
1%
#517320000000
0!
0%
#517325000000
1!
1%
#517330000000
0!
0%
#517335000000
1!
1%
#517340000000
0!
0%
#517345000000
1!
1%
#517350000000
0!
0%
#517355000000
1!
1%
#517360000000
0!
0%
#517365000000
1!
1%
#517370000000
0!
0%
#517375000000
1!
1%
#517380000000
0!
0%
#517385000000
1!
1%
#517390000000
0!
0%
#517395000000
1!
1%
#517400000000
0!
0%
#517405000000
1!
1%
#517410000000
0!
0%
#517415000000
1!
1%
#517420000000
0!
0%
#517425000000
1!
1%
#517430000000
0!
0%
#517435000000
1!
1%
#517440000000
0!
0%
#517445000000
1!
1%
#517450000000
0!
0%
#517455000000
1!
1%
#517460000000
0!
0%
#517465000000
1!
1%
#517470000000
0!
0%
#517475000000
1!
1%
#517480000000
0!
0%
#517485000000
1!
1%
#517490000000
0!
0%
#517495000000
1!
1%
#517500000000
0!
0%
#517505000000
1!
1%
#517510000000
0!
0%
#517515000000
1!
1%
#517520000000
0!
0%
#517525000000
1!
1%
#517530000000
0!
0%
#517535000000
1!
1%
#517540000000
0!
0%
#517545000000
1!
1%
#517550000000
0!
0%
#517555000000
1!
1%
#517560000000
0!
0%
#517565000000
1!
1%
#517570000000
0!
0%
#517575000000
1!
1%
#517580000000
0!
0%
#517585000000
1!
1%
#517590000000
0!
0%
#517595000000
1!
1%
#517600000000
0!
0%
#517605000000
1!
1%
#517610000000
0!
0%
#517615000000
1!
1%
#517620000000
0!
0%
#517625000000
1!
1%
#517630000000
0!
0%
#517635000000
1!
1%
#517640000000
0!
0%
#517645000000
1!
1%
#517650000000
0!
0%
#517655000000
1!
1%
#517660000000
0!
0%
#517665000000
1!
1%
#517670000000
0!
0%
#517675000000
1!
1%
#517680000000
0!
0%
#517685000000
1!
1%
#517690000000
0!
0%
#517695000000
1!
1%
#517700000000
0!
0%
#517705000000
1!
1%
#517710000000
0!
0%
#517715000000
1!
1%
#517720000000
0!
0%
#517725000000
1!
1%
#517730000000
0!
0%
#517735000000
1!
1%
#517740000000
0!
0%
#517745000000
1!
1%
#517750000000
0!
0%
#517755000000
1!
1%
#517760000000
0!
0%
#517765000000
1!
1%
#517770000000
0!
0%
#517775000000
1!
1%
#517780000000
0!
0%
#517785000000
1!
1%
#517790000000
0!
0%
#517795000000
1!
1%
#517800000000
0!
0%
#517805000000
1!
1%
#517810000000
0!
0%
#517815000000
1!
1%
#517820000000
0!
0%
#517825000000
1!
1%
#517830000000
0!
0%
#517835000000
1!
1%
#517840000000
0!
0%
#517845000000
1!
1%
#517850000000
0!
0%
#517855000000
1!
1%
#517860000000
0!
0%
#517865000000
1!
1%
#517870000000
0!
0%
#517875000000
1!
1%
#517880000000
0!
0%
#517885000000
1!
1%
#517890000000
0!
0%
#517895000000
1!
1%
#517900000000
0!
0%
#517905000000
1!
1%
#517910000000
0!
0%
#517915000000
1!
1%
#517920000000
0!
0%
#517925000000
1!
1%
#517930000000
0!
0%
#517935000000
1!
1%
#517940000000
0!
0%
#517945000000
1!
1%
#517950000000
0!
0%
#517955000000
1!
1%
#517960000000
0!
0%
#517965000000
1!
1%
#517970000000
0!
0%
#517975000000
1!
1%
#517980000000
0!
0%
#517985000000
1!
1%
#517990000000
0!
0%
#517995000000
1!
1%
#518000000000
0!
0%
#518005000000
1!
1%
#518010000000
0!
0%
#518015000000
1!
1%
#518020000000
0!
0%
#518025000000
1!
1%
#518030000000
0!
0%
#518035000000
1!
1%
#518040000000
0!
0%
#518045000000
1!
1%
#518050000000
0!
0%
#518055000000
1!
1%
#518060000000
0!
0%
#518065000000
1!
1%
#518070000000
0!
0%
#518075000000
1!
1%
#518080000000
0!
0%
#518085000000
1!
1%
#518090000000
0!
0%
#518095000000
1!
1%
#518100000000
0!
0%
#518105000000
1!
1%
#518110000000
0!
0%
#518115000000
1!
1%
#518120000000
0!
0%
#518125000000
1!
1%
#518130000000
0!
0%
#518135000000
1!
1%
#518140000000
0!
0%
#518145000000
1!
1%
#518150000000
0!
0%
#518155000000
1!
1%
#518160000000
0!
0%
#518165000000
1!
1%
#518170000000
0!
0%
#518175000000
1!
1%
#518180000000
0!
0%
#518185000000
1!
1%
#518190000000
0!
0%
#518195000000
1!
1%
#518200000000
0!
0%
#518205000000
1!
1%
#518210000000
0!
0%
#518215000000
1!
1%
#518220000000
0!
0%
#518225000000
1!
1%
#518230000000
0!
0%
#518235000000
1!
1%
#518240000000
0!
0%
#518245000000
1!
1%
#518250000000
0!
0%
#518255000000
1!
1%
#518260000000
0!
0%
#518265000000
1!
1%
#518270000000
0!
0%
#518275000000
1!
1%
#518280000000
0!
0%
#518285000000
1!
1%
#518290000000
0!
0%
#518295000000
1!
1%
#518300000000
0!
0%
#518305000000
1!
1%
#518310000000
0!
0%
#518315000000
1!
1%
#518320000000
0!
0%
#518325000000
1!
1%
#518330000000
0!
0%
#518335000000
1!
1%
#518340000000
0!
0%
#518345000000
1!
1%
#518350000000
0!
0%
#518355000000
1!
1%
#518360000000
0!
0%
#518365000000
1!
1%
#518370000000
0!
0%
#518375000000
1!
1%
#518380000000
0!
0%
#518385000000
1!
1%
#518390000000
0!
0%
#518395000000
1!
1%
#518400000000
0!
0%
#518405000000
1!
1%
#518410000000
0!
0%
#518415000000
1!
1%
#518420000000
0!
0%
#518425000000
1!
1%
#518430000000
0!
0%
#518435000000
1!
1%
#518440000000
0!
0%
#518445000000
1!
1%
#518450000000
0!
0%
#518455000000
1!
1%
#518460000000
0!
0%
#518465000000
1!
1%
#518470000000
0!
0%
#518475000000
1!
1%
#518480000000
0!
0%
#518485000000
1!
1%
#518490000000
0!
0%
#518495000000
1!
1%
#518500000000
0!
0%
#518505000000
1!
1%
#518510000000
0!
0%
#518515000000
1!
1%
#518520000000
0!
0%
#518525000000
1!
1%
#518530000000
0!
0%
#518535000000
1!
1%
#518540000000
0!
0%
#518545000000
1!
1%
#518550000000
0!
0%
#518555000000
1!
1%
#518560000000
0!
0%
#518565000000
1!
1%
#518570000000
0!
0%
#518575000000
1!
1%
#518580000000
0!
0%
#518585000000
1!
1%
#518590000000
0!
0%
#518595000000
1!
1%
#518600000000
0!
0%
#518605000000
1!
1%
#518610000000
0!
0%
#518615000000
1!
1%
#518620000000
0!
0%
#518625000000
1!
1%
#518630000000
0!
0%
#518635000000
1!
1%
#518640000000
0!
0%
#518645000000
1!
1%
#518650000000
0!
0%
#518655000000
1!
1%
#518660000000
0!
0%
#518665000000
1!
1%
#518670000000
0!
0%
#518675000000
1!
1%
#518680000000
0!
0%
#518685000000
1!
1%
#518690000000
0!
0%
#518695000000
1!
1%
#518700000000
0!
0%
#518705000000
1!
1%
#518710000000
0!
0%
#518715000000
1!
1%
#518720000000
0!
0%
#518725000000
1!
1%
#518730000000
0!
0%
#518735000000
1!
1%
#518740000000
0!
0%
#518745000000
1!
1%
#518750000000
0!
0%
#518755000000
1!
1%
#518760000000
0!
0%
#518765000000
1!
1%
#518770000000
0!
0%
#518775000000
1!
1%
#518780000000
0!
0%
#518785000000
1!
1%
#518790000000
0!
0%
#518795000000
1!
1%
#518800000000
0!
0%
#518805000000
1!
1%
#518810000000
0!
0%
#518815000000
1!
1%
#518820000000
0!
0%
#518825000000
1!
1%
#518830000000
0!
0%
#518835000000
1!
1%
#518840000000
0!
0%
#518845000000
1!
1%
#518850000000
0!
0%
#518855000000
1!
1%
#518860000000
0!
0%
#518865000000
1!
1%
#518870000000
0!
0%
#518875000000
1!
1%
#518880000000
0!
0%
#518885000000
1!
1%
#518890000000
0!
0%
#518895000000
1!
1%
#518900000000
0!
0%
#518905000000
1!
1%
#518910000000
0!
0%
#518915000000
1!
1%
#518920000000
0!
0%
#518925000000
1!
1%
#518930000000
0!
0%
#518935000000
1!
1%
#518940000000
0!
0%
#518945000000
1!
1%
#518950000000
0!
0%
#518955000000
1!
1%
#518960000000
0!
0%
#518965000000
1!
1%
#518970000000
0!
0%
#518975000000
1!
1%
#518980000000
0!
0%
#518985000000
1!
1%
#518990000000
0!
0%
#518995000000
1!
1%
#519000000000
0!
0%
#519005000000
1!
1%
#519010000000
0!
0%
#519015000000
1!
1%
#519020000000
0!
0%
#519025000000
1!
1%
#519030000000
0!
0%
#519035000000
1!
1%
#519040000000
0!
0%
#519045000000
1!
1%
#519050000000
0!
0%
#519055000000
1!
1%
#519060000000
0!
0%
#519065000000
1!
1%
#519070000000
0!
0%
#519075000000
1!
1%
#519080000000
0!
0%
#519085000000
1!
1%
#519090000000
0!
0%
#519095000000
1!
1%
#519100000000
0!
0%
#519105000000
1!
1%
#519110000000
0!
0%
#519115000000
1!
1%
#519120000000
0!
0%
#519125000000
1!
1%
#519130000000
0!
0%
#519135000000
1!
1%
#519140000000
0!
0%
#519145000000
1!
1%
#519150000000
0!
0%
#519155000000
1!
1%
#519160000000
0!
0%
#519165000000
1!
1%
#519170000000
0!
0%
#519175000000
1!
1%
#519180000000
0!
0%
#519185000000
1!
1%
#519190000000
0!
0%
#519195000000
1!
1%
#519200000000
0!
0%
#519205000000
1!
1%
#519210000000
0!
0%
#519215000000
1!
1%
#519220000000
0!
0%
#519225000000
1!
1%
#519230000000
0!
0%
#519235000000
1!
1%
#519240000000
0!
0%
#519245000000
1!
1%
#519250000000
0!
0%
#519255000000
1!
1%
#519260000000
0!
0%
#519265000000
1!
1%
#519270000000
0!
0%
#519275000000
1!
1%
#519280000000
0!
0%
#519285000000
1!
1%
#519290000000
0!
0%
#519295000000
1!
1%
#519300000000
0!
0%
#519305000000
1!
1%
#519310000000
0!
0%
#519315000000
1!
1%
#519320000000
0!
0%
#519325000000
1!
1%
#519330000000
0!
0%
#519335000000
1!
1%
#519340000000
0!
0%
#519345000000
1!
1%
#519350000000
0!
0%
#519355000000
1!
1%
#519360000000
0!
0%
#519365000000
1!
1%
#519370000000
0!
0%
#519375000000
1!
1%
#519380000000
0!
0%
#519385000000
1!
1%
#519390000000
0!
0%
#519395000000
1!
1%
#519400000000
0!
0%
#519405000000
1!
1%
#519410000000
0!
0%
#519415000000
1!
1%
#519420000000
0!
0%
#519425000000
1!
1%
#519430000000
0!
0%
#519435000000
1!
1%
#519440000000
0!
0%
#519445000000
1!
1%
#519450000000
0!
0%
#519455000000
1!
1%
#519460000000
0!
0%
#519465000000
1!
1%
#519470000000
0!
0%
#519475000000
1!
1%
#519480000000
0!
0%
#519485000000
1!
1%
#519490000000
0!
0%
#519495000000
1!
1%
#519500000000
0!
0%
#519505000000
1!
1%
#519510000000
0!
0%
#519515000000
1!
1%
#519520000000
0!
0%
#519525000000
1!
1%
#519530000000
0!
0%
#519535000000
1!
1%
#519540000000
0!
0%
#519545000000
1!
1%
#519550000000
0!
0%
#519555000000
1!
1%
#519560000000
0!
0%
#519565000000
1!
1%
#519570000000
0!
0%
#519575000000
1!
1%
#519580000000
0!
0%
#519585000000
1!
1%
#519590000000
0!
0%
#519595000000
1!
1%
#519600000000
0!
0%
#519605000000
1!
1%
#519610000000
0!
0%
#519615000000
1!
1%
#519620000000
0!
0%
#519625000000
1!
1%
#519630000000
0!
0%
#519635000000
1!
1%
#519640000000
0!
0%
#519645000000
1!
1%
#519650000000
0!
0%
#519655000000
1!
1%
#519660000000
0!
0%
#519665000000
1!
1%
#519670000000
0!
0%
#519675000000
1!
1%
#519680000000
0!
0%
#519685000000
1!
1%
#519690000000
0!
0%
#519695000000
1!
1%
#519700000000
0!
0%
#519705000000
1!
1%
#519710000000
0!
0%
#519715000000
1!
1%
#519720000000
0!
0%
#519725000000
1!
1%
#519730000000
0!
0%
#519735000000
1!
1%
#519740000000
0!
0%
#519745000000
1!
1%
#519750000000
0!
0%
#519755000000
1!
1%
#519760000000
0!
0%
#519765000000
1!
1%
#519770000000
0!
0%
#519775000000
1!
1%
#519780000000
0!
0%
#519785000000
1!
1%
#519790000000
0!
0%
#519795000000
1!
1%
#519800000000
0!
0%
#519805000000
1!
1%
#519810000000
0!
0%
#519815000000
1!
1%
#519820000000
0!
0%
#519825000000
1!
1%
#519830000000
0!
0%
#519835000000
1!
1%
#519840000000
0!
0%
#519845000000
1!
1%
#519850000000
0!
0%
#519855000000
1!
1%
#519860000000
0!
0%
#519865000000
1!
1%
#519870000000
0!
0%
#519875000000
1!
1%
#519880000000
0!
0%
#519885000000
1!
1%
#519890000000
0!
0%
#519895000000
1!
1%
#519900000000
0!
0%
#519905000000
1!
1%
#519910000000
0!
0%
#519915000000
1!
1%
#519920000000
0!
0%
#519925000000
1!
1%
#519930000000
0!
0%
#519935000000
1!
1%
#519940000000
0!
0%
#519945000000
1!
1%
#519950000000
0!
0%
#519955000000
1!
1%
#519960000000
0!
0%
#519965000000
1!
1%
#519970000000
0!
0%
#519975000000
1!
1%
#519980000000
0!
0%
#519985000000
1!
1%
#519990000000
0!
0%
#519995000000
1!
1%
#520000000000
0!
0%
#520005000000
1!
1%
#520010000000
0!
0%
#520015000000
1!
1%
#520020000000
0!
0%
#520025000000
1!
1%
#520030000000
0!
0%
#520035000000
1!
1%
#520040000000
0!
0%
#520045000000
1!
1%
#520050000000
0!
0%
#520055000000
1!
1%
#520060000000
0!
0%
#520065000000
1!
1%
#520070000000
0!
0%
#520075000000
1!
1%
#520080000000
0!
0%
#520085000000
1!
1%
#520090000000
0!
0%
#520095000000
1!
1%
#520100000000
0!
0%
#520105000000
1!
1%
#520110000000
0!
0%
#520115000000
1!
1%
#520120000000
0!
0%
#520125000000
1!
1%
#520130000000
0!
0%
#520135000000
1!
1%
#520140000000
0!
0%
#520145000000
1!
1%
#520150000000
0!
0%
#520155000000
1!
1%
#520160000000
0!
0%
#520165000000
1!
1%
#520170000000
0!
0%
#520175000000
1!
1%
#520180000000
0!
0%
#520185000000
1!
1%
#520190000000
0!
0%
#520195000000
1!
1%
#520200000000
0!
0%
#520205000000
1!
1%
#520210000000
0!
0%
#520215000000
1!
1%
#520220000000
0!
0%
#520225000000
1!
1%
#520230000000
0!
0%
#520235000000
1!
1%
#520240000000
0!
0%
#520245000000
1!
1%
#520250000000
0!
0%
#520255000000
1!
1%
#520260000000
0!
0%
#520265000000
1!
1%
#520270000000
0!
0%
#520275000000
1!
1%
#520280000000
0!
0%
#520285000000
1!
1%
#520290000000
0!
0%
#520295000000
1!
1%
#520300000000
0!
0%
#520305000000
1!
1%
#520310000000
0!
0%
#520315000000
1!
1%
#520320000000
0!
0%
#520325000000
1!
1%
#520330000000
0!
0%
#520335000000
1!
1%
#520340000000
0!
0%
#520345000000
1!
1%
#520350000000
0!
0%
#520355000000
1!
1%
#520360000000
0!
0%
#520365000000
1!
1%
#520370000000
0!
0%
#520375000000
1!
1%
#520380000000
0!
0%
#520385000000
1!
1%
#520390000000
0!
0%
#520395000000
1!
1%
#520400000000
0!
0%
#520405000000
1!
1%
#520410000000
0!
0%
#520415000000
1!
1%
#520420000000
0!
0%
#520425000000
1!
1%
#520430000000
0!
0%
#520435000000
1!
1%
#520440000000
0!
0%
#520445000000
1!
1%
#520450000000
0!
0%
#520455000000
1!
1%
#520460000000
0!
0%
#520465000000
1!
1%
#520470000000
0!
0%
#520475000000
1!
1%
#520480000000
0!
0%
#520485000000
1!
1%
#520490000000
0!
0%
#520495000000
1!
1%
#520500000000
0!
0%
#520505000000
1!
1%
#520510000000
0!
0%
#520515000000
1!
1%
#520520000000
0!
0%
#520525000000
1!
1%
#520530000000
0!
0%
#520535000000
1!
1%
#520540000000
0!
0%
#520545000000
1!
1%
#520550000000
0!
0%
#520555000000
1!
1%
#520560000000
0!
0%
#520565000000
1!
1%
#520570000000
0!
0%
#520575000000
1!
1%
#520580000000
0!
0%
#520585000000
1!
1%
#520590000000
0!
0%
#520595000000
1!
1%
#520600000000
0!
0%
#520605000000
1!
1%
#520610000000
0!
0%
#520615000000
1!
1%
#520620000000
0!
0%
#520625000000
1!
1%
#520630000000
0!
0%
#520635000000
1!
1%
#520640000000
0!
0%
#520645000000
1!
1%
#520650000000
0!
0%
#520655000000
1!
1%
#520660000000
0!
0%
#520665000000
1!
1%
#520670000000
0!
0%
#520675000000
1!
1%
#520680000000
0!
0%
#520685000000
1!
1%
#520690000000
0!
0%
#520695000000
1!
1%
#520700000000
0!
0%
#520705000000
1!
1%
#520710000000
0!
0%
#520715000000
1!
1%
#520720000000
0!
0%
#520725000000
1!
1%
#520730000000
0!
0%
#520735000000
1!
1%
#520740000000
0!
0%
#520745000000
1!
1%
#520750000000
0!
0%
#520755000000
1!
1%
#520760000000
0!
0%
#520765000000
1!
1%
#520770000000
0!
0%
#520775000000
1!
1%
#520780000000
0!
0%
#520785000000
1!
1%
#520790000000
0!
0%
#520795000000
1!
1%
#520800000000
0!
0%
#520805000000
1!
1%
#520810000000
0!
0%
#520815000000
1!
1%
#520820000000
0!
0%
#520825000000
1!
1%
#520830000000
0!
0%
#520835000000
1!
1%
#520840000000
0!
0%
#520845000000
1!
1%
#520850000000
0!
0%
#520855000000
1!
1%
#520860000000
0!
0%
#520865000000
1!
1%
#520870000000
0!
0%
#520875000000
1!
1%
#520880000000
0!
0%
#520885000000
1!
1%
#520890000000
0!
0%
#520895000000
1!
1%
#520900000000
0!
0%
#520905000000
1!
1%
#520910000000
0!
0%
#520915000000
1!
1%
#520920000000
0!
0%
#520925000000
1!
1%
#520930000000
0!
0%
#520935000000
1!
1%
#520940000000
0!
0%
#520945000000
1!
1%
#520950000000
0!
0%
#520955000000
1!
1%
#520960000000
0!
0%
#520965000000
1!
1%
#520970000000
0!
0%
#520975000000
1!
1%
#520980000000
0!
0%
#520985000000
1!
1%
#520990000000
0!
0%
#520995000000
1!
1%
#521000000000
0!
0%
#521005000000
1!
1%
#521010000000
0!
0%
#521015000000
1!
1%
#521020000000
0!
0%
#521025000000
1!
1%
#521030000000
0!
0%
#521035000000
1!
1%
#521040000000
0!
0%
#521045000000
1!
1%
#521050000000
0!
0%
#521055000000
1!
1%
#521060000000
0!
0%
#521065000000
1!
1%
#521070000000
0!
0%
#521075000000
1!
1%
#521080000000
0!
0%
#521085000000
1!
1%
#521090000000
0!
0%
#521095000000
1!
1%
#521100000000
0!
0%
#521105000000
1!
1%
#521110000000
0!
0%
#521115000000
1!
1%
#521120000000
0!
0%
#521125000000
1!
1%
#521130000000
0!
0%
#521135000000
1!
1%
#521140000000
0!
0%
#521145000000
1!
1%
#521150000000
0!
0%
#521155000000
1!
1%
#521160000000
0!
0%
#521165000000
1!
1%
#521170000000
0!
0%
#521175000000
1!
1%
#521180000000
0!
0%
#521185000000
1!
1%
#521190000000
0!
0%
#521195000000
1!
1%
#521200000000
0!
0%
#521205000000
1!
1%
#521210000000
0!
0%
#521215000000
1!
1%
#521220000000
0!
0%
#521225000000
1!
1%
#521230000000
0!
0%
#521235000000
1!
1%
#521240000000
0!
0%
#521245000000
1!
1%
#521250000000
0!
0%
#521255000000
1!
1%
#521260000000
0!
0%
#521265000000
1!
1%
#521270000000
0!
0%
#521275000000
1!
1%
#521280000000
0!
0%
#521285000000
1!
1%
#521290000000
0!
0%
#521295000000
1!
1%
#521300000000
0!
0%
#521305000000
1!
1%
#521310000000
0!
0%
#521315000000
1!
1%
#521320000000
0!
0%
#521325000000
1!
1%
#521330000000
0!
0%
#521335000000
1!
1%
#521340000000
0!
0%
#521345000000
1!
1%
#521350000000
0!
0%
#521355000000
1!
1%
#521360000000
0!
0%
#521365000000
1!
1%
#521370000000
0!
0%
#521375000000
1!
1%
#521380000000
0!
0%
#521385000000
1!
1%
#521390000000
0!
0%
#521395000000
1!
1%
#521400000000
0!
0%
#521405000000
1!
1%
#521410000000
0!
0%
#521415000000
1!
1%
#521420000000
0!
0%
#521425000000
1!
1%
#521430000000
0!
0%
#521435000000
1!
1%
#521440000000
0!
0%
#521445000000
1!
1%
#521450000000
0!
0%
#521455000000
1!
1%
#521460000000
0!
0%
#521465000000
1!
1%
#521470000000
0!
0%
#521475000000
1!
1%
#521480000000
0!
0%
#521485000000
1!
1%
#521490000000
0!
0%
#521495000000
1!
1%
#521500000000
0!
0%
#521505000000
1!
1%
#521510000000
0!
0%
#521515000000
1!
1%
#521520000000
0!
0%
#521525000000
1!
1%
#521530000000
0!
0%
#521535000000
1!
1%
#521540000000
0!
0%
#521545000000
1!
1%
#521550000000
0!
0%
#521555000000
1!
1%
#521560000000
0!
0%
#521565000000
1!
1%
#521570000000
0!
0%
#521575000000
1!
1%
#521580000000
0!
0%
#521585000000
1!
1%
#521590000000
0!
0%
#521595000000
1!
1%
#521600000000
0!
0%
#521605000000
1!
1%
#521610000000
0!
0%
#521615000000
1!
1%
#521620000000
0!
0%
#521625000000
1!
1%
#521630000000
0!
0%
#521635000000
1!
1%
#521640000000
0!
0%
#521645000000
1!
1%
#521650000000
0!
0%
#521655000000
1!
1%
#521660000000
0!
0%
#521665000000
1!
1%
#521670000000
0!
0%
#521675000000
1!
1%
#521680000000
0!
0%
#521685000000
1!
1%
#521690000000
0!
0%
#521695000000
1!
1%
#521700000000
0!
0%
#521705000000
1!
1%
#521710000000
0!
0%
#521715000000
1!
1%
#521720000000
0!
0%
#521725000000
1!
1%
#521730000000
0!
0%
#521735000000
1!
1%
#521740000000
0!
0%
#521745000000
1!
1%
#521750000000
0!
0%
#521755000000
1!
1%
#521760000000
0!
0%
#521765000000
1!
1%
#521770000000
0!
0%
#521775000000
1!
1%
#521780000000
0!
0%
#521785000000
1!
1%
#521790000000
0!
0%
#521795000000
1!
1%
#521800000000
0!
0%
#521805000000
1!
1%
#521810000000
0!
0%
#521815000000
1!
1%
#521820000000
0!
0%
#521825000000
1!
1%
#521830000000
0!
0%
#521835000000
1!
1%
#521840000000
0!
0%
#521845000000
1!
1%
#521850000000
0!
0%
#521855000000
1!
1%
#521860000000
0!
0%
#521865000000
1!
1%
#521870000000
0!
0%
#521875000000
1!
1%
#521880000000
0!
0%
#521885000000
1!
1%
#521890000000
0!
0%
#521895000000
1!
1%
#521900000000
0!
0%
#521905000000
1!
1%
#521910000000
0!
0%
#521915000000
1!
1%
#521920000000
0!
0%
#521925000000
1!
1%
#521930000000
0!
0%
#521935000000
1!
1%
#521940000000
0!
0%
#521945000000
1!
1%
#521950000000
0!
0%
#521955000000
1!
1%
#521960000000
0!
0%
#521965000000
1!
1%
#521970000000
0!
0%
#521975000000
1!
1%
#521980000000
0!
0%
#521985000000
1!
1%
#521990000000
0!
0%
#521995000000
1!
1%
#522000000000
0!
0%
#522005000000
1!
1%
#522010000000
0!
0%
#522015000000
1!
1%
#522020000000
0!
0%
#522025000000
1!
1%
#522030000000
0!
0%
#522035000000
1!
1%
#522040000000
0!
0%
#522045000000
1!
1%
#522050000000
0!
0%
#522055000000
1!
1%
#522060000000
0!
0%
#522065000000
1!
1%
#522070000000
0!
0%
#522075000000
1!
1%
#522080000000
0!
0%
#522085000000
1!
1%
#522090000000
0!
0%
#522095000000
1!
1%
#522100000000
0!
0%
#522105000000
1!
1%
#522110000000
0!
0%
#522115000000
1!
1%
#522120000000
0!
0%
#522125000000
1!
1%
#522130000000
0!
0%
#522135000000
1!
1%
#522140000000
0!
0%
#522145000000
1!
1%
#522150000000
0!
0%
#522155000000
1!
1%
#522160000000
0!
0%
#522165000000
1!
1%
#522170000000
0!
0%
#522175000000
1!
1%
#522180000000
0!
0%
#522185000000
1!
1%
#522190000000
0!
0%
#522195000000
1!
1%
#522200000000
0!
0%
#522205000000
1!
1%
#522210000000
0!
0%
#522215000000
1!
1%
#522220000000
0!
0%
#522225000000
1!
1%
#522230000000
0!
0%
#522235000000
1!
1%
#522240000000
0!
0%
#522245000000
1!
1%
#522250000000
0!
0%
#522255000000
1!
1%
#522260000000
0!
0%
#522265000000
1!
1%
#522270000000
0!
0%
#522275000000
1!
1%
#522280000000
0!
0%
#522285000000
1!
1%
#522290000000
0!
0%
#522295000000
1!
1%
#522300000000
0!
0%
#522305000000
1!
1%
#522310000000
0!
0%
#522315000000
1!
1%
#522320000000
0!
0%
#522325000000
1!
1%
#522330000000
0!
0%
#522335000000
1!
1%
#522340000000
0!
0%
#522345000000
1!
1%
#522350000000
0!
0%
#522355000000
1!
1%
#522360000000
0!
0%
#522365000000
1!
1%
#522370000000
0!
0%
#522375000000
1!
1%
#522380000000
0!
0%
#522385000000
1!
1%
#522390000000
0!
0%
#522395000000
1!
1%
#522400000000
0!
0%
#522405000000
1!
1%
#522410000000
0!
0%
#522415000000
1!
1%
#522420000000
0!
0%
#522425000000
1!
1%
#522430000000
0!
0%
#522435000000
1!
1%
#522440000000
0!
0%
#522445000000
1!
1%
#522450000000
0!
0%
#522455000000
1!
1%
#522460000000
0!
0%
#522465000000
1!
1%
#522470000000
0!
0%
#522475000000
1!
1%
#522480000000
0!
0%
#522485000000
1!
1%
#522490000000
0!
0%
#522495000000
1!
1%
#522500000000
0!
0%
#522505000000
1!
1%
#522510000000
0!
0%
#522515000000
1!
1%
#522520000000
0!
0%
#522525000000
1!
1%
#522530000000
0!
0%
#522535000000
1!
1%
#522540000000
0!
0%
#522545000000
1!
1%
#522550000000
0!
0%
#522555000000
1!
1%
#522560000000
0!
0%
#522565000000
1!
1%
#522570000000
0!
0%
#522575000000
1!
1%
#522580000000
0!
0%
#522585000000
1!
1%
#522590000000
0!
0%
#522595000000
1!
1%
#522600000000
0!
0%
#522605000000
1!
1%
#522610000000
0!
0%
#522615000000
1!
1%
#522620000000
0!
0%
#522625000000
1!
1%
#522630000000
0!
0%
#522635000000
1!
1%
#522640000000
0!
0%
#522645000000
1!
1%
#522650000000
0!
0%
#522655000000
1!
1%
#522660000000
0!
0%
#522665000000
1!
1%
#522670000000
0!
0%
#522675000000
1!
1%
#522680000000
0!
0%
#522685000000
1!
1%
#522690000000
0!
0%
#522695000000
1!
1%
#522700000000
0!
0%
#522705000000
1!
1%
#522710000000
0!
0%
#522715000000
1!
1%
#522720000000
0!
0%
#522725000000
1!
1%
#522730000000
0!
0%
#522735000000
1!
1%
#522740000000
0!
0%
#522745000000
1!
1%
#522750000000
0!
0%
#522755000000
1!
1%
#522760000000
0!
0%
#522765000000
1!
1%
#522770000000
0!
0%
#522775000000
1!
1%
#522780000000
0!
0%
#522785000000
1!
1%
#522790000000
0!
0%
#522795000000
1!
1%
#522800000000
0!
0%
#522805000000
1!
1%
#522810000000
0!
0%
#522815000000
1!
1%
#522820000000
0!
0%
#522825000000
1!
1%
#522830000000
0!
0%
#522835000000
1!
1%
#522840000000
0!
0%
#522845000000
1!
1%
#522850000000
0!
0%
#522855000000
1!
1%
#522860000000
0!
0%
#522865000000
1!
1%
#522870000000
0!
0%
#522875000000
1!
1%
#522880000000
0!
0%
#522885000000
1!
1%
#522890000000
0!
0%
#522895000000
1!
1%
#522900000000
0!
0%
#522905000000
1!
1%
#522910000000
0!
0%
#522915000000
1!
1%
#522920000000
0!
0%
#522925000000
1!
1%
#522930000000
0!
0%
#522935000000
1!
1%
#522940000000
0!
0%
#522945000000
1!
1%
#522950000000
0!
0%
#522955000000
1!
1%
#522960000000
0!
0%
#522965000000
1!
1%
#522970000000
0!
0%
#522975000000
1!
1%
#522980000000
0!
0%
#522985000000
1!
1%
#522990000000
0!
0%
#522995000000
1!
1%
#523000000000
0!
0%
#523005000000
1!
1%
#523010000000
0!
0%
#523015000000
1!
1%
#523020000000
0!
0%
#523025000000
1!
1%
#523030000000
0!
0%
#523035000000
1!
1%
#523040000000
0!
0%
#523045000000
1!
1%
#523050000000
0!
0%
#523055000000
1!
1%
#523060000000
0!
0%
#523065000000
1!
1%
#523070000000
0!
0%
#523075000000
1!
1%
#523080000000
0!
0%
#523085000000
1!
1%
#523090000000
0!
0%
#523095000000
1!
1%
#523100000000
0!
0%
#523105000000
1!
1%
#523110000000
0!
0%
#523115000000
1!
1%
#523120000000
0!
0%
#523125000000
1!
1%
#523130000000
0!
0%
#523135000000
1!
1%
#523140000000
0!
0%
#523145000000
1!
1%
#523150000000
0!
0%
#523155000000
1!
1%
#523160000000
0!
0%
#523165000000
1!
1%
#523170000000
0!
0%
#523175000000
1!
1%
#523180000000
0!
0%
#523185000000
1!
1%
#523190000000
0!
0%
#523195000000
1!
1%
#523200000000
0!
0%
#523205000000
1!
1%
#523210000000
0!
0%
#523215000000
1!
1%
#523220000000
0!
0%
#523225000000
1!
1%
#523230000000
0!
0%
#523235000000
1!
1%
#523240000000
0!
0%
#523245000000
1!
1%
#523250000000
0!
0%
#523255000000
1!
1%
#523260000000
0!
0%
#523265000000
1!
1%
#523270000000
0!
0%
#523275000000
1!
1%
#523280000000
0!
0%
#523285000000
1!
1%
#523290000000
0!
0%
#523295000000
1!
1%
#523300000000
0!
0%
#523305000000
1!
1%
#523310000000
0!
0%
#523315000000
1!
1%
#523320000000
0!
0%
#523325000000
1!
1%
#523330000000
0!
0%
#523335000000
1!
1%
#523340000000
0!
0%
#523345000000
1!
1%
#523350000000
0!
0%
#523355000000
1!
1%
#523360000000
0!
0%
#523365000000
1!
1%
#523370000000
0!
0%
#523375000000
1!
1%
#523380000000
0!
0%
#523385000000
1!
1%
#523390000000
0!
0%
#523395000000
1!
1%
#523400000000
0!
0%
#523405000000
1!
1%
#523410000000
0!
0%
#523415000000
1!
1%
#523420000000
0!
0%
#523425000000
1!
1%
#523430000000
0!
0%
#523435000000
1!
1%
#523440000000
0!
0%
#523445000000
1!
1%
#523450000000
0!
0%
#523455000000
1!
1%
#523460000000
0!
0%
#523465000000
1!
1%
#523470000000
0!
0%
#523475000000
1!
1%
#523480000000
0!
0%
#523485000000
1!
1%
#523490000000
0!
0%
#523495000000
1!
1%
#523500000000
0!
0%
#523505000000
1!
1%
#523510000000
0!
0%
#523515000000
1!
1%
#523520000000
0!
0%
#523525000000
1!
1%
#523530000000
0!
0%
#523535000000
1!
1%
#523540000000
0!
0%
#523545000000
1!
1%
#523550000000
0!
0%
#523555000000
1!
1%
#523560000000
0!
0%
#523565000000
1!
1%
#523570000000
0!
0%
#523575000000
1!
1%
#523580000000
0!
0%
#523585000000
1!
1%
#523590000000
0!
0%
#523595000000
1!
1%
#523600000000
0!
0%
#523605000000
1!
1%
#523610000000
0!
0%
#523615000000
1!
1%
#523620000000
0!
0%
#523625000000
1!
1%
#523630000000
0!
0%
#523635000000
1!
1%
#523640000000
0!
0%
#523645000000
1!
1%
#523650000000
0!
0%
#523655000000
1!
1%
#523660000000
0!
0%
#523665000000
1!
1%
#523670000000
0!
0%
#523675000000
1!
1%
#523680000000
0!
0%
#523685000000
1!
1%
#523690000000
0!
0%
#523695000000
1!
1%
#523700000000
0!
0%
#523705000000
1!
1%
#523710000000
0!
0%
#523715000000
1!
1%
#523720000000
0!
0%
#523725000000
1!
1%
#523730000000
0!
0%
#523735000000
1!
1%
#523740000000
0!
0%
#523745000000
1!
1%
#523750000000
0!
0%
#523755000000
1!
1%
#523760000000
0!
0%
#523765000000
1!
1%
#523770000000
0!
0%
#523775000000
1!
1%
#523780000000
0!
0%
#523785000000
1!
1%
#523790000000
0!
0%
#523795000000
1!
1%
#523800000000
0!
0%
#523805000000
1!
1%
#523810000000
0!
0%
#523815000000
1!
1%
#523820000000
0!
0%
#523825000000
1!
1%
#523830000000
0!
0%
#523835000000
1!
1%
#523840000000
0!
0%
#523845000000
1!
1%
#523850000000
0!
0%
#523855000000
1!
1%
#523860000000
0!
0%
#523865000000
1!
1%
#523870000000
0!
0%
#523875000000
1!
1%
#523880000000
0!
0%
#523885000000
1!
1%
#523890000000
0!
0%
#523895000000
1!
1%
#523900000000
0!
0%
#523905000000
1!
1%
#523910000000
0!
0%
#523915000000
1!
1%
#523920000000
0!
0%
#523925000000
1!
1%
#523930000000
0!
0%
#523935000000
1!
1%
#523940000000
0!
0%
#523945000000
1!
1%
#523950000000
0!
0%
#523955000000
1!
1%
#523960000000
0!
0%
#523965000000
1!
1%
#523970000000
0!
0%
#523975000000
1!
1%
#523980000000
0!
0%
#523985000000
1!
1%
#523990000000
0!
0%
#523995000000
1!
1%
#524000000000
0!
0%
#524005000000
1!
1%
#524010000000
0!
0%
#524015000000
1!
1%
#524020000000
0!
0%
#524025000000
1!
1%
#524030000000
0!
0%
#524035000000
1!
1%
#524040000000
0!
0%
#524045000000
1!
1%
#524050000000
0!
0%
#524055000000
1!
1%
#524060000000
0!
0%
#524065000000
1!
1%
#524070000000
0!
0%
#524075000000
1!
1%
#524080000000
0!
0%
#524085000000
1!
1%
#524090000000
0!
0%
#524095000000
1!
1%
#524100000000
0!
0%
#524105000000
1!
1%
#524110000000
0!
0%
#524115000000
1!
1%
#524120000000
0!
0%
#524125000000
1!
1%
#524130000000
0!
0%
#524135000000
1!
1%
#524140000000
0!
0%
#524145000000
1!
1%
#524150000000
0!
0%
#524155000000
1!
1%
#524160000000
0!
0%
#524165000000
1!
1%
#524170000000
0!
0%
#524175000000
1!
1%
#524180000000
0!
0%
#524185000000
1!
1%
#524190000000
0!
0%
#524195000000
1!
1%
#524200000000
0!
0%
#524205000000
1!
1%
#524210000000
0!
0%
#524215000000
1!
1%
#524220000000
0!
0%
#524225000000
1!
1%
#524230000000
0!
0%
#524235000000
1!
1%
#524240000000
0!
0%
#524245000000
1!
1%
#524250000000
0!
0%
#524255000000
1!
1%
#524260000000
0!
0%
#524265000000
1!
1%
#524270000000
0!
0%
#524275000000
1!
1%
#524280000000
0!
0%
#524285000000
1!
1%
#524290000000
0!
0%
#524295000000
1!
1%
#524300000000
0!
0%
#524305000000
1!
1%
#524310000000
0!
0%
#524315000000
1!
1%
#524320000000
0!
0%
#524325000000
1!
1%
#524330000000
0!
0%
#524335000000
1!
1%
#524340000000
0!
0%
#524345000000
1!
1%
#524350000000
0!
0%
#524355000000
1!
1%
#524360000000
0!
0%
#524365000000
1!
1%
#524370000000
0!
0%
#524375000000
1!
1%
#524380000000
0!
0%
#524385000000
1!
1%
#524390000000
0!
0%
#524395000000
1!
1%
#524400000000
0!
0%
#524405000000
1!
1%
#524410000000
0!
0%
#524415000000
1!
1%
#524420000000
0!
0%
#524425000000
1!
1%
#524430000000
0!
0%
#524435000000
1!
1%
#524440000000
0!
0%
#524445000000
1!
1%
#524450000000
0!
0%
#524455000000
1!
1%
#524460000000
0!
0%
#524465000000
1!
1%
#524470000000
0!
0%
#524475000000
1!
1%
#524480000000
0!
0%
#524485000000
1!
1%
#524490000000
0!
0%
#524495000000
1!
1%
#524500000000
0!
0%
#524505000000
1!
1%
#524510000000
0!
0%
#524515000000
1!
1%
#524520000000
0!
0%
#524525000000
1!
1%
#524530000000
0!
0%
#524535000000
1!
1%
#524540000000
0!
0%
#524545000000
1!
1%
#524550000000
0!
0%
#524555000000
1!
1%
#524560000000
0!
0%
#524565000000
1!
1%
#524570000000
0!
0%
#524575000000
1!
1%
#524580000000
0!
0%
#524585000000
1!
1%
#524590000000
0!
0%
#524595000000
1!
1%
#524600000000
0!
0%
#524605000000
1!
1%
#524610000000
0!
0%
#524615000000
1!
1%
#524620000000
0!
0%
#524625000000
1!
1%
#524630000000
0!
0%
#524635000000
1!
1%
#524640000000
0!
0%
#524645000000
1!
1%
#524650000000
0!
0%
#524655000000
1!
1%
#524660000000
0!
0%
#524665000000
1!
1%
#524670000000
0!
0%
#524675000000
1!
1%
#524680000000
0!
0%
#524685000000
1!
1%
#524690000000
0!
0%
#524695000000
1!
1%
#524700000000
0!
0%
#524705000000
1!
1%
#524710000000
0!
0%
#524715000000
1!
1%
#524720000000
0!
0%
#524725000000
1!
1%
#524730000000
0!
0%
#524735000000
1!
1%
#524740000000
0!
0%
#524745000000
1!
1%
#524750000000
0!
0%
#524755000000
1!
1%
#524760000000
0!
0%
#524765000000
1!
1%
#524770000000
0!
0%
#524775000000
1!
1%
#524780000000
0!
0%
#524785000000
1!
1%
#524790000000
0!
0%
#524795000000
1!
1%
#524800000000
0!
0%
#524805000000
1!
1%
#524810000000
0!
0%
#524815000000
1!
1%
#524820000000
0!
0%
#524825000000
1!
1%
#524830000000
0!
0%
#524835000000
1!
1%
#524840000000
0!
0%
#524845000000
1!
1%
#524850000000
0!
0%
#524855000000
1!
1%
#524860000000
0!
0%
#524865000000
1!
1%
#524870000000
0!
0%
#524875000000
1!
1%
#524880000000
0!
0%
#524885000000
1!
1%
#524890000000
0!
0%
#524895000000
1!
1%
#524900000000
0!
0%
#524905000000
1!
1%
#524910000000
0!
0%
#524915000000
1!
1%
#524920000000
0!
0%
#524925000000
1!
1%
#524930000000
0!
0%
#524935000000
1!
1%
#524940000000
0!
0%
#524945000000
1!
1%
#524950000000
0!
0%
#524955000000
1!
1%
#524960000000
0!
0%
#524965000000
1!
1%
#524970000000
0!
0%
#524975000000
1!
1%
#524980000000
0!
0%
#524985000000
1!
1%
#524990000000
0!
0%
#524995000000
1!
1%
#525000000000
0!
0%
#525005000000
1!
1%
#525010000000
0!
0%
#525015000000
1!
1%
#525020000000
0!
0%
#525025000000
1!
1%
#525030000000
0!
0%
#525035000000
1!
1%
#525040000000
0!
0%
#525045000000
1!
1%
#525050000000
0!
0%
#525055000000
1!
1%
#525060000000
0!
0%
#525065000000
1!
1%
#525070000000
0!
0%
#525075000000
1!
1%
#525080000000
0!
0%
#525085000000
1!
1%
#525090000000
0!
0%
#525095000000
1!
1%
#525100000000
0!
0%
#525105000000
1!
1%
#525110000000
0!
0%
#525115000000
1!
1%
#525120000000
0!
0%
#525125000000
1!
1%
#525130000000
0!
0%
#525135000000
1!
1%
#525140000000
0!
0%
#525145000000
1!
1%
#525150000000
0!
0%
#525155000000
1!
1%
#525160000000
0!
0%
#525165000000
1!
1%
#525170000000
0!
0%
#525175000000
1!
1%
#525180000000
0!
0%
#525185000000
1!
1%
#525190000000
0!
0%
#525195000000
1!
1%
#525200000000
0!
0%
#525205000000
1!
1%
#525210000000
0!
0%
#525215000000
1!
1%
#525220000000
0!
0%
#525225000000
1!
1%
#525230000000
0!
0%
#525235000000
1!
1%
#525240000000
0!
0%
#525245000000
1!
1%
#525250000000
0!
0%
#525255000000
1!
1%
#525260000000
0!
0%
#525265000000
1!
1%
#525270000000
0!
0%
#525275000000
1!
1%
#525280000000
0!
0%
#525285000000
1!
1%
#525290000000
0!
0%
#525295000000
1!
1%
#525300000000
0!
0%
#525305000000
1!
1%
#525310000000
0!
0%
#525315000000
1!
1%
#525320000000
0!
0%
#525325000000
1!
1%
#525330000000
0!
0%
#525335000000
1!
1%
#525340000000
0!
0%
#525345000000
1!
1%
#525350000000
0!
0%
#525355000000
1!
1%
#525360000000
0!
0%
#525365000000
1!
1%
#525370000000
0!
0%
#525375000000
1!
1%
#525380000000
0!
0%
#525385000000
1!
1%
#525390000000
0!
0%
#525395000000
1!
1%
#525400000000
0!
0%
#525405000000
1!
1%
#525410000000
0!
0%
#525415000000
1!
1%
#525420000000
0!
0%
#525425000000
1!
1%
#525430000000
0!
0%
#525435000000
1!
1%
#525440000000
0!
0%
#525445000000
1!
1%
#525450000000
0!
0%
#525455000000
1!
1%
#525460000000
0!
0%
#525465000000
1!
1%
#525470000000
0!
0%
#525475000000
1!
1%
#525480000000
0!
0%
#525485000000
1!
1%
#525490000000
0!
0%
#525495000000
1!
1%
#525500000000
0!
0%
#525505000000
1!
1%
#525510000000
0!
0%
#525515000000
1!
1%
#525520000000
0!
0%
#525525000000
1!
1%
#525530000000
0!
0%
#525535000000
1!
1%
#525540000000
0!
0%
#525545000000
1!
1%
#525550000000
0!
0%
#525555000000
1!
1%
#525560000000
0!
0%
#525565000000
1!
1%
#525570000000
0!
0%
#525575000000
1!
1%
#525580000000
0!
0%
#525585000000
1!
1%
#525590000000
0!
0%
#525595000000
1!
1%
#525600000000
0!
0%
#525605000000
1!
1%
#525610000000
0!
0%
#525615000000
1!
1%
#525620000000
0!
0%
#525625000000
1!
1%
#525630000000
0!
0%
#525635000000
1!
1%
#525640000000
0!
0%
#525645000000
1!
1%
#525650000000
0!
0%
#525655000000
1!
1%
#525660000000
0!
0%
#525665000000
1!
1%
#525670000000
0!
0%
#525675000000
1!
1%
#525680000000
0!
0%
#525685000000
1!
1%
#525690000000
0!
0%
#525695000000
1!
1%
#525700000000
0!
0%
#525705000000
1!
1%
#525710000000
0!
0%
#525715000000
1!
1%
#525720000000
0!
0%
#525725000000
1!
1%
#525730000000
0!
0%
#525735000000
1!
1%
#525740000000
0!
0%
#525745000000
1!
1%
#525750000000
0!
0%
#525755000000
1!
1%
#525760000000
0!
0%
#525765000000
1!
1%
#525770000000
0!
0%
#525775000000
1!
1%
#525780000000
0!
0%
#525785000000
1!
1%
#525790000000
0!
0%
#525795000000
1!
1%
#525800000000
0!
0%
#525805000000
1!
1%
#525810000000
0!
0%
#525815000000
1!
1%
#525820000000
0!
0%
#525825000000
1!
1%
#525830000000
0!
0%
#525835000000
1!
1%
#525840000000
0!
0%
#525845000000
1!
1%
#525850000000
0!
0%
#525855000000
1!
1%
#525860000000
0!
0%
#525865000000
1!
1%
#525870000000
0!
0%
#525875000000
1!
1%
#525880000000
0!
0%
#525885000000
1!
1%
#525890000000
0!
0%
#525895000000
1!
1%
#525900000000
0!
0%
#525905000000
1!
1%
#525910000000
0!
0%
#525915000000
1!
1%
#525920000000
0!
0%
#525925000000
1!
1%
#525930000000
0!
0%
#525935000000
1!
1%
#525940000000
0!
0%
#525945000000
1!
1%
#525950000000
0!
0%
#525955000000
1!
1%
#525960000000
0!
0%
#525965000000
1!
1%
#525970000000
0!
0%
#525975000000
1!
1%
#525980000000
0!
0%
#525985000000
1!
1%
#525990000000
0!
0%
#525995000000
1!
1%
#526000000000
0!
0%
#526005000000
1!
1%
#526010000000
0!
0%
#526015000000
1!
1%
#526020000000
0!
0%
#526025000000
1!
1%
#526030000000
0!
0%
#526035000000
1!
1%
#526040000000
0!
0%
#526045000000
1!
1%
#526050000000
0!
0%
#526055000000
1!
1%
#526060000000
0!
0%
#526065000000
1!
1%
#526070000000
0!
0%
#526075000000
1!
1%
#526080000000
0!
0%
#526085000000
1!
1%
#526090000000
0!
0%
#526095000000
1!
1%
#526100000000
0!
0%
#526105000000
1!
1%
#526110000000
0!
0%
#526115000000
1!
1%
#526120000000
0!
0%
#526125000000
1!
1%
#526130000000
0!
0%
#526135000000
1!
1%
#526140000000
0!
0%
#526145000000
1!
1%
#526150000000
0!
0%
#526155000000
1!
1%
#526160000000
0!
0%
#526165000000
1!
1%
#526170000000
0!
0%
#526175000000
1!
1%
#526180000000
0!
0%
#526185000000
1!
1%
#526190000000
0!
0%
#526195000000
1!
1%
#526200000000
0!
0%
#526205000000
1!
1%
#526210000000
0!
0%
#526215000000
1!
1%
#526220000000
0!
0%
#526225000000
1!
1%
#526230000000
0!
0%
#526235000000
1!
1%
#526240000000
0!
0%
#526245000000
1!
1%
#526250000000
0!
0%
#526255000000
1!
1%
#526260000000
0!
0%
#526265000000
1!
1%
#526270000000
0!
0%
#526275000000
1!
1%
#526280000000
0!
0%
#526285000000
1!
1%
#526290000000
0!
0%
#526295000000
1!
1%
#526300000000
0!
0%
#526305000000
1!
1%
#526310000000
0!
0%
#526315000000
1!
1%
#526320000000
0!
0%
#526325000000
1!
1%
#526330000000
0!
0%
#526335000000
1!
1%
#526340000000
0!
0%
#526345000000
1!
1%
#526350000000
0!
0%
#526355000000
1!
1%
#526360000000
0!
0%
#526365000000
1!
1%
#526370000000
0!
0%
#526375000000
1!
1%
#526380000000
0!
0%
#526385000000
1!
1%
#526390000000
0!
0%
#526395000000
1!
1%
#526400000000
0!
0%
#526405000000
1!
1%
#526410000000
0!
0%
#526415000000
1!
1%
#526420000000
0!
0%
#526425000000
1!
1%
#526430000000
0!
0%
#526435000000
1!
1%
#526440000000
0!
0%
#526445000000
1!
1%
#526450000000
0!
0%
#526455000000
1!
1%
#526460000000
0!
0%
#526465000000
1!
1%
#526470000000
0!
0%
#526475000000
1!
1%
#526480000000
0!
0%
#526485000000
1!
1%
#526490000000
0!
0%
#526495000000
1!
1%
#526500000000
0!
0%
#526505000000
1!
1%
#526510000000
0!
0%
#526515000000
1!
1%
#526520000000
0!
0%
#526525000000
1!
1%
#526530000000
0!
0%
#526535000000
1!
1%
#526540000000
0!
0%
#526545000000
1!
1%
#526550000000
0!
0%
#526555000000
1!
1%
#526560000000
0!
0%
#526565000000
1!
1%
#526570000000
0!
0%
#526575000000
1!
1%
#526580000000
0!
0%
#526585000000
1!
1%
#526590000000
0!
0%
#526595000000
1!
1%
#526600000000
0!
0%
#526605000000
1!
1%
#526610000000
0!
0%
#526615000000
1!
1%
#526620000000
0!
0%
#526625000000
1!
1%
#526630000000
0!
0%
#526635000000
1!
1%
#526640000000
0!
0%
#526645000000
1!
1%
#526650000000
0!
0%
#526655000000
1!
1%
#526660000000
0!
0%
#526665000000
1!
1%
#526670000000
0!
0%
#526675000000
1!
1%
#526680000000
0!
0%
#526685000000
1!
1%
#526690000000
0!
0%
#526695000000
1!
1%
#526700000000
0!
0%
#526705000000
1!
1%
#526710000000
0!
0%
#526715000000
1!
1%
#526720000000
0!
0%
#526725000000
1!
1%
#526730000000
0!
0%
#526735000000
1!
1%
#526740000000
0!
0%
#526745000000
1!
1%
#526750000000
0!
0%
#526755000000
1!
1%
#526760000000
0!
0%
#526765000000
1!
1%
#526770000000
0!
0%
#526775000000
1!
1%
#526780000000
0!
0%
#526785000000
1!
1%
#526790000000
0!
0%
#526795000000
1!
1%
#526800000000
0!
0%
#526805000000
1!
1%
#526810000000
0!
0%
#526815000000
1!
1%
#526820000000
0!
0%
#526825000000
1!
1%
#526830000000
0!
0%
#526835000000
1!
1%
#526840000000
0!
0%
#526845000000
1!
1%
#526850000000
0!
0%
#526855000000
1!
1%
#526860000000
0!
0%
#526865000000
1!
1%
#526870000000
0!
0%
#526875000000
1!
1%
#526880000000
0!
0%
#526885000000
1!
1%
#526890000000
0!
0%
#526895000000
1!
1%
#526900000000
0!
0%
#526905000000
1!
1%
#526910000000
0!
0%
#526915000000
1!
1%
#526920000000
0!
0%
#526925000000
1!
1%
#526930000000
0!
0%
#526935000000
1!
1%
#526940000000
0!
0%
#526945000000
1!
1%
#526950000000
0!
0%
#526955000000
1!
1%
#526960000000
0!
0%
#526965000000
1!
1%
#526970000000
0!
0%
#526975000000
1!
1%
#526980000000
0!
0%
#526985000000
1!
1%
#526990000000
0!
0%
#526995000000
1!
1%
#527000000000
0!
0%
#527005000000
1!
1%
#527010000000
0!
0%
#527015000000
1!
1%
#527020000000
0!
0%
#527025000000
1!
1%
#527030000000
0!
0%
#527035000000
1!
1%
#527040000000
0!
0%
#527045000000
1!
1%
#527050000000
0!
0%
#527055000000
1!
1%
#527060000000
0!
0%
#527065000000
1!
1%
#527070000000
0!
0%
#527075000000
1!
1%
#527080000000
0!
0%
#527085000000
1!
1%
#527090000000
0!
0%
#527095000000
1!
1%
#527100000000
0!
0%
#527105000000
1!
1%
#527110000000
0!
0%
#527115000000
1!
1%
#527120000000
0!
0%
#527125000000
1!
1%
#527130000000
0!
0%
#527135000000
1!
1%
#527140000000
0!
0%
#527145000000
1!
1%
#527150000000
0!
0%
#527155000000
1!
1%
#527160000000
0!
0%
#527165000000
1!
1%
#527170000000
0!
0%
#527175000000
1!
1%
#527180000000
0!
0%
#527185000000
1!
1%
#527190000000
0!
0%
#527195000000
1!
1%
#527200000000
0!
0%
#527205000000
1!
1%
#527210000000
0!
0%
#527215000000
1!
1%
#527220000000
0!
0%
#527225000000
1!
1%
#527230000000
0!
0%
#527235000000
1!
1%
#527240000000
0!
0%
#527245000000
1!
1%
#527250000000
0!
0%
#527255000000
1!
1%
#527260000000
0!
0%
#527265000000
1!
1%
#527270000000
0!
0%
#527275000000
1!
1%
#527280000000
0!
0%
#527285000000
1!
1%
#527290000000
0!
0%
#527295000000
1!
1%
#527300000000
0!
0%
#527305000000
1!
1%
#527310000000
0!
0%
#527315000000
1!
1%
#527320000000
0!
0%
#527325000000
1!
1%
#527330000000
0!
0%
#527335000000
1!
1%
#527340000000
0!
0%
#527345000000
1!
1%
#527350000000
0!
0%
#527355000000
1!
1%
#527360000000
0!
0%
#527365000000
1!
1%
#527370000000
0!
0%
#527375000000
1!
1%
#527380000000
0!
0%
#527385000000
1!
1%
#527390000000
0!
0%
#527395000000
1!
1%
#527400000000
0!
0%
#527405000000
1!
1%
#527410000000
0!
0%
#527415000000
1!
1%
#527420000000
0!
0%
#527425000000
1!
1%
#527430000000
0!
0%
#527435000000
1!
1%
#527440000000
0!
0%
#527445000000
1!
1%
#527450000000
0!
0%
#527455000000
1!
1%
#527460000000
0!
0%
#527465000000
1!
1%
#527470000000
0!
0%
#527475000000
1!
1%
#527480000000
0!
0%
#527485000000
1!
1%
#527490000000
0!
0%
#527495000000
1!
1%
#527500000000
0!
0%
#527505000000
1!
1%
#527510000000
0!
0%
#527515000000
1!
1%
#527520000000
0!
0%
#527525000000
1!
1%
#527530000000
0!
0%
#527535000000
1!
1%
#527540000000
0!
0%
#527545000000
1!
1%
#527550000000
0!
0%
#527555000000
1!
1%
#527560000000
0!
0%
#527565000000
1!
1%
#527570000000
0!
0%
#527575000000
1!
1%
#527580000000
0!
0%
#527585000000
1!
1%
#527590000000
0!
0%
#527595000000
1!
1%
#527600000000
0!
0%
#527605000000
1!
1%
#527610000000
0!
0%
#527615000000
1!
1%
#527620000000
0!
0%
#527625000000
1!
1%
#527630000000
0!
0%
#527635000000
1!
1%
#527640000000
0!
0%
#527645000000
1!
1%
#527650000000
0!
0%
#527655000000
1!
1%
#527660000000
0!
0%
#527665000000
1!
1%
#527670000000
0!
0%
#527675000000
1!
1%
#527680000000
0!
0%
#527685000000
1!
1%
#527690000000
0!
0%
#527695000000
1!
1%
#527700000000
0!
0%
#527705000000
1!
1%
#527710000000
0!
0%
#527715000000
1!
1%
#527720000000
0!
0%
#527725000000
1!
1%
#527730000000
0!
0%
#527735000000
1!
1%
#527740000000
0!
0%
#527745000000
1!
1%
#527750000000
0!
0%
#527755000000
1!
1%
#527760000000
0!
0%
#527765000000
1!
1%
#527770000000
0!
0%
#527775000000
1!
1%
#527780000000
0!
0%
#527785000000
1!
1%
#527790000000
0!
0%
#527795000000
1!
1%
#527800000000
0!
0%
#527805000000
1!
1%
#527810000000
0!
0%
#527815000000
1!
1%
#527820000000
0!
0%
#527825000000
1!
1%
#527830000000
0!
0%
#527835000000
1!
1%
#527840000000
0!
0%
#527845000000
1!
1%
#527850000000
0!
0%
#527855000000
1!
1%
#527860000000
0!
0%
#527865000000
1!
1%
#527870000000
0!
0%
#527875000000
1!
1%
#527880000000
0!
0%
#527885000000
1!
1%
#527890000000
0!
0%
#527895000000
1!
1%
#527900000000
0!
0%
#527905000000
1!
1%
#527910000000
0!
0%
#527915000000
1!
1%
#527920000000
0!
0%
#527925000000
1!
1%
#527930000000
0!
0%
#527935000000
1!
1%
#527940000000
0!
0%
#527945000000
1!
1%
#527950000000
0!
0%
#527955000000
1!
1%
#527960000000
0!
0%
#527965000000
1!
1%
#527970000000
0!
0%
#527975000000
1!
1%
#527980000000
0!
0%
#527985000000
1!
1%
#527990000000
0!
0%
#527995000000
1!
1%
#528000000000
0!
0%
#528005000000
1!
1%
#528010000000
0!
0%
#528015000000
1!
1%
#528020000000
0!
0%
#528025000000
1!
1%
#528030000000
0!
0%
#528035000000
1!
1%
#528040000000
0!
0%
#528045000000
1!
1%
#528050000000
0!
0%
#528055000000
1!
1%
#528060000000
0!
0%
#528065000000
1!
1%
#528070000000
0!
0%
#528075000000
1!
1%
#528080000000
0!
0%
#528085000000
1!
1%
#528090000000
0!
0%
#528095000000
1!
1%
#528100000000
0!
0%
#528105000000
1!
1%
#528110000000
0!
0%
#528115000000
1!
1%
#528120000000
0!
0%
#528125000000
1!
1%
#528130000000
0!
0%
#528135000000
1!
1%
#528140000000
0!
0%
#528145000000
1!
1%
#528150000000
0!
0%
#528155000000
1!
1%
#528160000000
0!
0%
#528165000000
1!
1%
#528170000000
0!
0%
#528175000000
1!
1%
#528180000000
0!
0%
#528185000000
1!
1%
#528190000000
0!
0%
#528195000000
1!
1%
#528200000000
0!
0%
#528205000000
1!
1%
#528210000000
0!
0%
#528215000000
1!
1%
#528220000000
0!
0%
#528225000000
1!
1%
#528230000000
0!
0%
#528235000000
1!
1%
#528240000000
0!
0%
#528245000000
1!
1%
#528250000000
0!
0%
#528255000000
1!
1%
#528260000000
0!
0%
#528265000000
1!
1%
#528270000000
0!
0%
#528275000000
1!
1%
#528280000000
0!
0%
#528285000000
1!
1%
#528290000000
0!
0%
#528295000000
1!
1%
#528300000000
0!
0%
#528305000000
1!
1%
#528310000000
0!
0%
#528315000000
1!
1%
#528320000000
0!
0%
#528325000000
1!
1%
#528330000000
0!
0%
#528335000000
1!
1%
#528340000000
0!
0%
#528345000000
1!
1%
#528350000000
0!
0%
#528355000000
1!
1%
#528360000000
0!
0%
#528365000000
1!
1%
#528370000000
0!
0%
#528375000000
1!
1%
#528380000000
0!
0%
#528385000000
1!
1%
#528390000000
0!
0%
#528395000000
1!
1%
#528400000000
0!
0%
#528405000000
1!
1%
#528410000000
0!
0%
#528415000000
1!
1%
#528420000000
0!
0%
#528425000000
1!
1%
#528430000000
0!
0%
#528435000000
1!
1%
#528440000000
0!
0%
#528445000000
1!
1%
#528450000000
0!
0%
#528455000000
1!
1%
#528460000000
0!
0%
#528465000000
1!
1%
#528470000000
0!
0%
#528475000000
1!
1%
#528480000000
0!
0%
#528485000000
1!
1%
#528490000000
0!
0%
#528495000000
1!
1%
#528500000000
0!
0%
#528505000000
1!
1%
#528510000000
0!
0%
#528515000000
1!
1%
#528520000000
0!
0%
#528525000000
1!
1%
#528530000000
0!
0%
#528535000000
1!
1%
#528540000000
0!
0%
#528545000000
1!
1%
#528550000000
0!
0%
#528555000000
1!
1%
#528560000000
0!
0%
#528565000000
1!
1%
#528570000000
0!
0%
#528575000000
1!
1%
#528580000000
0!
0%
#528585000000
1!
1%
#528590000000
0!
0%
#528595000000
1!
1%
#528600000000
0!
0%
#528605000000
1!
1%
#528610000000
0!
0%
#528615000000
1!
1%
#528620000000
0!
0%
#528625000000
1!
1%
#528630000000
0!
0%
#528635000000
1!
1%
#528640000000
0!
0%
#528645000000
1!
1%
#528650000000
0!
0%
#528655000000
1!
1%
#528660000000
0!
0%
#528665000000
1!
1%
#528670000000
0!
0%
#528675000000
1!
1%
#528680000000
0!
0%
#528685000000
1!
1%
#528690000000
0!
0%
#528695000000
1!
1%
#528700000000
0!
0%
#528705000000
1!
1%
#528710000000
0!
0%
#528715000000
1!
1%
#528720000000
0!
0%
#528725000000
1!
1%
#528730000000
0!
0%
#528735000000
1!
1%
#528740000000
0!
0%
#528745000000
1!
1%
#528750000000
0!
0%
#528755000000
1!
1%
#528760000000
0!
0%
#528765000000
1!
1%
#528770000000
0!
0%
#528775000000
1!
1%
#528780000000
0!
0%
#528785000000
1!
1%
#528790000000
0!
0%
#528795000000
1!
1%
#528800000000
0!
0%
#528805000000
1!
1%
#528810000000
0!
0%
#528815000000
1!
1%
#528820000000
0!
0%
#528825000000
1!
1%
#528830000000
0!
0%
#528835000000
1!
1%
#528840000000
0!
0%
#528845000000
1!
1%
#528850000000
0!
0%
#528855000000
1!
1%
#528860000000
0!
0%
#528865000000
1!
1%
#528870000000
0!
0%
#528875000000
1!
1%
#528880000000
0!
0%
#528885000000
1!
1%
#528890000000
0!
0%
#528895000000
1!
1%
#528900000000
0!
0%
#528905000000
1!
1%
#528910000000
0!
0%
#528915000000
1!
1%
#528920000000
0!
0%
#528925000000
1!
1%
#528930000000
0!
0%
#528935000000
1!
1%
#528940000000
0!
0%
#528945000000
1!
1%
#528950000000
0!
0%
#528955000000
1!
1%
#528960000000
0!
0%
#528965000000
1!
1%
#528970000000
0!
0%
#528975000000
1!
1%
#528980000000
0!
0%
#528985000000
1!
1%
#528990000000
0!
0%
#528995000000
1!
1%
#529000000000
0!
0%
#529005000000
1!
1%
#529010000000
0!
0%
#529015000000
1!
1%
#529020000000
0!
0%
#529025000000
1!
1%
#529030000000
0!
0%
#529035000000
1!
1%
#529040000000
0!
0%
#529045000000
1!
1%
#529050000000
0!
0%
#529055000000
1!
1%
#529060000000
0!
0%
#529065000000
1!
1%
#529070000000
0!
0%
#529075000000
1!
1%
#529080000000
0!
0%
#529085000000
1!
1%
#529090000000
0!
0%
#529095000000
1!
1%
#529100000000
0!
0%
#529105000000
1!
1%
#529110000000
0!
0%
#529115000000
1!
1%
#529120000000
0!
0%
#529125000000
1!
1%
#529130000000
0!
0%
#529135000000
1!
1%
#529140000000
0!
0%
#529145000000
1!
1%
#529150000000
0!
0%
#529155000000
1!
1%
#529160000000
0!
0%
#529165000000
1!
1%
#529170000000
0!
0%
#529175000000
1!
1%
#529180000000
0!
0%
#529185000000
1!
1%
#529190000000
0!
0%
#529195000000
1!
1%
#529200000000
0!
0%
#529205000000
1!
1%
#529210000000
0!
0%
#529215000000
1!
1%
#529220000000
0!
0%
#529225000000
1!
1%
#529230000000
0!
0%
#529235000000
1!
1%
#529240000000
0!
0%
#529245000000
1!
1%
#529250000000
0!
0%
#529255000000
1!
1%
#529260000000
0!
0%
#529265000000
1!
1%
#529270000000
0!
0%
#529275000000
1!
1%
#529280000000
0!
0%
#529285000000
1!
1%
#529290000000
0!
0%
#529295000000
1!
1%
#529300000000
0!
0%
#529305000000
1!
1%
#529310000000
0!
0%
#529315000000
1!
1%
#529320000000
0!
0%
#529325000000
1!
1%
#529330000000
0!
0%
#529335000000
1!
1%
#529340000000
0!
0%
#529345000000
1!
1%
#529350000000
0!
0%
#529355000000
1!
1%
#529360000000
0!
0%
#529365000000
1!
1%
#529370000000
0!
0%
#529375000000
1!
1%
#529380000000
0!
0%
#529385000000
1!
1%
#529390000000
0!
0%
#529395000000
1!
1%
#529400000000
0!
0%
#529405000000
1!
1%
#529410000000
0!
0%
#529415000000
1!
1%
#529420000000
0!
0%
#529425000000
1!
1%
#529430000000
0!
0%
#529435000000
1!
1%
#529440000000
0!
0%
#529445000000
1!
1%
#529450000000
0!
0%
#529455000000
1!
1%
#529460000000
0!
0%
#529465000000
1!
1%
#529470000000
0!
0%
#529475000000
1!
1%
#529480000000
0!
0%
#529485000000
1!
1%
#529490000000
0!
0%
#529495000000
1!
1%
#529500000000
0!
0%
#529505000000
1!
1%
#529510000000
0!
0%
#529515000000
1!
1%
#529520000000
0!
0%
#529525000000
1!
1%
#529530000000
0!
0%
#529535000000
1!
1%
#529540000000
0!
0%
#529545000000
1!
1%
#529550000000
0!
0%
#529555000000
1!
1%
#529560000000
0!
0%
#529565000000
1!
1%
#529570000000
0!
0%
#529575000000
1!
1%
#529580000000
0!
0%
#529585000000
1!
1%
#529590000000
0!
0%
#529595000000
1!
1%
#529600000000
0!
0%
#529605000000
1!
1%
#529610000000
0!
0%
#529615000000
1!
1%
#529620000000
0!
0%
#529625000000
1!
1%
#529630000000
0!
0%
#529635000000
1!
1%
#529640000000
0!
0%
#529645000000
1!
1%
#529650000000
0!
0%
#529655000000
1!
1%
#529660000000
0!
0%
#529665000000
1!
1%
#529670000000
0!
0%
#529675000000
1!
1%
#529680000000
0!
0%
#529685000000
1!
1%
#529690000000
0!
0%
#529695000000
1!
1%
#529700000000
0!
0%
#529705000000
1!
1%
#529710000000
0!
0%
#529715000000
1!
1%
#529720000000
0!
0%
#529725000000
1!
1%
#529730000000
0!
0%
#529735000000
1!
1%
#529740000000
0!
0%
#529745000000
1!
1%
#529750000000
0!
0%
#529755000000
1!
1%
#529760000000
0!
0%
#529765000000
1!
1%
#529770000000
0!
0%
#529775000000
1!
1%
#529780000000
0!
0%
#529785000000
1!
1%
#529790000000
0!
0%
#529795000000
1!
1%
#529800000000
0!
0%
#529805000000
1!
1%
#529810000000
0!
0%
#529815000000
1!
1%
#529820000000
0!
0%
#529825000000
1!
1%
#529830000000
0!
0%
#529835000000
1!
1%
#529840000000
0!
0%
#529845000000
1!
1%
#529850000000
0!
0%
#529855000000
1!
1%
#529860000000
0!
0%
#529865000000
1!
1%
#529870000000
0!
0%
#529875000000
1!
1%
#529880000000
0!
0%
#529885000000
1!
1%
#529890000000
0!
0%
#529895000000
1!
1%
#529900000000
0!
0%
#529905000000
1!
1%
#529910000000
0!
0%
#529915000000
1!
1%
#529920000000
0!
0%
#529925000000
1!
1%
#529930000000
0!
0%
#529935000000
1!
1%
#529940000000
0!
0%
#529945000000
1!
1%
#529950000000
0!
0%
#529955000000
1!
1%
#529960000000
0!
0%
#529965000000
1!
1%
#529970000000
0!
0%
#529975000000
1!
1%
#529980000000
0!
0%
#529985000000
1!
1%
#529990000000
0!
0%
#529995000000
1!
1%
#530000000000
0!
0%
#530005000000
1!
1%
#530010000000
0!
0%
#530015000000
1!
1%
#530020000000
0!
0%
#530025000000
1!
1%
#530030000000
0!
0%
#530035000000
1!
1%
#530040000000
0!
0%
#530045000000
1!
1%
#530050000000
0!
0%
#530055000000
1!
1%
#530060000000
0!
0%
#530065000000
1!
1%
#530070000000
0!
0%
#530075000000
1!
1%
#530080000000
0!
0%
#530085000000
1!
1%
#530090000000
0!
0%
#530095000000
1!
1%
#530100000000
0!
0%
#530105000000
1!
1%
#530110000000
0!
0%
#530115000000
1!
1%
#530120000000
0!
0%
#530125000000
1!
1%
#530130000000
0!
0%
#530135000000
1!
1%
#530140000000
0!
0%
#530145000000
1!
1%
#530150000000
0!
0%
#530155000000
1!
1%
#530160000000
0!
0%
#530165000000
1!
1%
#530170000000
0!
0%
#530175000000
1!
1%
#530180000000
0!
0%
#530185000000
1!
1%
#530190000000
0!
0%
#530195000000
1!
1%
#530200000000
0!
0%
#530205000000
1!
1%
#530210000000
0!
0%
#530215000000
1!
1%
#530220000000
0!
0%
#530225000000
1!
1%
#530230000000
0!
0%
#530235000000
1!
1%
#530240000000
0!
0%
#530245000000
1!
1%
#530250000000
0!
0%
#530255000000
1!
1%
#530260000000
0!
0%
#530265000000
1!
1%
#530270000000
0!
0%
#530275000000
1!
1%
#530280000000
0!
0%
#530285000000
1!
1%
#530290000000
0!
0%
#530295000000
1!
1%
#530300000000
0!
0%
#530305000000
1!
1%
#530310000000
0!
0%
#530315000000
1!
1%
#530320000000
0!
0%
#530325000000
1!
1%
#530330000000
0!
0%
#530335000000
1!
1%
#530340000000
0!
0%
#530345000000
1!
1%
#530350000000
0!
0%
#530355000000
1!
1%
#530360000000
0!
0%
#530365000000
1!
1%
#530370000000
0!
0%
#530375000000
1!
1%
#530380000000
0!
0%
#530385000000
1!
1%
#530390000000
0!
0%
#530395000000
1!
1%
#530400000000
0!
0%
#530405000000
1!
1%
#530410000000
0!
0%
#530415000000
1!
1%
#530420000000
0!
0%
#530425000000
1!
1%
#530430000000
0!
0%
#530435000000
1!
1%
#530440000000
0!
0%
#530445000000
1!
1%
#530450000000
0!
0%
#530455000000
1!
1%
#530460000000
0!
0%
#530465000000
1!
1%
#530470000000
0!
0%
#530475000000
1!
1%
#530480000000
0!
0%
#530485000000
1!
1%
#530490000000
0!
0%
#530495000000
1!
1%
#530500000000
0!
0%
#530505000000
1!
1%
#530510000000
0!
0%
#530515000000
1!
1%
#530520000000
0!
0%
#530525000000
1!
1%
#530530000000
0!
0%
#530535000000
1!
1%
#530540000000
0!
0%
#530545000000
1!
1%
#530550000000
0!
0%
#530555000000
1!
1%
#530560000000
0!
0%
#530565000000
1!
1%
#530570000000
0!
0%
#530575000000
1!
1%
#530580000000
0!
0%
#530585000000
1!
1%
#530590000000
0!
0%
#530595000000
1!
1%
#530600000000
0!
0%
#530605000000
1!
1%
#530610000000
0!
0%
#530615000000
1!
1%
#530620000000
0!
0%
#530625000000
1!
1%
#530630000000
0!
0%
#530635000000
1!
1%
#530640000000
0!
0%
#530645000000
1!
1%
#530650000000
0!
0%
#530655000000
1!
1%
#530660000000
0!
0%
#530665000000
1!
1%
#530670000000
0!
0%
#530675000000
1!
1%
#530680000000
0!
0%
#530685000000
1!
1%
#530690000000
0!
0%
#530695000000
1!
1%
#530700000000
0!
0%
#530705000000
1!
1%
#530710000000
0!
0%
#530715000000
1!
1%
#530720000000
0!
0%
#530725000000
1!
1%
#530730000000
0!
0%
#530735000000
1!
1%
#530740000000
0!
0%
#530745000000
1!
1%
#530750000000
0!
0%
#530755000000
1!
1%
#530760000000
0!
0%
#530765000000
1!
1%
#530770000000
0!
0%
#530775000000
1!
1%
#530780000000
0!
0%
#530785000000
1!
1%
#530790000000
0!
0%
#530795000000
1!
1%
#530800000000
0!
0%
#530805000000
1!
1%
#530810000000
0!
0%
#530815000000
1!
1%
#530820000000
0!
0%
#530825000000
1!
1%
#530830000000
0!
0%
#530835000000
1!
1%
#530840000000
0!
0%
#530845000000
1!
1%
#530850000000
0!
0%
#530855000000
1!
1%
#530860000000
0!
0%
#530865000000
1!
1%
#530870000000
0!
0%
#530875000000
1!
1%
#530880000000
0!
0%
#530885000000
1!
1%
#530890000000
0!
0%
#530895000000
1!
1%
#530900000000
0!
0%
#530905000000
1!
1%
#530910000000
0!
0%
#530915000000
1!
1%
#530920000000
0!
0%
#530925000000
1!
1%
#530930000000
0!
0%
#530935000000
1!
1%
#530940000000
0!
0%
#530945000000
1!
1%
#530950000000
0!
0%
#530955000000
1!
1%
#530960000000
0!
0%
#530965000000
1!
1%
#530970000000
0!
0%
#530975000000
1!
1%
#530980000000
0!
0%
#530985000000
1!
1%
#530990000000
0!
0%
#530995000000
1!
1%
#531000000000
0!
0%
#531005000000
1!
1%
#531010000000
0!
0%
#531015000000
1!
1%
#531020000000
0!
0%
#531025000000
1!
1%
#531030000000
0!
0%
#531035000000
1!
1%
#531040000000
0!
0%
#531045000000
1!
1%
#531050000000
0!
0%
#531055000000
1!
1%
#531060000000
0!
0%
#531065000000
1!
1%
#531070000000
0!
0%
#531075000000
1!
1%
#531080000000
0!
0%
#531085000000
1!
1%
#531090000000
0!
0%
#531095000000
1!
1%
#531100000000
0!
0%
#531105000000
1!
1%
#531110000000
0!
0%
#531115000000
1!
1%
#531120000000
0!
0%
#531125000000
1!
1%
#531130000000
0!
0%
#531135000000
1!
1%
#531140000000
0!
0%
#531145000000
1!
1%
#531150000000
0!
0%
#531155000000
1!
1%
#531160000000
0!
0%
#531165000000
1!
1%
#531170000000
0!
0%
#531175000000
1!
1%
#531180000000
0!
0%
#531185000000
1!
1%
#531190000000
0!
0%
#531195000000
1!
1%
#531200000000
0!
0%
#531205000000
1!
1%
#531210000000
0!
0%
#531215000000
1!
1%
#531220000000
0!
0%
#531225000000
1!
1%
#531230000000
0!
0%
#531235000000
1!
1%
#531240000000
0!
0%
#531245000000
1!
1%
#531250000000
0!
0%
#531255000000
1!
1%
#531260000000
0!
0%
#531265000000
1!
1%
#531270000000
0!
0%
#531275000000
1!
1%
#531280000000
0!
0%
#531285000000
1!
1%
#531290000000
0!
0%
#531295000000
1!
1%
#531300000000
0!
0%
#531305000000
1!
1%
#531310000000
0!
0%
#531315000000
1!
1%
#531320000000
0!
0%
#531325000000
1!
1%
#531330000000
0!
0%
#531335000000
1!
1%
#531340000000
0!
0%
#531345000000
1!
1%
#531350000000
0!
0%
#531355000000
1!
1%
#531360000000
0!
0%
#531365000000
1!
1%
#531370000000
0!
0%
#531375000000
1!
1%
#531380000000
0!
0%
#531385000000
1!
1%
#531390000000
0!
0%
#531395000000
1!
1%
#531400000000
0!
0%
#531405000000
1!
1%
#531410000000
0!
0%
#531415000000
1!
1%
#531420000000
0!
0%
#531425000000
1!
1%
#531430000000
0!
0%
#531435000000
1!
1%
#531440000000
0!
0%
#531445000000
1!
1%
#531450000000
0!
0%
#531455000000
1!
1%
#531460000000
0!
0%
#531465000000
1!
1%
#531470000000
0!
0%
#531475000000
1!
1%
#531480000000
0!
0%
#531485000000
1!
1%
#531490000000
0!
0%
#531495000000
1!
1%
#531500000000
0!
0%
#531505000000
1!
1%
#531510000000
0!
0%
#531515000000
1!
1%
#531520000000
0!
0%
#531525000000
1!
1%
#531530000000
0!
0%
#531535000000
1!
1%
#531540000000
0!
0%
#531545000000
1!
1%
#531550000000
0!
0%
#531555000000
1!
1%
#531560000000
0!
0%
#531565000000
1!
1%
#531570000000
0!
0%
#531575000000
1!
1%
#531580000000
0!
0%
#531585000000
1!
1%
#531590000000
0!
0%
#531595000000
1!
1%
#531600000000
0!
0%
#531605000000
1!
1%
#531610000000
0!
0%
#531615000000
1!
1%
#531620000000
0!
0%
#531625000000
1!
1%
#531630000000
0!
0%
#531635000000
1!
1%
#531640000000
0!
0%
#531645000000
1!
1%
#531650000000
0!
0%
#531655000000
1!
1%
#531660000000
0!
0%
#531665000000
1!
1%
#531670000000
0!
0%
#531675000000
1!
1%
#531680000000
0!
0%
#531685000000
1!
1%
#531690000000
0!
0%
#531695000000
1!
1%
#531700000000
0!
0%
#531705000000
1!
1%
#531710000000
0!
0%
#531715000000
1!
1%
#531720000000
0!
0%
#531725000000
1!
1%
#531730000000
0!
0%
#531735000000
1!
1%
#531740000000
0!
0%
#531745000000
1!
1%
#531750000000
0!
0%
#531755000000
1!
1%
#531760000000
0!
0%
#531765000000
1!
1%
#531770000000
0!
0%
#531775000000
1!
1%
#531780000000
0!
0%
#531785000000
1!
1%
#531790000000
0!
0%
#531795000000
1!
1%
#531800000000
0!
0%
#531805000000
1!
1%
#531810000000
0!
0%
#531815000000
1!
1%
#531820000000
0!
0%
#531825000000
1!
1%
#531830000000
0!
0%
#531835000000
1!
1%
#531840000000
0!
0%
#531845000000
1!
1%
#531850000000
0!
0%
#531855000000
1!
1%
#531860000000
0!
0%
#531865000000
1!
1%
#531870000000
0!
0%
#531875000000
1!
1%
#531880000000
0!
0%
#531885000000
1!
1%
#531890000000
0!
0%
#531895000000
1!
1%
#531900000000
0!
0%
#531905000000
1!
1%
#531910000000
0!
0%
#531915000000
1!
1%
#531920000000
0!
0%
#531925000000
1!
1%
#531930000000
0!
0%
#531935000000
1!
1%
#531940000000
0!
0%
#531945000000
1!
1%
#531950000000
0!
0%
#531955000000
1!
1%
#531960000000
0!
0%
#531965000000
1!
1%
#531970000000
0!
0%
#531975000000
1!
1%
#531980000000
0!
0%
#531985000000
1!
1%
#531990000000
0!
0%
#531995000000
1!
1%
#532000000000
0!
0%
#532005000000
1!
1%
#532010000000
0!
0%
#532015000000
1!
1%
#532020000000
0!
0%
#532025000000
1!
1%
#532030000000
0!
0%
#532035000000
1!
1%
#532040000000
0!
0%
#532045000000
1!
1%
#532050000000
0!
0%
#532055000000
1!
1%
#532060000000
0!
0%
#532065000000
1!
1%
#532070000000
0!
0%
#532075000000
1!
1%
#532080000000
0!
0%
#532085000000
1!
1%
#532090000000
0!
0%
#532095000000
1!
1%
#532100000000
0!
0%
#532105000000
1!
1%
#532110000000
0!
0%
#532115000000
1!
1%
#532120000000
0!
0%
#532125000000
1!
1%
#532130000000
0!
0%
#532135000000
1!
1%
#532140000000
0!
0%
#532145000000
1!
1%
#532150000000
0!
0%
#532155000000
1!
1%
#532160000000
0!
0%
#532165000000
1!
1%
#532170000000
0!
0%
#532175000000
1!
1%
#532180000000
0!
0%
#532185000000
1!
1%
#532190000000
0!
0%
#532195000000
1!
1%
#532200000000
0!
0%
#532205000000
1!
1%
#532210000000
0!
0%
#532215000000
1!
1%
#532220000000
0!
0%
#532225000000
1!
1%
#532230000000
0!
0%
#532235000000
1!
1%
#532240000000
0!
0%
#532245000000
1!
1%
#532250000000
0!
0%
#532255000000
1!
1%
#532260000000
0!
0%
#532265000000
1!
1%
#532270000000
0!
0%
#532275000000
1!
1%
#532280000000
0!
0%
#532285000000
1!
1%
#532290000000
0!
0%
#532295000000
1!
1%
#532300000000
0!
0%
#532305000000
1!
1%
#532310000000
0!
0%
#532315000000
1!
1%
#532320000000
0!
0%
#532325000000
1!
1%
#532330000000
0!
0%
#532335000000
1!
1%
#532340000000
0!
0%
#532345000000
1!
1%
#532350000000
0!
0%
#532355000000
1!
1%
#532360000000
0!
0%
#532365000000
1!
1%
#532370000000
0!
0%
#532375000000
1!
1%
#532380000000
0!
0%
#532385000000
1!
1%
#532390000000
0!
0%
#532395000000
1!
1%
#532400000000
0!
0%
#532405000000
1!
1%
#532410000000
0!
0%
#532415000000
1!
1%
#532420000000
0!
0%
#532425000000
1!
1%
#532430000000
0!
0%
#532435000000
1!
1%
#532440000000
0!
0%
#532445000000
1!
1%
#532450000000
0!
0%
#532455000000
1!
1%
#532460000000
0!
0%
#532465000000
1!
1%
#532470000000
0!
0%
#532475000000
1!
1%
#532480000000
0!
0%
#532485000000
1!
1%
#532490000000
0!
0%
#532495000000
1!
1%
#532500000000
0!
0%
#532505000000
1!
1%
#532510000000
0!
0%
#532515000000
1!
1%
#532520000000
0!
0%
#532525000000
1!
1%
#532530000000
0!
0%
#532535000000
1!
1%
#532540000000
0!
0%
#532545000000
1!
1%
#532550000000
0!
0%
#532555000000
1!
1%
#532560000000
0!
0%
#532565000000
1!
1%
#532570000000
0!
0%
#532575000000
1!
1%
#532580000000
0!
0%
#532585000000
1!
1%
#532590000000
0!
0%
#532595000000
1!
1%
#532600000000
0!
0%
#532605000000
1!
1%
#532610000000
0!
0%
#532615000000
1!
1%
#532620000000
0!
0%
#532625000000
1!
1%
#532630000000
0!
0%
#532635000000
1!
1%
#532640000000
0!
0%
#532645000000
1!
1%
#532650000000
0!
0%
#532655000000
1!
1%
#532660000000
0!
0%
#532665000000
1!
1%
#532670000000
0!
0%
#532675000000
1!
1%
#532680000000
0!
0%
#532685000000
1!
1%
#532690000000
0!
0%
#532695000000
1!
1%
#532700000000
0!
0%
#532705000000
1!
1%
#532710000000
0!
0%
#532715000000
1!
1%
#532720000000
0!
0%
#532725000000
1!
1%
#532730000000
0!
0%
#532735000000
1!
1%
#532740000000
0!
0%
#532745000000
1!
1%
#532750000000
0!
0%
#532755000000
1!
1%
#532760000000
0!
0%
#532765000000
1!
1%
#532770000000
0!
0%
#532775000000
1!
1%
#532780000000
0!
0%
#532785000000
1!
1%
#532790000000
0!
0%
#532795000000
1!
1%
#532800000000
0!
0%
#532805000000
1!
1%
#532810000000
0!
0%
#532815000000
1!
1%
#532820000000
0!
0%
#532825000000
1!
1%
#532830000000
0!
0%
#532835000000
1!
1%
#532840000000
0!
0%
#532845000000
1!
1%
#532850000000
0!
0%
#532855000000
1!
1%
#532860000000
0!
0%
#532865000000
1!
1%
#532870000000
0!
0%
#532875000000
1!
1%
#532880000000
0!
0%
#532885000000
1!
1%
#532890000000
0!
0%
#532895000000
1!
1%
#532900000000
0!
0%
#532905000000
1!
1%
#532910000000
0!
0%
#532915000000
1!
1%
#532920000000
0!
0%
#532925000000
1!
1%
#532930000000
0!
0%
#532935000000
1!
1%
#532940000000
0!
0%
#532945000000
1!
1%
#532950000000
0!
0%
#532955000000
1!
1%
#532960000000
0!
0%
#532965000000
1!
1%
#532970000000
0!
0%
#532975000000
1!
1%
#532980000000
0!
0%
#532985000000
1!
1%
#532990000000
0!
0%
#532995000000
1!
1%
#533000000000
0!
0%
#533005000000
1!
1%
#533010000000
0!
0%
#533015000000
1!
1%
#533020000000
0!
0%
#533025000000
1!
1%
#533030000000
0!
0%
#533035000000
1!
1%
#533040000000
0!
0%
#533045000000
1!
1%
#533050000000
0!
0%
#533055000000
1!
1%
#533060000000
0!
0%
#533065000000
1!
1%
#533070000000
0!
0%
#533075000000
1!
1%
#533080000000
0!
0%
#533085000000
1!
1%
#533090000000
0!
0%
#533095000000
1!
1%
#533100000000
0!
0%
#533105000000
1!
1%
#533110000000
0!
0%
#533115000000
1!
1%
#533120000000
0!
0%
#533125000000
1!
1%
#533130000000
0!
0%
#533135000000
1!
1%
#533140000000
0!
0%
#533145000000
1!
1%
#533150000000
0!
0%
#533155000000
1!
1%
#533160000000
0!
0%
#533165000000
1!
1%
#533170000000
0!
0%
#533175000000
1!
1%
#533180000000
0!
0%
#533185000000
1!
1%
#533190000000
0!
0%
#533195000000
1!
1%
#533200000000
0!
0%
#533205000000
1!
1%
#533210000000
0!
0%
#533215000000
1!
1%
#533220000000
0!
0%
#533225000000
1!
1%
#533230000000
0!
0%
#533235000000
1!
1%
#533240000000
0!
0%
#533245000000
1!
1%
#533250000000
0!
0%
#533255000000
1!
1%
#533260000000
0!
0%
#533265000000
1!
1%
#533270000000
0!
0%
#533275000000
1!
1%
#533280000000
0!
0%
#533285000000
1!
1%
#533290000000
0!
0%
#533295000000
1!
1%
#533300000000
0!
0%
#533305000000
1!
1%
#533310000000
0!
0%
#533315000000
1!
1%
#533320000000
0!
0%
#533325000000
1!
1%
#533330000000
0!
0%
#533335000000
1!
1%
#533340000000
0!
0%
#533345000000
1!
1%
#533350000000
0!
0%
#533355000000
1!
1%
#533360000000
0!
0%
#533365000000
1!
1%
#533370000000
0!
0%
#533375000000
1!
1%
#533380000000
0!
0%
#533385000000
1!
1%
#533390000000
0!
0%
#533395000000
1!
1%
#533400000000
0!
0%
#533405000000
1!
1%
#533410000000
0!
0%
#533415000000
1!
1%
#533420000000
0!
0%
#533425000000
1!
1%
#533430000000
0!
0%
#533435000000
1!
1%
#533440000000
0!
0%
#533445000000
1!
1%
#533450000000
0!
0%
#533455000000
1!
1%
#533460000000
0!
0%
#533465000000
1!
1%
#533470000000
0!
0%
#533475000000
1!
1%
#533480000000
0!
0%
#533485000000
1!
1%
#533490000000
0!
0%
#533495000000
1!
1%
#533500000000
0!
0%
#533505000000
1!
1%
#533510000000
0!
0%
#533515000000
1!
1%
#533520000000
0!
0%
#533525000000
1!
1%
#533530000000
0!
0%
#533535000000
1!
1%
#533540000000
0!
0%
#533545000000
1!
1%
#533550000000
0!
0%
#533555000000
1!
1%
#533560000000
0!
0%
#533565000000
1!
1%
#533570000000
0!
0%
#533575000000
1!
1%
#533580000000
0!
0%
#533585000000
1!
1%
#533590000000
0!
0%
#533595000000
1!
1%
#533600000000
0!
0%
#533605000000
1!
1%
#533610000000
0!
0%
#533615000000
1!
1%
#533620000000
0!
0%
#533625000000
1!
1%
#533630000000
0!
0%
#533635000000
1!
1%
#533640000000
0!
0%
#533645000000
1!
1%
#533650000000
0!
0%
#533655000000
1!
1%
#533660000000
0!
0%
#533665000000
1!
1%
#533670000000
0!
0%
#533675000000
1!
1%
#533680000000
0!
0%
#533685000000
1!
1%
#533690000000
0!
0%
#533695000000
1!
1%
#533700000000
0!
0%
#533705000000
1!
1%
#533710000000
0!
0%
#533715000000
1!
1%
#533720000000
0!
0%
#533725000000
1!
1%
#533730000000
0!
0%
#533735000000
1!
1%
#533740000000
0!
0%
#533745000000
1!
1%
#533750000000
0!
0%
#533755000000
1!
1%
#533760000000
0!
0%
#533765000000
1!
1%
#533770000000
0!
0%
#533775000000
1!
1%
#533780000000
0!
0%
#533785000000
1!
1%
#533790000000
0!
0%
#533795000000
1!
1%
#533800000000
0!
0%
#533805000000
1!
1%
#533810000000
0!
0%
#533815000000
1!
1%
#533820000000
0!
0%
#533825000000
1!
1%
#533830000000
0!
0%
#533835000000
1!
1%
#533840000000
0!
0%
#533845000000
1!
1%
#533850000000
0!
0%
#533855000000
1!
1%
#533860000000
0!
0%
#533865000000
1!
1%
#533870000000
0!
0%
#533875000000
1!
1%
#533880000000
0!
0%
#533885000000
1!
1%
#533890000000
0!
0%
#533895000000
1!
1%
#533900000000
0!
0%
#533905000000
1!
1%
#533910000000
0!
0%
#533915000000
1!
1%
#533920000000
0!
0%
#533925000000
1!
1%
#533930000000
0!
0%
#533935000000
1!
1%
#533940000000
0!
0%
#533945000000
1!
1%
#533950000000
0!
0%
#533955000000
1!
1%
#533960000000
0!
0%
#533965000000
1!
1%
#533970000000
0!
0%
#533975000000
1!
1%
#533980000000
0!
0%
#533985000000
1!
1%
#533990000000
0!
0%
#533995000000
1!
1%
#534000000000
0!
0%
#534005000000
1!
1%
#534010000000
0!
0%
#534015000000
1!
1%
#534020000000
0!
0%
#534025000000
1!
1%
#534030000000
0!
0%
#534035000000
1!
1%
#534040000000
0!
0%
#534045000000
1!
1%
#534050000000
0!
0%
#534055000000
1!
1%
#534060000000
0!
0%
#534065000000
1!
1%
#534070000000
0!
0%
#534075000000
1!
1%
#534080000000
0!
0%
#534085000000
1!
1%
#534090000000
0!
0%
#534095000000
1!
1%
#534100000000
0!
0%
#534105000000
1!
1%
#534110000000
0!
0%
#534115000000
1!
1%
#534120000000
0!
0%
#534125000000
1!
1%
#534130000000
0!
0%
#534135000000
1!
1%
#534140000000
0!
0%
#534145000000
1!
1%
#534150000000
0!
0%
#534155000000
1!
1%
#534160000000
0!
0%
#534165000000
1!
1%
#534170000000
0!
0%
#534175000000
1!
1%
#534180000000
0!
0%
#534185000000
1!
1%
#534190000000
0!
0%
#534195000000
1!
1%
#534200000000
0!
0%
#534205000000
1!
1%
#534210000000
0!
0%
#534215000000
1!
1%
#534220000000
0!
0%
#534225000000
1!
1%
#534230000000
0!
0%
#534235000000
1!
1%
#534240000000
0!
0%
#534245000000
1!
1%
#534250000000
0!
0%
#534255000000
1!
1%
#534260000000
0!
0%
#534265000000
1!
1%
#534270000000
0!
0%
#534275000000
1!
1%
#534280000000
0!
0%
#534285000000
1!
1%
#534290000000
0!
0%
#534295000000
1!
1%
#534300000000
0!
0%
#534305000000
1!
1%
#534310000000
0!
0%
#534315000000
1!
1%
#534320000000
0!
0%
#534325000000
1!
1%
#534330000000
0!
0%
#534335000000
1!
1%
#534340000000
0!
0%
#534345000000
1!
1%
#534350000000
0!
0%
#534355000000
1!
1%
#534360000000
0!
0%
#534365000000
1!
1%
#534370000000
0!
0%
#534375000000
1!
1%
#534380000000
0!
0%
#534385000000
1!
1%
#534390000000
0!
0%
#534395000000
1!
1%
#534400000000
0!
0%
#534405000000
1!
1%
#534410000000
0!
0%
#534415000000
1!
1%
#534420000000
0!
0%
#534425000000
1!
1%
#534430000000
0!
0%
#534435000000
1!
1%
#534440000000
0!
0%
#534445000000
1!
1%
#534450000000
0!
0%
#534455000000
1!
1%
#534460000000
0!
0%
#534465000000
1!
1%
#534470000000
0!
0%
#534475000000
1!
1%
#534480000000
0!
0%
#534485000000
1!
1%
#534490000000
0!
0%
#534495000000
1!
1%
#534500000000
0!
0%
#534505000000
1!
1%
#534510000000
0!
0%
#534515000000
1!
1%
#534520000000
0!
0%
#534525000000
1!
1%
#534530000000
0!
0%
#534535000000
1!
1%
#534540000000
0!
0%
#534545000000
1!
1%
#534550000000
0!
0%
#534555000000
1!
1%
#534560000000
0!
0%
#534565000000
1!
1%
#534570000000
0!
0%
#534575000000
1!
1%
#534580000000
0!
0%
#534585000000
1!
1%
#534590000000
0!
0%
#534595000000
1!
1%
#534600000000
0!
0%
#534605000000
1!
1%
#534610000000
0!
0%
#534615000000
1!
1%
#534620000000
0!
0%
#534625000000
1!
1%
#534630000000
0!
0%
#534635000000
1!
1%
#534640000000
0!
0%
#534645000000
1!
1%
#534650000000
0!
0%
#534655000000
1!
1%
#534660000000
0!
0%
#534665000000
1!
1%
#534670000000
0!
0%
#534675000000
1!
1%
#534680000000
0!
0%
#534685000000
1!
1%
#534690000000
0!
0%
#534695000000
1!
1%
#534700000000
0!
0%
#534705000000
1!
1%
#534710000000
0!
0%
#534715000000
1!
1%
#534720000000
0!
0%
#534725000000
1!
1%
#534730000000
0!
0%
#534735000000
1!
1%
#534740000000
0!
0%
#534745000000
1!
1%
#534750000000
0!
0%
#534755000000
1!
1%
#534760000000
0!
0%
#534765000000
1!
1%
#534770000000
0!
0%
#534775000000
1!
1%
#534780000000
0!
0%
#534785000000
1!
1%
#534790000000
0!
0%
#534795000000
1!
1%
#534800000000
0!
0%
#534805000000
1!
1%
#534810000000
0!
0%
#534815000000
1!
1%
#534820000000
0!
0%
#534825000000
1!
1%
#534830000000
0!
0%
#534835000000
1!
1%
#534840000000
0!
0%
#534845000000
1!
1%
#534850000000
0!
0%
#534855000000
1!
1%
#534860000000
0!
0%
#534865000000
1!
1%
#534870000000
0!
0%
#534875000000
1!
1%
#534880000000
0!
0%
#534885000000
1!
1%
#534890000000
0!
0%
#534895000000
1!
1%
#534900000000
0!
0%
#534905000000
1!
1%
#534910000000
0!
0%
#534915000000
1!
1%
#534920000000
0!
0%
#534925000000
1!
1%
#534930000000
0!
0%
#534935000000
1!
1%
#534940000000
0!
0%
#534945000000
1!
1%
#534950000000
0!
0%
#534955000000
1!
1%
#534960000000
0!
0%
#534965000000
1!
1%
#534970000000
0!
0%
#534975000000
1!
1%
#534980000000
0!
0%
#534985000000
1!
1%
#534990000000
0!
0%
#534995000000
1!
1%
#535000000000
0!
0%
#535005000000
1!
1%
#535010000000
0!
0%
#535015000000
1!
1%
#535020000000
0!
0%
#535025000000
1!
1%
#535030000000
0!
0%
#535035000000
1!
1%
#535040000000
0!
0%
#535045000000
1!
1%
#535050000000
0!
0%
#535055000000
1!
1%
#535060000000
0!
0%
#535065000000
1!
1%
#535070000000
0!
0%
#535075000000
1!
1%
#535080000000
0!
0%
#535085000000
1!
1%
#535090000000
0!
0%
#535095000000
1!
1%
#535100000000
0!
0%
#535105000000
1!
1%
#535110000000
0!
0%
#535115000000
1!
1%
#535120000000
0!
0%
#535125000000
1!
1%
#535130000000
0!
0%
#535135000000
1!
1%
#535140000000
0!
0%
#535145000000
1!
1%
#535150000000
0!
0%
#535155000000
1!
1%
#535160000000
0!
0%
#535165000000
1!
1%
#535170000000
0!
0%
#535175000000
1!
1%
#535180000000
0!
0%
#535185000000
1!
1%
#535190000000
0!
0%
#535195000000
1!
1%
#535200000000
0!
0%
#535205000000
1!
1%
#535210000000
0!
0%
#535215000000
1!
1%
#535220000000
0!
0%
#535225000000
1!
1%
#535230000000
0!
0%
#535235000000
1!
1%
#535240000000
0!
0%
#535245000000
1!
1%
#535250000000
0!
0%
#535255000000
1!
1%
#535260000000
0!
0%
#535265000000
1!
1%
#535270000000
0!
0%
#535275000000
1!
1%
#535280000000
0!
0%
#535285000000
1!
1%
#535290000000
0!
0%
#535295000000
1!
1%
#535300000000
0!
0%
#535305000000
1!
1%
#535310000000
0!
0%
#535315000000
1!
1%
#535320000000
0!
0%
#535325000000
1!
1%
#535330000000
0!
0%
#535335000000
1!
1%
#535340000000
0!
0%
#535345000000
1!
1%
#535350000000
0!
0%
#535355000000
1!
1%
#535360000000
0!
0%
#535365000000
1!
1%
#535370000000
0!
0%
#535375000000
1!
1%
#535380000000
0!
0%
#535385000000
1!
1%
#535390000000
0!
0%
#535395000000
1!
1%
#535400000000
0!
0%
#535405000000
1!
1%
#535410000000
0!
0%
#535415000000
1!
1%
#535420000000
0!
0%
#535425000000
1!
1%
#535430000000
0!
0%
#535435000000
1!
1%
#535440000000
0!
0%
#535445000000
1!
1%
#535450000000
0!
0%
#535455000000
1!
1%
#535460000000
0!
0%
#535465000000
1!
1%
#535470000000
0!
0%
#535475000000
1!
1%
#535480000000
0!
0%
#535485000000
1!
1%
#535490000000
0!
0%
#535495000000
1!
1%
#535500000000
0!
0%
#535505000000
1!
1%
#535510000000
0!
0%
#535515000000
1!
1%
#535520000000
0!
0%
#535525000000
1!
1%
#535530000000
0!
0%
#535535000000
1!
1%
#535540000000
0!
0%
#535545000000
1!
1%
#535550000000
0!
0%
#535555000000
1!
1%
#535560000000
0!
0%
#535565000000
1!
1%
#535570000000
0!
0%
#535575000000
1!
1%
#535580000000
0!
0%
#535585000000
1!
1%
#535590000000
0!
0%
#535595000000
1!
1%
#535600000000
0!
0%
#535605000000
1!
1%
#535610000000
0!
0%
#535615000000
1!
1%
#535620000000
0!
0%
#535625000000
1!
1%
#535630000000
0!
0%
#535635000000
1!
1%
#535640000000
0!
0%
#535645000000
1!
1%
#535650000000
0!
0%
#535655000000
1!
1%
#535660000000
0!
0%
#535665000000
1!
1%
#535670000000
0!
0%
#535675000000
1!
1%
#535680000000
0!
0%
#535685000000
1!
1%
#535690000000
0!
0%
#535695000000
1!
1%
#535700000000
0!
0%
#535705000000
1!
1%
#535710000000
0!
0%
#535715000000
1!
1%
#535720000000
0!
0%
#535725000000
1!
1%
#535730000000
0!
0%
#535735000000
1!
1%
#535740000000
0!
0%
#535745000000
1!
1%
#535750000000
0!
0%
#535755000000
1!
1%
#535760000000
0!
0%
#535765000000
1!
1%
#535770000000
0!
0%
#535775000000
1!
1%
#535780000000
0!
0%
#535785000000
1!
1%
#535790000000
0!
0%
#535795000000
1!
1%
#535800000000
0!
0%
#535805000000
1!
1%
#535810000000
0!
0%
#535815000000
1!
1%
#535820000000
0!
0%
#535825000000
1!
1%
#535830000000
0!
0%
#535835000000
1!
1%
#535840000000
0!
0%
#535845000000
1!
1%
#535850000000
0!
0%
#535855000000
1!
1%
#535860000000
0!
0%
#535865000000
1!
1%
#535870000000
0!
0%
#535875000000
1!
1%
#535880000000
0!
0%
#535885000000
1!
1%
#535890000000
0!
0%
#535895000000
1!
1%
#535900000000
0!
0%
#535905000000
1!
1%
#535910000000
0!
0%
#535915000000
1!
1%
#535920000000
0!
0%
#535925000000
1!
1%
#535930000000
0!
0%
#535935000000
1!
1%
#535940000000
0!
0%
#535945000000
1!
1%
#535950000000
0!
0%
#535955000000
1!
1%
#535960000000
0!
0%
#535965000000
1!
1%
#535970000000
0!
0%
#535975000000
1!
1%
#535980000000
0!
0%
#535985000000
1!
1%
#535990000000
0!
0%
#535995000000
1!
1%
#536000000000
0!
0%
#536005000000
1!
1%
#536010000000
0!
0%
#536015000000
1!
1%
#536020000000
0!
0%
#536025000000
1!
1%
#536030000000
0!
0%
#536035000000
1!
1%
#536040000000
0!
0%
#536045000000
1!
1%
#536050000000
0!
0%
#536055000000
1!
1%
#536060000000
0!
0%
#536065000000
1!
1%
#536070000000
0!
0%
#536075000000
1!
1%
#536080000000
0!
0%
#536085000000
1!
1%
#536090000000
0!
0%
#536095000000
1!
1%
#536100000000
0!
0%
#536105000000
1!
1%
#536110000000
0!
0%
#536115000000
1!
1%
#536120000000
0!
0%
#536125000000
1!
1%
#536130000000
0!
0%
#536135000000
1!
1%
#536140000000
0!
0%
#536145000000
1!
1%
#536150000000
0!
0%
#536155000000
1!
1%
#536160000000
0!
0%
#536165000000
1!
1%
#536170000000
0!
0%
#536175000000
1!
1%
#536180000000
0!
0%
#536185000000
1!
1%
#536190000000
0!
0%
#536195000000
1!
1%
#536200000000
0!
0%
#536205000000
1!
1%
#536210000000
0!
0%
#536215000000
1!
1%
#536220000000
0!
0%
#536225000000
1!
1%
#536230000000
0!
0%
#536235000000
1!
1%
#536240000000
0!
0%
#536245000000
1!
1%
#536250000000
0!
0%
#536255000000
1!
1%
#536260000000
0!
0%
#536265000000
1!
1%
#536270000000
0!
0%
#536275000000
1!
1%
#536280000000
0!
0%
#536285000000
1!
1%
#536290000000
0!
0%
#536295000000
1!
1%
#536300000000
0!
0%
#536305000000
1!
1%
#536310000000
0!
0%
#536315000000
1!
1%
#536320000000
0!
0%
#536325000000
1!
1%
#536330000000
0!
0%
#536335000000
1!
1%
#536340000000
0!
0%
#536345000000
1!
1%
#536350000000
0!
0%
#536355000000
1!
1%
#536360000000
0!
0%
#536365000000
1!
1%
#536370000000
0!
0%
#536375000000
1!
1%
#536380000000
0!
0%
#536385000000
1!
1%
#536390000000
0!
0%
#536395000000
1!
1%
#536400000000
0!
0%
#536405000000
1!
1%
#536410000000
0!
0%
#536415000000
1!
1%
#536420000000
0!
0%
#536425000000
1!
1%
#536430000000
0!
0%
#536435000000
1!
1%
#536440000000
0!
0%
#536445000000
1!
1%
#536450000000
0!
0%
#536455000000
1!
1%
#536460000000
0!
0%
#536465000000
1!
1%
#536470000000
0!
0%
#536475000000
1!
1%
#536480000000
0!
0%
#536485000000
1!
1%
#536490000000
0!
0%
#536495000000
1!
1%
#536500000000
0!
0%
#536505000000
1!
1%
#536510000000
0!
0%
#536515000000
1!
1%
#536520000000
0!
0%
#536525000000
1!
1%
#536530000000
0!
0%
#536535000000
1!
1%
#536540000000
0!
0%
#536545000000
1!
1%
#536550000000
0!
0%
#536555000000
1!
1%
#536560000000
0!
0%
#536565000000
1!
1%
#536570000000
0!
0%
#536575000000
1!
1%
#536580000000
0!
0%
#536585000000
1!
1%
#536590000000
0!
0%
#536595000000
1!
1%
#536600000000
0!
0%
#536605000000
1!
1%
#536610000000
0!
0%
#536615000000
1!
1%
#536620000000
0!
0%
#536625000000
1!
1%
#536630000000
0!
0%
#536635000000
1!
1%
#536640000000
0!
0%
#536645000000
1!
1%
#536650000000
0!
0%
#536655000000
1!
1%
#536660000000
0!
0%
#536665000000
1!
1%
#536670000000
0!
0%
#536675000000
1!
1%
#536680000000
0!
0%
#536685000000
1!
1%
#536690000000
0!
0%
#536695000000
1!
1%
#536700000000
0!
0%
#536705000000
1!
1%
#536710000000
0!
0%
#536715000000
1!
1%
#536720000000
0!
0%
#536725000000
1!
1%
#536730000000
0!
0%
#536735000000
1!
1%
#536740000000
0!
0%
#536745000000
1!
1%
#536750000000
0!
0%
#536755000000
1!
1%
#536760000000
0!
0%
#536765000000
1!
1%
#536770000000
0!
0%
#536775000000
1!
1%
#536780000000
0!
0%
#536785000000
1!
1%
#536790000000
0!
0%
#536795000000
1!
1%
#536800000000
0!
0%
#536805000000
1!
1%
#536810000000
0!
0%
#536815000000
1!
1%
#536820000000
0!
0%
#536825000000
1!
1%
#536830000000
0!
0%
#536835000000
1!
1%
#536840000000
0!
0%
#536845000000
1!
1%
#536850000000
0!
0%
#536855000000
1!
1%
#536860000000
0!
0%
#536865000000
1!
1%
#536870000000
0!
0%
#536875000000
1!
1%
#536880000000
0!
0%
#536885000000
1!
1%
#536890000000
0!
0%
#536895000000
1!
1%
#536900000000
0!
0%
#536905000000
1!
1%
#536910000000
0!
0%
#536915000000
1!
1%
#536920000000
0!
0%
#536925000000
1!
1%
#536930000000
0!
0%
#536935000000
1!
1%
#536940000000
0!
0%
#536945000000
1!
1%
#536950000000
0!
0%
#536955000000
1!
1%
#536960000000
0!
0%
#536965000000
1!
1%
#536970000000
0!
0%
#536975000000
1!
1%
#536980000000
0!
0%
#536985000000
1!
1%
#536990000000
0!
0%
#536995000000
1!
1%
#537000000000
0!
0%
#537005000000
1!
1%
#537010000000
0!
0%
#537015000000
1!
1%
#537020000000
0!
0%
#537025000000
1!
1%
#537030000000
0!
0%
#537035000000
1!
1%
#537040000000
0!
0%
#537045000000
1!
1%
#537050000000
0!
0%
#537055000000
1!
1%
#537060000000
0!
0%
#537065000000
1!
1%
#537070000000
0!
0%
#537075000000
1!
1%
#537080000000
0!
0%
#537085000000
1!
1%
#537090000000
0!
0%
#537095000000
1!
1%
#537100000000
0!
0%
#537105000000
1!
1%
#537110000000
0!
0%
#537115000000
1!
1%
#537120000000
0!
0%
#537125000000
1!
1%
#537130000000
0!
0%
#537135000000
1!
1%
#537140000000
0!
0%
#537145000000
1!
1%
#537150000000
0!
0%
#537155000000
1!
1%
#537160000000
0!
0%
#537165000000
1!
1%
#537170000000
0!
0%
#537175000000
1!
1%
#537180000000
0!
0%
#537185000000
1!
1%
#537190000000
0!
0%
#537195000000
1!
1%
#537200000000
0!
0%
#537205000000
1!
1%
#537210000000
0!
0%
#537215000000
1!
1%
#537220000000
0!
0%
#537225000000
1!
1%
#537230000000
0!
0%
#537235000000
1!
1%
#537240000000
0!
0%
#537245000000
1!
1%
#537250000000
0!
0%
#537255000000
1!
1%
#537260000000
0!
0%
#537265000000
1!
1%
#537270000000
0!
0%
#537275000000
1!
1%
#537280000000
0!
0%
#537285000000
1!
1%
#537290000000
0!
0%
#537295000000
1!
1%
#537300000000
0!
0%
#537305000000
1!
1%
#537310000000
0!
0%
#537315000000
1!
1%
#537320000000
0!
0%
#537325000000
1!
1%
#537330000000
0!
0%
#537335000000
1!
1%
#537340000000
0!
0%
#537345000000
1!
1%
#537350000000
0!
0%
#537355000000
1!
1%
#537360000000
0!
0%
#537365000000
1!
1%
#537370000000
0!
0%
#537375000000
1!
1%
#537380000000
0!
0%
#537385000000
1!
1%
#537390000000
0!
0%
#537395000000
1!
1%
#537400000000
0!
0%
#537405000000
1!
1%
#537410000000
0!
0%
#537415000000
1!
1%
#537420000000
0!
0%
#537425000000
1!
1%
#537430000000
0!
0%
#537435000000
1!
1%
#537440000000
0!
0%
#537445000000
1!
1%
#537450000000
0!
0%
#537455000000
1!
1%
#537460000000
0!
0%
#537465000000
1!
1%
#537470000000
0!
0%
#537475000000
1!
1%
#537480000000
0!
0%
#537485000000
1!
1%
#537490000000
0!
0%
#537495000000
1!
1%
#537500000000
0!
0%
#537505000000
1!
1%
#537510000000
0!
0%
#537515000000
1!
1%
#537520000000
0!
0%
#537525000000
1!
1%
#537530000000
0!
0%
#537535000000
1!
1%
#537540000000
0!
0%
#537545000000
1!
1%
#537550000000
0!
0%
#537555000000
1!
1%
#537560000000
0!
0%
#537565000000
1!
1%
#537570000000
0!
0%
#537575000000
1!
1%
#537580000000
0!
0%
#537585000000
1!
1%
#537590000000
0!
0%
#537595000000
1!
1%
#537600000000
0!
0%
#537605000000
1!
1%
#537610000000
0!
0%
#537615000000
1!
1%
#537620000000
0!
0%
#537625000000
1!
1%
#537630000000
0!
0%
#537635000000
1!
1%
#537640000000
0!
0%
#537645000000
1!
1%
#537650000000
0!
0%
#537655000000
1!
1%
#537660000000
0!
0%
#537665000000
1!
1%
#537670000000
0!
0%
#537675000000
1!
1%
#537680000000
0!
0%
#537685000000
1!
1%
#537690000000
0!
0%
#537695000000
1!
1%
#537700000000
0!
0%
#537705000000
1!
1%
#537710000000
0!
0%
#537715000000
1!
1%
#537720000000
0!
0%
#537725000000
1!
1%
#537730000000
0!
0%
#537735000000
1!
1%
#537740000000
0!
0%
#537745000000
1!
1%
#537750000000
0!
0%
#537755000000
1!
1%
#537760000000
0!
0%
#537765000000
1!
1%
#537770000000
0!
0%
#537775000000
1!
1%
#537780000000
0!
0%
#537785000000
1!
1%
#537790000000
0!
0%
#537795000000
1!
1%
#537800000000
0!
0%
#537805000000
1!
1%
#537810000000
0!
0%
#537815000000
1!
1%
#537820000000
0!
0%
#537825000000
1!
1%
#537830000000
0!
0%
#537835000000
1!
1%
#537840000000
0!
0%
#537845000000
1!
1%
#537850000000
0!
0%
#537855000000
1!
1%
#537860000000
0!
0%
#537865000000
1!
1%
#537870000000
0!
0%
#537875000000
1!
1%
#537880000000
0!
0%
#537885000000
1!
1%
#537890000000
0!
0%
#537895000000
1!
1%
#537900000000
0!
0%
#537905000000
1!
1%
#537910000000
0!
0%
#537915000000
1!
1%
#537920000000
0!
0%
#537925000000
1!
1%
#537930000000
0!
0%
#537935000000
1!
1%
#537940000000
0!
0%
#537945000000
1!
1%
#537950000000
0!
0%
#537955000000
1!
1%
#537960000000
0!
0%
#537965000000
1!
1%
#537970000000
0!
0%
#537975000000
1!
1%
#537980000000
0!
0%
#537985000000
1!
1%
#537990000000
0!
0%
#537995000000
1!
1%
#538000000000
0!
0%
#538005000000
1!
1%
#538010000000
0!
0%
#538015000000
1!
1%
#538020000000
0!
0%
#538025000000
1!
1%
#538030000000
0!
0%
#538035000000
1!
1%
#538040000000
0!
0%
#538045000000
1!
1%
#538050000000
0!
0%
#538055000000
1!
1%
#538060000000
0!
0%
#538065000000
1!
1%
#538070000000
0!
0%
#538075000000
1!
1%
#538080000000
0!
0%
#538085000000
1!
1%
#538090000000
0!
0%
#538095000000
1!
1%
#538100000000
0!
0%
#538105000000
1!
1%
#538110000000
0!
0%
#538115000000
1!
1%
#538120000000
0!
0%
#538125000000
1!
1%
#538130000000
0!
0%
#538135000000
1!
1%
#538140000000
0!
0%
#538145000000
1!
1%
#538150000000
0!
0%
#538155000000
1!
1%
#538160000000
0!
0%
#538165000000
1!
1%
#538170000000
0!
0%
#538175000000
1!
1%
#538180000000
0!
0%
#538185000000
1!
1%
#538190000000
0!
0%
#538195000000
1!
1%
#538200000000
0!
0%
#538205000000
1!
1%
#538210000000
0!
0%
#538215000000
1!
1%
#538220000000
0!
0%
#538225000000
1!
1%
#538230000000
0!
0%
#538235000000
1!
1%
#538240000000
0!
0%
#538245000000
1!
1%
#538250000000
0!
0%
#538255000000
1!
1%
#538260000000
0!
0%
#538265000000
1!
1%
#538270000000
0!
0%
#538275000000
1!
1%
#538280000000
0!
0%
#538285000000
1!
1%
#538290000000
0!
0%
#538295000000
1!
1%
#538300000000
0!
0%
#538305000000
1!
1%
#538310000000
0!
0%
#538315000000
1!
1%
#538320000000
0!
0%
#538325000000
1!
1%
#538330000000
0!
0%
#538335000000
1!
1%
#538340000000
0!
0%
#538345000000
1!
1%
#538350000000
0!
0%
#538355000000
1!
1%
#538360000000
0!
0%
#538365000000
1!
1%
#538370000000
0!
0%
#538375000000
1!
1%
#538380000000
0!
0%
#538385000000
1!
1%
#538390000000
0!
0%
#538395000000
1!
1%
#538400000000
0!
0%
#538405000000
1!
1%
#538410000000
0!
0%
#538415000000
1!
1%
#538420000000
0!
0%
#538425000000
1!
1%
#538430000000
0!
0%
#538435000000
1!
1%
#538440000000
0!
0%
#538445000000
1!
1%
#538450000000
0!
0%
#538455000000
1!
1%
#538460000000
0!
0%
#538465000000
1!
1%
#538470000000
0!
0%
#538475000000
1!
1%
#538480000000
0!
0%
#538485000000
1!
1%
#538490000000
0!
0%
#538495000000
1!
1%
#538500000000
0!
0%
#538505000000
1!
1%
#538510000000
0!
0%
#538515000000
1!
1%
#538520000000
0!
0%
#538525000000
1!
1%
#538530000000
0!
0%
#538535000000
1!
1%
#538540000000
0!
0%
#538545000000
1!
1%
#538550000000
0!
0%
#538555000000
1!
1%
#538560000000
0!
0%
#538565000000
1!
1%
#538570000000
0!
0%
#538575000000
1!
1%
#538580000000
0!
0%
#538585000000
1!
1%
#538590000000
0!
0%
#538595000000
1!
1%
#538600000000
0!
0%
#538605000000
1!
1%
#538610000000
0!
0%
#538615000000
1!
1%
#538620000000
0!
0%
#538625000000
1!
1%
#538630000000
0!
0%
#538635000000
1!
1%
#538640000000
0!
0%
#538645000000
1!
1%
#538650000000
0!
0%
#538655000000
1!
1%
#538660000000
0!
0%
#538665000000
1!
1%
#538670000000
0!
0%
#538675000000
1!
1%
#538680000000
0!
0%
#538685000000
1!
1%
#538690000000
0!
0%
#538695000000
1!
1%
#538700000000
0!
0%
#538705000000
1!
1%
#538710000000
0!
0%
#538715000000
1!
1%
#538720000000
0!
0%
#538725000000
1!
1%
#538730000000
0!
0%
#538735000000
1!
1%
#538740000000
0!
0%
#538745000000
1!
1%
#538750000000
0!
0%
#538755000000
1!
1%
#538760000000
0!
0%
#538765000000
1!
1%
#538770000000
0!
0%
#538775000000
1!
1%
#538780000000
0!
0%
#538785000000
1!
1%
#538790000000
0!
0%
#538795000000
1!
1%
#538800000000
0!
0%
#538805000000
1!
1%
#538810000000
0!
0%
#538815000000
1!
1%
#538820000000
0!
0%
#538825000000
1!
1%
#538830000000
0!
0%
#538835000000
1!
1%
#538840000000
0!
0%
#538845000000
1!
1%
#538850000000
0!
0%
#538855000000
1!
1%
#538860000000
0!
0%
#538865000000
1!
1%
#538870000000
0!
0%
#538875000000
1!
1%
#538880000000
0!
0%
#538885000000
1!
1%
#538890000000
0!
0%
#538895000000
1!
1%
#538900000000
0!
0%
#538905000000
1!
1%
#538910000000
0!
0%
#538915000000
1!
1%
#538920000000
0!
0%
#538925000000
1!
1%
#538930000000
0!
0%
#538935000000
1!
1%
#538940000000
0!
0%
#538945000000
1!
1%
#538950000000
0!
0%
#538955000000
1!
1%
#538960000000
0!
0%
#538965000000
1!
1%
#538970000000
0!
0%
#538975000000
1!
1%
#538980000000
0!
0%
#538985000000
1!
1%
#538990000000
0!
0%
#538995000000
1!
1%
#539000000000
0!
0%
#539005000000
1!
1%
#539010000000
0!
0%
#539015000000
1!
1%
#539020000000
0!
0%
#539025000000
1!
1%
#539030000000
0!
0%
#539035000000
1!
1%
#539040000000
0!
0%
#539045000000
1!
1%
#539050000000
0!
0%
#539055000000
1!
1%
#539060000000
0!
0%
#539065000000
1!
1%
#539070000000
0!
0%
#539075000000
1!
1%
#539080000000
0!
0%
#539085000000
1!
1%
#539090000000
0!
0%
#539095000000
1!
1%
#539100000000
0!
0%
#539105000000
1!
1%
#539110000000
0!
0%
#539115000000
1!
1%
#539120000000
0!
0%
#539125000000
1!
1%
#539130000000
0!
0%
#539135000000
1!
1%
#539140000000
0!
0%
#539145000000
1!
1%
#539150000000
0!
0%
#539155000000
1!
1%
#539160000000
0!
0%
#539165000000
1!
1%
#539170000000
0!
0%
#539175000000
1!
1%
#539180000000
0!
0%
#539185000000
1!
1%
#539190000000
0!
0%
#539195000000
1!
1%
#539200000000
0!
0%
#539205000000
1!
1%
#539210000000
0!
0%
#539215000000
1!
1%
#539220000000
0!
0%
#539225000000
1!
1%
#539230000000
0!
0%
#539235000000
1!
1%
#539240000000
0!
0%
#539245000000
1!
1%
#539250000000
0!
0%
#539255000000
1!
1%
#539260000000
0!
0%
#539265000000
1!
1%
#539270000000
0!
0%
#539275000000
1!
1%
#539280000000
0!
0%
#539285000000
1!
1%
#539290000000
0!
0%
#539295000000
1!
1%
#539300000000
0!
0%
#539305000000
1!
1%
#539310000000
0!
0%
#539315000000
1!
1%
#539320000000
0!
0%
#539325000000
1!
1%
#539330000000
0!
0%
#539335000000
1!
1%
#539340000000
0!
0%
#539345000000
1!
1%
#539350000000
0!
0%
#539355000000
1!
1%
#539360000000
0!
0%
#539365000000
1!
1%
#539370000000
0!
0%
#539375000000
1!
1%
#539380000000
0!
0%
#539385000000
1!
1%
#539390000000
0!
0%
#539395000000
1!
1%
#539400000000
0!
0%
#539405000000
1!
1%
#539410000000
0!
0%
#539415000000
1!
1%
#539420000000
0!
0%
#539425000000
1!
1%
#539430000000
0!
0%
#539435000000
1!
1%
#539440000000
0!
0%
#539445000000
1!
1%
#539450000000
0!
0%
#539455000000
1!
1%
#539460000000
0!
0%
#539465000000
1!
1%
#539470000000
0!
0%
#539475000000
1!
1%
#539480000000
0!
0%
#539485000000
1!
1%
#539490000000
0!
0%
#539495000000
1!
1%
#539500000000
0!
0%
#539505000000
1!
1%
#539510000000
0!
0%
#539515000000
1!
1%
#539520000000
0!
0%
#539525000000
1!
1%
#539530000000
0!
0%
#539535000000
1!
1%
#539540000000
0!
0%
#539545000000
1!
1%
#539550000000
0!
0%
#539555000000
1!
1%
#539560000000
0!
0%
#539565000000
1!
1%
#539570000000
0!
0%
#539575000000
1!
1%
#539580000000
0!
0%
#539585000000
1!
1%
#539590000000
0!
0%
#539595000000
1!
1%
#539600000000
0!
0%
#539605000000
1!
1%
#539610000000
0!
0%
#539615000000
1!
1%
#539620000000
0!
0%
#539625000000
1!
1%
#539630000000
0!
0%
#539635000000
1!
1%
#539640000000
0!
0%
#539645000000
1!
1%
#539650000000
0!
0%
#539655000000
1!
1%
#539660000000
0!
0%
#539665000000
1!
1%
#539670000000
0!
0%
#539675000000
1!
1%
#539680000000
0!
0%
#539685000000
1!
1%
#539690000000
0!
0%
#539695000000
1!
1%
#539700000000
0!
0%
#539705000000
1!
1%
#539710000000
0!
0%
#539715000000
1!
1%
#539720000000
0!
0%
#539725000000
1!
1%
#539730000000
0!
0%
#539735000000
1!
1%
#539740000000
0!
0%
#539745000000
1!
1%
#539750000000
0!
0%
#539755000000
1!
1%
#539760000000
0!
0%
#539765000000
1!
1%
#539770000000
0!
0%
#539775000000
1!
1%
#539780000000
0!
0%
#539785000000
1!
1%
#539790000000
0!
0%
#539795000000
1!
1%
#539800000000
0!
0%
#539805000000
1!
1%
#539810000000
0!
0%
#539815000000
1!
1%
#539820000000
0!
0%
#539825000000
1!
1%
#539830000000
0!
0%
#539835000000
1!
1%
#539840000000
0!
0%
#539845000000
1!
1%
#539850000000
0!
0%
#539855000000
1!
1%
#539860000000
0!
0%
#539865000000
1!
1%
#539870000000
0!
0%
#539875000000
1!
1%
#539880000000
0!
0%
#539885000000
1!
1%
#539890000000
0!
0%
#539895000000
1!
1%
#539900000000
0!
0%
#539905000000
1!
1%
#539910000000
0!
0%
#539915000000
1!
1%
#539920000000
0!
0%
#539925000000
1!
1%
#539930000000
0!
0%
#539935000000
1!
1%
#539940000000
0!
0%
#539945000000
1!
1%
#539950000000
0!
0%
#539955000000
1!
1%
#539960000000
0!
0%
#539965000000
1!
1%
#539970000000
0!
0%
#539975000000
1!
1%
#539980000000
0!
0%
#539985000000
1!
1%
#539990000000
0!
0%
#539995000000
1!
1%
#540000000000
0!
0%
#540005000000
1!
1%
#540010000000
0!
0%
#540015000000
1!
1%
#540020000000
0!
0%
#540025000000
1!
1%
#540030000000
0!
0%
#540035000000
1!
1%
#540040000000
0!
0%
#540045000000
1!
1%
#540050000000
0!
0%
#540055000000
1!
1%
#540060000000
0!
0%
#540065000000
1!
1%
#540070000000
0!
0%
#540075000000
1!
1%
#540080000000
0!
0%
#540085000000
1!
1%
#540090000000
0!
0%
#540095000000
1!
1%
#540100000000
0!
0%
#540105000000
1!
1%
#540110000000
0!
0%
#540115000000
1!
1%
#540120000000
0!
0%
#540125000000
1!
1%
#540130000000
0!
0%
#540135000000
1!
1%
#540140000000
0!
0%
#540145000000
1!
1%
#540150000000
0!
0%
#540155000000
1!
1%
#540160000000
0!
0%
#540165000000
1!
1%
#540170000000
0!
0%
#540175000000
1!
1%
#540180000000
0!
0%
#540185000000
1!
1%
#540190000000
0!
0%
#540195000000
1!
1%
#540200000000
0!
0%
#540205000000
1!
1%
#540210000000
0!
0%
#540215000000
1!
1%
#540220000000
0!
0%
#540225000000
1!
1%
#540230000000
0!
0%
#540235000000
1!
1%
#540240000000
0!
0%
#540245000000
1!
1%
#540250000000
0!
0%
#540255000000
1!
1%
#540260000000
0!
0%
#540265000000
1!
1%
#540270000000
0!
0%
#540275000000
1!
1%
#540280000000
0!
0%
#540285000000
1!
1%
#540290000000
0!
0%
#540295000000
1!
1%
#540300000000
0!
0%
#540305000000
1!
1%
#540310000000
0!
0%
#540315000000
1!
1%
#540320000000
0!
0%
#540325000000
1!
1%
#540330000000
0!
0%
#540335000000
1!
1%
#540340000000
0!
0%
#540345000000
1!
1%
#540350000000
0!
0%
#540355000000
1!
1%
#540360000000
0!
0%
#540365000000
1!
1%
#540370000000
0!
0%
#540375000000
1!
1%
#540380000000
0!
0%
#540385000000
1!
1%
#540390000000
0!
0%
#540395000000
1!
1%
#540400000000
0!
0%
#540405000000
1!
1%
#540410000000
0!
0%
#540415000000
1!
1%
#540420000000
0!
0%
#540425000000
1!
1%
#540430000000
0!
0%
#540435000000
1!
1%
#540440000000
0!
0%
#540445000000
1!
1%
#540450000000
0!
0%
#540455000000
1!
1%
#540460000000
0!
0%
#540465000000
1!
1%
#540470000000
0!
0%
#540475000000
1!
1%
#540480000000
0!
0%
#540485000000
1!
1%
#540490000000
0!
0%
#540495000000
1!
1%
#540500000000
0!
0%
#540505000000
1!
1%
#540510000000
0!
0%
#540515000000
1!
1%
#540520000000
0!
0%
#540525000000
1!
1%
#540530000000
0!
0%
#540535000000
1!
1%
#540540000000
0!
0%
#540545000000
1!
1%
#540550000000
0!
0%
#540555000000
1!
1%
#540560000000
0!
0%
#540565000000
1!
1%
#540570000000
0!
0%
#540575000000
1!
1%
#540580000000
0!
0%
#540585000000
1!
1%
#540590000000
0!
0%
#540595000000
1!
1%
#540600000000
0!
0%
#540605000000
1!
1%
#540610000000
0!
0%
#540615000000
1!
1%
#540620000000
0!
0%
#540625000000
1!
1%
#540630000000
0!
0%
#540635000000
1!
1%
#540640000000
0!
0%
#540645000000
1!
1%
#540650000000
0!
0%
#540655000000
1!
1%
#540660000000
0!
0%
#540665000000
1!
1%
#540670000000
0!
0%
#540675000000
1!
1%
#540680000000
0!
0%
#540685000000
1!
1%
#540690000000
0!
0%
#540695000000
1!
1%
#540700000000
0!
0%
#540705000000
1!
1%
#540710000000
0!
0%
#540715000000
1!
1%
#540720000000
0!
0%
#540725000000
1!
1%
#540730000000
0!
0%
#540735000000
1!
1%
#540740000000
0!
0%
#540745000000
1!
1%
#540750000000
0!
0%
#540755000000
1!
1%
#540760000000
0!
0%
#540765000000
1!
1%
#540770000000
0!
0%
#540775000000
1!
1%
#540780000000
0!
0%
#540785000000
1!
1%
#540790000000
0!
0%
#540795000000
1!
1%
#540800000000
0!
0%
#540805000000
1!
1%
#540810000000
0!
0%
#540815000000
1!
1%
#540820000000
0!
0%
#540825000000
1!
1%
#540830000000
0!
0%
#540835000000
1!
1%
#540840000000
0!
0%
#540845000000
1!
1%
#540850000000
0!
0%
#540855000000
1!
1%
#540860000000
0!
0%
#540865000000
1!
1%
#540870000000
0!
0%
#540875000000
1!
1%
#540880000000
0!
0%
#540885000000
1!
1%
#540890000000
0!
0%
#540895000000
1!
1%
#540900000000
0!
0%
#540905000000
1!
1%
#540910000000
0!
0%
#540915000000
1!
1%
#540920000000
0!
0%
#540925000000
1!
1%
#540930000000
0!
0%
#540935000000
1!
1%
#540940000000
0!
0%
#540945000000
1!
1%
#540950000000
0!
0%
#540955000000
1!
1%
#540960000000
0!
0%
#540965000000
1!
1%
#540970000000
0!
0%
#540975000000
1!
1%
#540980000000
0!
0%
#540985000000
1!
1%
#540990000000
0!
0%
#540995000000
1!
1%
#541000000000
0!
0%
#541005000000
1!
1%
#541010000000
0!
0%
#541015000000
1!
1%
#541020000000
0!
0%
#541025000000
1!
1%
#541030000000
0!
0%
#541035000000
1!
1%
#541040000000
0!
0%
#541045000000
1!
1%
#541050000000
0!
0%
#541055000000
1!
1%
#541060000000
0!
0%
#541065000000
1!
1%
#541070000000
0!
0%
#541075000000
1!
1%
#541080000000
0!
0%
#541085000000
1!
1%
#541090000000
0!
0%
#541095000000
1!
1%
#541100000000
0!
0%
#541105000000
1!
1%
#541110000000
0!
0%
#541115000000
1!
1%
#541120000000
0!
0%
#541125000000
1!
1%
#541130000000
0!
0%
#541135000000
1!
1%
#541140000000
0!
0%
#541145000000
1!
1%
#541150000000
0!
0%
#541155000000
1!
1%
#541160000000
0!
0%
#541165000000
1!
1%
#541170000000
0!
0%
#541175000000
1!
1%
#541180000000
0!
0%
#541185000000
1!
1%
#541190000000
0!
0%
#541195000000
1!
1%
#541200000000
0!
0%
#541205000000
1!
1%
#541210000000
0!
0%
#541215000000
1!
1%
#541220000000
0!
0%
#541225000000
1!
1%
#541230000000
0!
0%
#541235000000
1!
1%
#541240000000
0!
0%
#541245000000
1!
1%
#541250000000
0!
0%
#541255000000
1!
1%
#541260000000
0!
0%
#541265000000
1!
1%
#541270000000
0!
0%
#541275000000
1!
1%
#541280000000
0!
0%
#541285000000
1!
1%
#541290000000
0!
0%
#541295000000
1!
1%
#541300000000
0!
0%
#541305000000
1!
1%
#541310000000
0!
0%
#541315000000
1!
1%
#541320000000
0!
0%
#541325000000
1!
1%
#541330000000
0!
0%
#541335000000
1!
1%
#541340000000
0!
0%
#541345000000
1!
1%
#541350000000
0!
0%
#541355000000
1!
1%
#541360000000
0!
0%
#541365000000
1!
1%
#541370000000
0!
0%
#541375000000
1!
1%
#541380000000
0!
0%
#541385000000
1!
1%
#541390000000
0!
0%
#541395000000
1!
1%
#541400000000
0!
0%
#541405000000
1!
1%
#541410000000
0!
0%
#541415000000
1!
1%
#541420000000
0!
0%
#541425000000
1!
1%
#541430000000
0!
0%
#541435000000
1!
1%
#541440000000
0!
0%
#541445000000
1!
1%
#541450000000
0!
0%
#541455000000
1!
1%
#541460000000
0!
0%
#541465000000
1!
1%
#541470000000
0!
0%
#541475000000
1!
1%
#541480000000
0!
0%
#541485000000
1!
1%
#541490000000
0!
0%
#541495000000
1!
1%
#541500000000
0!
0%
#541505000000
1!
1%
#541510000000
0!
0%
#541515000000
1!
1%
#541520000000
0!
0%
#541525000000
1!
1%
#541530000000
0!
0%
#541535000000
1!
1%
#541540000000
0!
0%
#541545000000
1!
1%
#541550000000
0!
0%
#541555000000
1!
1%
#541560000000
0!
0%
#541565000000
1!
1%
#541570000000
0!
0%
#541575000000
1!
1%
#541580000000
0!
0%
#541585000000
1!
1%
#541590000000
0!
0%
#541595000000
1!
1%
#541600000000
0!
0%
#541605000000
1!
1%
#541610000000
0!
0%
#541615000000
1!
1%
#541620000000
0!
0%
#541625000000
1!
1%
#541630000000
0!
0%
#541635000000
1!
1%
#541640000000
0!
0%
#541645000000
1!
1%
#541650000000
0!
0%
#541655000000
1!
1%
#541660000000
0!
0%
#541665000000
1!
1%
#541670000000
0!
0%
#541675000000
1!
1%
#541680000000
0!
0%
#541685000000
1!
1%
#541690000000
0!
0%
#541695000000
1!
1%
#541700000000
0!
0%
#541705000000
1!
1%
#541710000000
0!
0%
#541715000000
1!
1%
#541720000000
0!
0%
#541725000000
1!
1%
#541730000000
0!
0%
#541735000000
1!
1%
#541740000000
0!
0%
#541745000000
1!
1%
#541750000000
0!
0%
#541755000000
1!
1%
#541760000000
0!
0%
#541765000000
1!
1%
#541770000000
0!
0%
#541775000000
1!
1%
#541780000000
0!
0%
#541785000000
1!
1%
#541790000000
0!
0%
#541795000000
1!
1%
#541800000000
0!
0%
#541805000000
1!
1%
#541810000000
0!
0%
#541815000000
1!
1%
#541820000000
0!
0%
#541825000000
1!
1%
#541830000000
0!
0%
#541835000000
1!
1%
#541840000000
0!
0%
#541845000000
1!
1%
#541850000000
0!
0%
#541855000000
1!
1%
#541860000000
0!
0%
#541865000000
1!
1%
#541870000000
0!
0%
#541875000000
1!
1%
#541880000000
0!
0%
#541885000000
1!
1%
#541890000000
0!
0%
#541895000000
1!
1%
#541900000000
0!
0%
#541905000000
1!
1%
#541910000000
0!
0%
#541915000000
1!
1%
#541920000000
0!
0%
#541925000000
1!
1%
#541930000000
0!
0%
#541935000000
1!
1%
#541940000000
0!
0%
#541945000000
1!
1%
#541950000000
0!
0%
#541955000000
1!
1%
#541960000000
0!
0%
#541965000000
1!
1%
#541970000000
0!
0%
#541975000000
1!
1%
#541980000000
0!
0%
#541985000000
1!
1%
#541990000000
0!
0%
#541995000000
1!
1%
#542000000000
0!
0%
#542005000000
1!
1%
#542010000000
0!
0%
#542015000000
1!
1%
#542020000000
0!
0%
#542025000000
1!
1%
#542030000000
0!
0%
#542035000000
1!
1%
#542040000000
0!
0%
#542045000000
1!
1%
#542050000000
0!
0%
#542055000000
1!
1%
#542060000000
0!
0%
#542065000000
1!
1%
#542070000000
0!
0%
#542075000000
1!
1%
#542080000000
0!
0%
#542085000000
1!
1%
#542090000000
0!
0%
#542095000000
1!
1%
#542100000000
0!
0%
#542105000000
1!
1%
#542110000000
0!
0%
#542115000000
1!
1%
#542120000000
0!
0%
#542125000000
1!
1%
#542130000000
0!
0%
#542135000000
1!
1%
#542140000000
0!
0%
#542145000000
1!
1%
#542150000000
0!
0%
#542155000000
1!
1%
#542160000000
0!
0%
#542165000000
1!
1%
#542170000000
0!
0%
#542175000000
1!
1%
#542180000000
0!
0%
#542185000000
1!
1%
#542190000000
0!
0%
#542195000000
1!
1%
#542200000000
0!
0%
#542205000000
1!
1%
#542210000000
0!
0%
#542215000000
1!
1%
#542220000000
0!
0%
#542225000000
1!
1%
#542230000000
0!
0%
#542235000000
1!
1%
#542240000000
0!
0%
#542245000000
1!
1%
#542250000000
0!
0%
#542255000000
1!
1%
#542260000000
0!
0%
#542265000000
1!
1%
#542270000000
0!
0%
#542275000000
1!
1%
#542280000000
0!
0%
#542285000000
1!
1%
#542290000000
0!
0%
#542295000000
1!
1%
#542300000000
0!
0%
#542305000000
1!
1%
#542310000000
0!
0%
#542315000000
1!
1%
#542320000000
0!
0%
#542325000000
1!
1%
#542330000000
0!
0%
#542335000000
1!
1%
#542340000000
0!
0%
#542345000000
1!
1%
#542350000000
0!
0%
#542355000000
1!
1%
#542360000000
0!
0%
#542365000000
1!
1%
#542370000000
0!
0%
#542375000000
1!
1%
#542380000000
0!
0%
#542385000000
1!
1%
#542390000000
0!
0%
#542395000000
1!
1%
#542400000000
0!
0%
#542405000000
1!
1%
#542410000000
0!
0%
#542415000000
1!
1%
#542420000000
0!
0%
#542425000000
1!
1%
#542430000000
0!
0%
#542435000000
1!
1%
#542440000000
0!
0%
#542445000000
1!
1%
#542450000000
0!
0%
#542455000000
1!
1%
#542460000000
0!
0%
#542465000000
1!
1%
#542470000000
0!
0%
#542475000000
1!
1%
#542480000000
0!
0%
#542485000000
1!
1%
#542490000000
0!
0%
#542495000000
1!
1%
#542500000000
0!
0%
#542505000000
1!
1%
#542510000000
0!
0%
#542515000000
1!
1%
#542520000000
0!
0%
#542525000000
1!
1%
#542530000000
0!
0%
#542535000000
1!
1%
#542540000000
0!
0%
#542545000000
1!
1%
#542550000000
0!
0%
#542555000000
1!
1%
#542560000000
0!
0%
#542565000000
1!
1%
#542570000000
0!
0%
#542575000000
1!
1%
#542580000000
0!
0%
#542585000000
1!
1%
#542590000000
0!
0%
#542595000000
1!
1%
#542600000000
0!
0%
#542605000000
1!
1%
#542610000000
0!
0%
#542615000000
1!
1%
#542620000000
0!
0%
#542625000000
1!
1%
#542630000000
0!
0%
#542635000000
1!
1%
#542640000000
0!
0%
#542645000000
1!
1%
#542650000000
0!
0%
#542655000000
1!
1%
#542660000000
0!
0%
#542665000000
1!
1%
#542670000000
0!
0%
#542675000000
1!
1%
#542680000000
0!
0%
#542685000000
1!
1%
#542690000000
0!
0%
#542695000000
1!
1%
#542700000000
0!
0%
#542705000000
1!
1%
#542710000000
0!
0%
#542715000000
1!
1%
#542720000000
0!
0%
#542725000000
1!
1%
#542730000000
0!
0%
#542735000000
1!
1%
#542740000000
0!
0%
#542745000000
1!
1%
#542750000000
0!
0%
#542755000000
1!
1%
#542760000000
0!
0%
#542765000000
1!
1%
#542770000000
0!
0%
#542775000000
1!
1%
#542780000000
0!
0%
#542785000000
1!
1%
#542790000000
0!
0%
#542795000000
1!
1%
#542800000000
0!
0%
#542805000000
1!
1%
#542810000000
0!
0%
#542815000000
1!
1%
#542820000000
0!
0%
#542825000000
1!
1%
#542830000000
0!
0%
#542835000000
1!
1%
#542840000000
0!
0%
#542845000000
1!
1%
#542850000000
0!
0%
#542855000000
1!
1%
#542860000000
0!
0%
#542865000000
1!
1%
#542870000000
0!
0%
#542875000000
1!
1%
#542880000000
0!
0%
#542885000000
1!
1%
#542890000000
0!
0%
#542895000000
1!
1%
#542900000000
0!
0%
#542905000000
1!
1%
#542910000000
0!
0%
#542915000000
1!
1%
#542920000000
0!
0%
#542925000000
1!
1%
#542930000000
0!
0%
#542935000000
1!
1%
#542940000000
0!
0%
#542945000000
1!
1%
#542950000000
0!
0%
#542955000000
1!
1%
#542960000000
0!
0%
#542965000000
1!
1%
#542970000000
0!
0%
#542975000000
1!
1%
#542980000000
0!
0%
#542985000000
1!
1%
#542990000000
0!
0%
#542995000000
1!
1%
#543000000000
0!
0%
#543005000000
1!
1%
#543010000000
0!
0%
#543015000000
1!
1%
#543020000000
0!
0%
#543025000000
1!
1%
#543030000000
0!
0%
#543035000000
1!
1%
#543040000000
0!
0%
#543045000000
1!
1%
#543050000000
0!
0%
#543055000000
1!
1%
#543060000000
0!
0%
#543065000000
1!
1%
#543070000000
0!
0%
#543075000000
1!
1%
#543080000000
0!
0%
#543085000000
1!
1%
#543090000000
0!
0%
#543095000000
1!
1%
#543100000000
0!
0%
#543105000000
1!
1%
#543110000000
0!
0%
#543115000000
1!
1%
#543120000000
0!
0%
#543125000000
1!
1%
#543130000000
0!
0%
#543135000000
1!
1%
#543140000000
0!
0%
#543145000000
1!
1%
#543150000000
0!
0%
#543155000000
1!
1%
#543160000000
0!
0%
#543165000000
1!
1%
#543170000000
0!
0%
#543175000000
1!
1%
#543180000000
0!
0%
#543185000000
1!
1%
#543190000000
0!
0%
#543195000000
1!
1%
#543200000000
0!
0%
#543205000000
1!
1%
#543210000000
0!
0%
#543215000000
1!
1%
#543220000000
0!
0%
#543225000000
1!
1%
#543230000000
0!
0%
#543235000000
1!
1%
#543240000000
0!
0%
#543245000000
1!
1%
#543250000000
0!
0%
#543255000000
1!
1%
#543260000000
0!
0%
#543265000000
1!
1%
#543270000000
0!
0%
#543275000000
1!
1%
#543280000000
0!
0%
#543285000000
1!
1%
#543290000000
0!
0%
#543295000000
1!
1%
#543300000000
0!
0%
#543305000000
1!
1%
#543310000000
0!
0%
#543315000000
1!
1%
#543320000000
0!
0%
#543325000000
1!
1%
#543330000000
0!
0%
#543335000000
1!
1%
#543340000000
0!
0%
#543345000000
1!
1%
#543350000000
0!
0%
#543355000000
1!
1%
#543360000000
0!
0%
#543365000000
1!
1%
#543370000000
0!
0%
#543375000000
1!
1%
#543380000000
0!
0%
#543385000000
1!
1%
#543390000000
0!
0%
#543395000000
1!
1%
#543400000000
0!
0%
#543405000000
1!
1%
#543410000000
0!
0%
#543415000000
1!
1%
#543420000000
0!
0%
#543425000000
1!
1%
#543430000000
0!
0%
#543435000000
1!
1%
#543440000000
0!
0%
#543445000000
1!
1%
#543450000000
0!
0%
#543455000000
1!
1%
#543460000000
0!
0%
#543465000000
1!
1%
#543470000000
0!
0%
#543475000000
1!
1%
#543480000000
0!
0%
#543485000000
1!
1%
#543490000000
0!
0%
#543495000000
1!
1%
#543500000000
0!
0%
#543505000000
1!
1%
#543510000000
0!
0%
#543515000000
1!
1%
#543520000000
0!
0%
#543525000000
1!
1%
#543530000000
0!
0%
#543535000000
1!
1%
#543540000000
0!
0%
#543545000000
1!
1%
#543550000000
0!
0%
#543555000000
1!
1%
#543560000000
0!
0%
#543565000000
1!
1%
#543570000000
0!
0%
#543575000000
1!
1%
#543580000000
0!
0%
#543585000000
1!
1%
#543590000000
0!
0%
#543595000000
1!
1%
#543600000000
0!
0%
#543605000000
1!
1%
#543610000000
0!
0%
#543615000000
1!
1%
#543620000000
0!
0%
#543625000000
1!
1%
#543630000000
0!
0%
#543635000000
1!
1%
#543640000000
0!
0%
#543645000000
1!
1%
#543650000000
0!
0%
#543655000000
1!
1%
#543660000000
0!
0%
#543665000000
1!
1%
#543670000000
0!
0%
#543675000000
1!
1%
#543680000000
0!
0%
#543685000000
1!
1%
#543690000000
0!
0%
#543695000000
1!
1%
#543700000000
0!
0%
#543705000000
1!
1%
#543710000000
0!
0%
#543715000000
1!
1%
#543720000000
0!
0%
#543725000000
1!
1%
#543730000000
0!
0%
#543735000000
1!
1%
#543740000000
0!
0%
#543745000000
1!
1%
#543750000000
0!
0%
#543755000000
1!
1%
#543760000000
0!
0%
#543765000000
1!
1%
#543770000000
0!
0%
#543775000000
1!
1%
#543780000000
0!
0%
#543785000000
1!
1%
#543790000000
0!
0%
#543795000000
1!
1%
#543800000000
0!
0%
#543805000000
1!
1%
#543810000000
0!
0%
#543815000000
1!
1%
#543820000000
0!
0%
#543825000000
1!
1%
#543830000000
0!
0%
#543835000000
1!
1%
#543840000000
0!
0%
#543845000000
1!
1%
#543850000000
0!
0%
#543855000000
1!
1%
#543860000000
0!
0%
#543865000000
1!
1%
#543870000000
0!
0%
#543875000000
1!
1%
#543880000000
0!
0%
#543885000000
1!
1%
#543890000000
0!
0%
#543895000000
1!
1%
#543900000000
0!
0%
#543905000000
1!
1%
#543910000000
0!
0%
#543915000000
1!
1%
#543920000000
0!
0%
#543925000000
1!
1%
#543930000000
0!
0%
#543935000000
1!
1%
#543940000000
0!
0%
#543945000000
1!
1%
#543950000000
0!
0%
#543955000000
1!
1%
#543960000000
0!
0%
#543965000000
1!
1%
#543970000000
0!
0%
#543975000000
1!
1%
#543980000000
0!
0%
#543985000000
1!
1%
#543990000000
0!
0%
#543995000000
1!
1%
#544000000000
0!
0%
#544005000000
1!
1%
#544010000000
0!
0%
#544015000000
1!
1%
#544020000000
0!
0%
#544025000000
1!
1%
#544030000000
0!
0%
#544035000000
1!
1%
#544040000000
0!
0%
#544045000000
1!
1%
#544050000000
0!
0%
#544055000000
1!
1%
#544060000000
0!
0%
#544065000000
1!
1%
#544070000000
0!
0%
#544075000000
1!
1%
#544080000000
0!
0%
#544085000000
1!
1%
#544090000000
0!
0%
#544095000000
1!
1%
#544100000000
0!
0%
#544105000000
1!
1%
#544110000000
0!
0%
#544115000000
1!
1%
#544120000000
0!
0%
#544125000000
1!
1%
#544130000000
0!
0%
#544135000000
1!
1%
#544140000000
0!
0%
#544145000000
1!
1%
#544150000000
0!
0%
#544155000000
1!
1%
#544160000000
0!
0%
#544165000000
1!
1%
#544170000000
0!
0%
#544175000000
1!
1%
#544180000000
0!
0%
#544185000000
1!
1%
#544190000000
0!
0%
#544195000000
1!
1%
#544200000000
0!
0%
#544205000000
1!
1%
#544210000000
0!
0%
#544215000000
1!
1%
#544220000000
0!
0%
#544225000000
1!
1%
#544230000000
0!
0%
#544235000000
1!
1%
#544240000000
0!
0%
#544245000000
1!
1%
#544250000000
0!
0%
#544255000000
1!
1%
#544260000000
0!
0%
#544265000000
1!
1%
#544270000000
0!
0%
#544275000000
1!
1%
#544280000000
0!
0%
#544285000000
1!
1%
#544290000000
0!
0%
#544295000000
1!
1%
#544300000000
0!
0%
#544305000000
1!
1%
#544310000000
0!
0%
#544315000000
1!
1%
#544320000000
0!
0%
#544325000000
1!
1%
#544330000000
0!
0%
#544335000000
1!
1%
#544340000000
0!
0%
#544345000000
1!
1%
#544350000000
0!
0%
#544355000000
1!
1%
#544360000000
0!
0%
#544365000000
1!
1%
#544370000000
0!
0%
#544375000000
1!
1%
#544380000000
0!
0%
#544385000000
1!
1%
#544390000000
0!
0%
#544395000000
1!
1%
#544400000000
0!
0%
#544405000000
1!
1%
#544410000000
0!
0%
#544415000000
1!
1%
#544420000000
0!
0%
#544425000000
1!
1%
#544430000000
0!
0%
#544435000000
1!
1%
#544440000000
0!
0%
#544445000000
1!
1%
#544450000000
0!
0%
#544455000000
1!
1%
#544460000000
0!
0%
#544465000000
1!
1%
#544470000000
0!
0%
#544475000000
1!
1%
#544480000000
0!
0%
#544485000000
1!
1%
#544490000000
0!
0%
#544495000000
1!
1%
#544500000000
0!
0%
#544505000000
1!
1%
#544510000000
0!
0%
#544515000000
1!
1%
#544520000000
0!
0%
#544525000000
1!
1%
#544530000000
0!
0%
#544535000000
1!
1%
#544540000000
0!
0%
#544545000000
1!
1%
#544550000000
0!
0%
#544555000000
1!
1%
#544560000000
0!
0%
#544565000000
1!
1%
#544570000000
0!
0%
#544575000000
1!
1%
#544580000000
0!
0%
#544585000000
1!
1%
#544590000000
0!
0%
#544595000000
1!
1%
#544600000000
0!
0%
#544605000000
1!
1%
#544610000000
0!
0%
#544615000000
1!
1%
#544620000000
0!
0%
#544625000000
1!
1%
#544630000000
0!
0%
#544635000000
1!
1%
#544640000000
0!
0%
#544645000000
1!
1%
#544650000000
0!
0%
#544655000000
1!
1%
#544660000000
0!
0%
#544665000000
1!
1%
#544670000000
0!
0%
#544675000000
1!
1%
#544680000000
0!
0%
#544685000000
1!
1%
#544690000000
0!
0%
#544695000000
1!
1%
#544700000000
0!
0%
#544705000000
1!
1%
#544710000000
0!
0%
#544715000000
1!
1%
#544720000000
0!
0%
#544725000000
1!
1%
#544730000000
0!
0%
#544735000000
1!
1%
#544740000000
0!
0%
#544745000000
1!
1%
#544750000000
0!
0%
#544755000000
1!
1%
#544760000000
0!
0%
#544765000000
1!
1%
#544770000000
0!
0%
#544775000000
1!
1%
#544780000000
0!
0%
#544785000000
1!
1%
#544790000000
0!
0%
#544795000000
1!
1%
#544800000000
0!
0%
#544805000000
1!
1%
#544810000000
0!
0%
#544815000000
1!
1%
#544820000000
0!
0%
#544825000000
1!
1%
#544830000000
0!
0%
#544835000000
1!
1%
#544840000000
0!
0%
#544845000000
1!
1%
#544850000000
0!
0%
#544855000000
1!
1%
#544860000000
0!
0%
#544865000000
1!
1%
#544870000000
0!
0%
#544875000000
1!
1%
#544880000000
0!
0%
#544885000000
1!
1%
#544890000000
0!
0%
#544895000000
1!
1%
#544900000000
0!
0%
#544905000000
1!
1%
#544910000000
0!
0%
#544915000000
1!
1%
#544920000000
0!
0%
#544925000000
1!
1%
#544930000000
0!
0%
#544935000000
1!
1%
#544940000000
0!
0%
#544945000000
1!
1%
#544950000000
0!
0%
#544955000000
1!
1%
#544960000000
0!
0%
#544965000000
1!
1%
#544970000000
0!
0%
#544975000000
1!
1%
#544980000000
0!
0%
#544985000000
1!
1%
#544990000000
0!
0%
#544995000000
1!
1%
#545000000000
0!
0%
#545005000000
1!
1%
#545010000000
0!
0%
#545015000000
1!
1%
#545020000000
0!
0%
#545025000000
1!
1%
#545030000000
0!
0%
#545035000000
1!
1%
#545040000000
0!
0%
#545045000000
1!
1%
#545050000000
0!
0%
#545055000000
1!
1%
#545060000000
0!
0%
#545065000000
1!
1%
#545070000000
0!
0%
#545075000000
1!
1%
#545080000000
0!
0%
#545085000000
1!
1%
#545090000000
0!
0%
#545095000000
1!
1%
#545100000000
0!
0%
#545105000000
1!
1%
#545110000000
0!
0%
#545115000000
1!
1%
#545120000000
0!
0%
#545125000000
1!
1%
#545130000000
0!
0%
#545135000000
1!
1%
#545140000000
0!
0%
#545145000000
1!
1%
#545150000000
0!
0%
#545155000000
1!
1%
#545160000000
0!
0%
#545165000000
1!
1%
#545170000000
0!
0%
#545175000000
1!
1%
#545180000000
0!
0%
#545185000000
1!
1%
#545190000000
0!
0%
#545195000000
1!
1%
#545200000000
0!
0%
#545205000000
1!
1%
#545210000000
0!
0%
#545215000000
1!
1%
#545220000000
0!
0%
#545225000000
1!
1%
#545230000000
0!
0%
#545235000000
1!
1%
#545240000000
0!
0%
#545245000000
1!
1%
#545250000000
0!
0%
#545255000000
1!
1%
#545260000000
0!
0%
#545265000000
1!
1%
#545270000000
0!
0%
#545275000000
1!
1%
#545280000000
0!
0%
#545285000000
1!
1%
#545290000000
0!
0%
#545295000000
1!
1%
#545300000000
0!
0%
#545305000000
1!
1%
#545310000000
0!
0%
#545315000000
1!
1%
#545320000000
0!
0%
#545325000000
1!
1%
#545330000000
0!
0%
#545335000000
1!
1%
#545340000000
0!
0%
#545345000000
1!
1%
#545350000000
0!
0%
#545355000000
1!
1%
#545360000000
0!
0%
#545365000000
1!
1%
#545370000000
0!
0%
#545375000000
1!
1%
#545380000000
0!
0%
#545385000000
1!
1%
#545390000000
0!
0%
#545395000000
1!
1%
#545400000000
0!
0%
#545405000000
1!
1%
#545410000000
0!
0%
#545415000000
1!
1%
#545420000000
0!
0%
#545425000000
1!
1%
#545430000000
0!
0%
#545435000000
1!
1%
#545440000000
0!
0%
#545445000000
1!
1%
#545450000000
0!
0%
#545455000000
1!
1%
#545460000000
0!
0%
#545465000000
1!
1%
#545470000000
0!
0%
#545475000000
1!
1%
#545480000000
0!
0%
#545485000000
1!
1%
#545490000000
0!
0%
#545495000000
1!
1%
#545500000000
0!
0%
#545505000000
1!
1%
#545510000000
0!
0%
#545515000000
1!
1%
#545520000000
0!
0%
#545525000000
1!
1%
#545530000000
0!
0%
#545535000000
1!
1%
#545540000000
0!
0%
#545545000000
1!
1%
#545550000000
0!
0%
#545555000000
1!
1%
#545560000000
0!
0%
#545565000000
1!
1%
#545570000000
0!
0%
#545575000000
1!
1%
#545580000000
0!
0%
#545585000000
1!
1%
#545590000000
0!
0%
#545595000000
1!
1%
#545600000000
0!
0%
#545605000000
1!
1%
#545610000000
0!
0%
#545615000000
1!
1%
#545620000000
0!
0%
#545625000000
1!
1%
#545630000000
0!
0%
#545635000000
1!
1%
#545640000000
0!
0%
#545645000000
1!
1%
#545650000000
0!
0%
#545655000000
1!
1%
#545660000000
0!
0%
#545665000000
1!
1%
#545670000000
0!
0%
#545675000000
1!
1%
#545680000000
0!
0%
#545685000000
1!
1%
#545690000000
0!
0%
#545695000000
1!
1%
#545700000000
0!
0%
#545705000000
1!
1%
#545710000000
0!
0%
#545715000000
1!
1%
#545720000000
0!
0%
#545725000000
1!
1%
#545730000000
0!
0%
#545735000000
1!
1%
#545740000000
0!
0%
#545745000000
1!
1%
#545750000000
0!
0%
#545755000000
1!
1%
#545760000000
0!
0%
#545765000000
1!
1%
#545770000000
0!
0%
#545775000000
1!
1%
#545780000000
0!
0%
#545785000000
1!
1%
#545790000000
0!
0%
#545795000000
1!
1%
#545800000000
0!
0%
#545805000000
1!
1%
#545810000000
0!
0%
#545815000000
1!
1%
#545820000000
0!
0%
#545825000000
1!
1%
#545830000000
0!
0%
#545835000000
1!
1%
#545840000000
0!
0%
#545845000000
1!
1%
#545850000000
0!
0%
#545855000000
1!
1%
#545860000000
0!
0%
#545865000000
1!
1%
#545870000000
0!
0%
#545875000000
1!
1%
#545880000000
0!
0%
#545885000000
1!
1%
#545890000000
0!
0%
#545895000000
1!
1%
#545900000000
0!
0%
#545905000000
1!
1%
#545910000000
0!
0%
#545915000000
1!
1%
#545920000000
0!
0%
#545925000000
1!
1%
#545930000000
0!
0%
#545935000000
1!
1%
#545940000000
0!
0%
#545945000000
1!
1%
#545950000000
0!
0%
#545955000000
1!
1%
#545960000000
0!
0%
#545965000000
1!
1%
#545970000000
0!
0%
#545975000000
1!
1%
#545980000000
0!
0%
#545985000000
1!
1%
#545990000000
0!
0%
#545995000000
1!
1%
#546000000000
0!
0%
#546005000000
1!
1%
#546010000000
0!
0%
#546015000000
1!
1%
#546020000000
0!
0%
#546025000000
1!
1%
#546030000000
0!
0%
#546035000000
1!
1%
#546040000000
0!
0%
#546045000000
1!
1%
#546050000000
0!
0%
#546055000000
1!
1%
#546060000000
0!
0%
#546065000000
1!
1%
#546070000000
0!
0%
#546075000000
1!
1%
#546080000000
0!
0%
#546085000000
1!
1%
#546090000000
0!
0%
#546095000000
1!
1%
#546100000000
0!
0%
#546105000000
1!
1%
#546110000000
0!
0%
#546115000000
1!
1%
#546120000000
0!
0%
#546125000000
1!
1%
#546130000000
0!
0%
#546135000000
1!
1%
#546140000000
0!
0%
#546145000000
1!
1%
#546150000000
0!
0%
#546155000000
1!
1%
#546160000000
0!
0%
#546165000000
1!
1%
#546170000000
0!
0%
#546175000000
1!
1%
#546180000000
0!
0%
#546185000000
1!
1%
#546190000000
0!
0%
#546195000000
1!
1%
#546200000000
0!
0%
#546205000000
1!
1%
#546210000000
0!
0%
#546215000000
1!
1%
#546220000000
0!
0%
#546225000000
1!
1%
#546230000000
0!
0%
#546235000000
1!
1%
#546240000000
0!
0%
#546245000000
1!
1%
#546250000000
0!
0%
#546255000000
1!
1%
#546260000000
0!
0%
#546265000000
1!
1%
#546270000000
0!
0%
#546275000000
1!
1%
#546280000000
0!
0%
#546285000000
1!
1%
#546290000000
0!
0%
#546295000000
1!
1%
#546300000000
0!
0%
#546305000000
1!
1%
#546310000000
0!
0%
#546315000000
1!
1%
#546320000000
0!
0%
#546325000000
1!
1%
#546330000000
0!
0%
#546335000000
1!
1%
#546340000000
0!
0%
#546345000000
1!
1%
#546350000000
0!
0%
#546355000000
1!
1%
#546360000000
0!
0%
#546365000000
1!
1%
#546370000000
0!
0%
#546375000000
1!
1%
#546380000000
0!
0%
#546385000000
1!
1%
#546390000000
0!
0%
#546395000000
1!
1%
#546400000000
0!
0%
#546405000000
1!
1%
#546410000000
0!
0%
#546415000000
1!
1%
#546420000000
0!
0%
#546425000000
1!
1%
#546430000000
0!
0%
#546435000000
1!
1%
#546440000000
0!
0%
#546445000000
1!
1%
#546450000000
0!
0%
#546455000000
1!
1%
#546460000000
0!
0%
#546465000000
1!
1%
#546470000000
0!
0%
#546475000000
1!
1%
#546480000000
0!
0%
#546485000000
1!
1%
#546490000000
0!
0%
#546495000000
1!
1%
#546500000000
0!
0%
#546505000000
1!
1%
#546510000000
0!
0%
#546515000000
1!
1%
#546520000000
0!
0%
#546525000000
1!
1%
#546530000000
0!
0%
#546535000000
1!
1%
#546540000000
0!
0%
#546545000000
1!
1%
#546550000000
0!
0%
#546555000000
1!
1%
#546560000000
0!
0%
#546565000000
1!
1%
#546570000000
0!
0%
#546575000000
1!
1%
#546580000000
0!
0%
#546585000000
1!
1%
#546590000000
0!
0%
#546595000000
1!
1%
#546600000000
0!
0%
#546605000000
1!
1%
#546610000000
0!
0%
#546615000000
1!
1%
#546620000000
0!
0%
#546625000000
1!
1%
#546630000000
0!
0%
#546635000000
1!
1%
#546640000000
0!
0%
#546645000000
1!
1%
#546650000000
0!
0%
#546655000000
1!
1%
#546660000000
0!
0%
#546665000000
1!
1%
#546670000000
0!
0%
#546675000000
1!
1%
#546680000000
0!
0%
#546685000000
1!
1%
#546690000000
0!
0%
#546695000000
1!
1%
#546700000000
0!
0%
#546705000000
1!
1%
#546710000000
0!
0%
#546715000000
1!
1%
#546720000000
0!
0%
#546725000000
1!
1%
#546730000000
0!
0%
#546735000000
1!
1%
#546740000000
0!
0%
#546745000000
1!
1%
#546750000000
0!
0%
#546755000000
1!
1%
#546760000000
0!
0%
#546765000000
1!
1%
#546770000000
0!
0%
#546775000000
1!
1%
#546780000000
0!
0%
#546785000000
1!
1%
#546790000000
0!
0%
#546795000000
1!
1%
#546800000000
0!
0%
#546805000000
1!
1%
#546810000000
0!
0%
#546815000000
1!
1%
#546820000000
0!
0%
#546825000000
1!
1%
#546830000000
0!
0%
#546835000000
1!
1%
#546840000000
0!
0%
#546845000000
1!
1%
#546850000000
0!
0%
#546855000000
1!
1%
#546860000000
0!
0%
#546865000000
1!
1%
#546870000000
0!
0%
#546875000000
1!
1%
#546880000000
0!
0%
#546885000000
1!
1%
#546890000000
0!
0%
#546895000000
1!
1%
#546900000000
0!
0%
#546905000000
1!
1%
#546910000000
0!
0%
#546915000000
1!
1%
#546920000000
0!
0%
#546925000000
1!
1%
#546930000000
0!
0%
#546935000000
1!
1%
#546940000000
0!
0%
#546945000000
1!
1%
#546950000000
0!
0%
#546955000000
1!
1%
#546960000000
0!
0%
#546965000000
1!
1%
#546970000000
0!
0%
#546975000000
1!
1%
#546980000000
0!
0%
#546985000000
1!
1%
#546990000000
0!
0%
#546995000000
1!
1%
#547000000000
0!
0%
#547005000000
1!
1%
#547010000000
0!
0%
#547015000000
1!
1%
#547020000000
0!
0%
#547025000000
1!
1%
#547030000000
0!
0%
#547035000000
1!
1%
#547040000000
0!
0%
#547045000000
1!
1%
#547050000000
0!
0%
#547055000000
1!
1%
#547060000000
0!
0%
#547065000000
1!
1%
#547070000000
0!
0%
#547075000000
1!
1%
#547080000000
0!
0%
#547085000000
1!
1%
#547090000000
0!
0%
#547095000000
1!
1%
#547100000000
0!
0%
#547105000000
1!
1%
#547110000000
0!
0%
#547115000000
1!
1%
#547120000000
0!
0%
#547125000000
1!
1%
#547130000000
0!
0%
#547135000000
1!
1%
#547140000000
0!
0%
#547145000000
1!
1%
#547150000000
0!
0%
#547155000000
1!
1%
#547160000000
0!
0%
#547165000000
1!
1%
#547170000000
0!
0%
#547175000000
1!
1%
#547180000000
0!
0%
#547185000000
1!
1%
#547190000000
0!
0%
#547195000000
1!
1%
#547200000000
0!
0%
#547205000000
1!
1%
#547210000000
0!
0%
#547215000000
1!
1%
#547220000000
0!
0%
#547225000000
1!
1%
#547230000000
0!
0%
#547235000000
1!
1%
#547240000000
0!
0%
#547245000000
1!
1%
#547250000000
0!
0%
#547255000000
1!
1%
#547260000000
0!
0%
#547265000000
1!
1%
#547270000000
0!
0%
#547275000000
1!
1%
#547280000000
0!
0%
#547285000000
1!
1%
#547290000000
0!
0%
#547295000000
1!
1%
#547300000000
0!
0%
#547305000000
1!
1%
#547310000000
0!
0%
#547315000000
1!
1%
#547320000000
0!
0%
#547325000000
1!
1%
#547330000000
0!
0%
#547335000000
1!
1%
#547340000000
0!
0%
#547345000000
1!
1%
#547350000000
0!
0%
#547355000000
1!
1%
#547360000000
0!
0%
#547365000000
1!
1%
#547370000000
0!
0%
#547375000000
1!
1%
#547380000000
0!
0%
#547385000000
1!
1%
#547390000000
0!
0%
#547395000000
1!
1%
#547400000000
0!
0%
#547405000000
1!
1%
#547410000000
0!
0%
#547415000000
1!
1%
#547420000000
0!
0%
#547425000000
1!
1%
#547430000000
0!
0%
#547435000000
1!
1%
#547440000000
0!
0%
#547445000000
1!
1%
#547450000000
0!
0%
#547455000000
1!
1%
#547460000000
0!
0%
#547465000000
1!
1%
#547470000000
0!
0%
#547475000000
1!
1%
#547480000000
0!
0%
#547485000000
1!
1%
#547490000000
0!
0%
#547495000000
1!
1%
#547500000000
0!
0%
#547505000000
1!
1%
#547510000000
0!
0%
#547515000000
1!
1%
#547520000000
0!
0%
#547525000000
1!
1%
#547530000000
0!
0%
#547535000000
1!
1%
#547540000000
0!
0%
#547545000000
1!
1%
#547550000000
0!
0%
#547555000000
1!
1%
#547560000000
0!
0%
#547565000000
1!
1%
#547570000000
0!
0%
#547575000000
1!
1%
#547580000000
0!
0%
#547585000000
1!
1%
#547590000000
0!
0%
#547595000000
1!
1%
#547600000000
0!
0%
#547605000000
1!
1%
#547610000000
0!
0%
#547615000000
1!
1%
#547620000000
0!
0%
#547625000000
1!
1%
#547630000000
0!
0%
#547635000000
1!
1%
#547640000000
0!
0%
#547645000000
1!
1%
#547650000000
0!
0%
#547655000000
1!
1%
#547660000000
0!
0%
#547665000000
1!
1%
#547670000000
0!
0%
#547675000000
1!
1%
#547680000000
0!
0%
#547685000000
1!
1%
#547690000000
0!
0%
#547695000000
1!
1%
#547700000000
0!
0%
#547705000000
1!
1%
#547710000000
0!
0%
#547715000000
1!
1%
#547720000000
0!
0%
#547725000000
1!
1%
#547730000000
0!
0%
#547735000000
1!
1%
#547740000000
0!
0%
#547745000000
1!
1%
#547750000000
0!
0%
#547755000000
1!
1%
#547760000000
0!
0%
#547765000000
1!
1%
#547770000000
0!
0%
#547775000000
1!
1%
#547780000000
0!
0%
#547785000000
1!
1%
#547790000000
0!
0%
#547795000000
1!
1%
#547800000000
0!
0%
#547805000000
1!
1%
#547810000000
0!
0%
#547815000000
1!
1%
#547820000000
0!
0%
#547825000000
1!
1%
#547830000000
0!
0%
#547835000000
1!
1%
#547840000000
0!
0%
#547845000000
1!
1%
#547850000000
0!
0%
#547855000000
1!
1%
#547860000000
0!
0%
#547865000000
1!
1%
#547870000000
0!
0%
#547875000000
1!
1%
#547880000000
0!
0%
#547885000000
1!
1%
#547890000000
0!
0%
#547895000000
1!
1%
#547900000000
0!
0%
#547905000000
1!
1%
#547910000000
0!
0%
#547915000000
1!
1%
#547920000000
0!
0%
#547925000000
1!
1%
#547930000000
0!
0%
#547935000000
1!
1%
#547940000000
0!
0%
#547945000000
1!
1%
#547950000000
0!
0%
#547955000000
1!
1%
#547960000000
0!
0%
#547965000000
1!
1%
#547970000000
0!
0%
#547975000000
1!
1%
#547980000000
0!
0%
#547985000000
1!
1%
#547990000000
0!
0%
#547995000000
1!
1%
#548000000000
0!
0%
#548005000000
1!
1%
#548010000000
0!
0%
#548015000000
1!
1%
#548020000000
0!
0%
#548025000000
1!
1%
#548030000000
0!
0%
#548035000000
1!
1%
#548040000000
0!
0%
#548045000000
1!
1%
#548050000000
0!
0%
#548055000000
1!
1%
#548060000000
0!
0%
#548065000000
1!
1%
#548070000000
0!
0%
#548075000000
1!
1%
#548080000000
0!
0%
#548085000000
1!
1%
#548090000000
0!
0%
#548095000000
1!
1%
#548100000000
0!
0%
#548105000000
1!
1%
#548110000000
0!
0%
#548115000000
1!
1%
#548120000000
0!
0%
#548125000000
1!
1%
#548130000000
0!
0%
#548135000000
1!
1%
#548140000000
0!
0%
#548145000000
1!
1%
#548150000000
0!
0%
#548155000000
1!
1%
#548160000000
0!
0%
#548165000000
1!
1%
#548170000000
0!
0%
#548175000000
1!
1%
#548180000000
0!
0%
#548185000000
1!
1%
#548190000000
0!
0%
#548195000000
1!
1%
#548200000000
0!
0%
#548205000000
1!
1%
#548210000000
0!
0%
#548215000000
1!
1%
#548220000000
0!
0%
#548225000000
1!
1%
#548230000000
0!
0%
#548235000000
1!
1%
#548240000000
0!
0%
#548245000000
1!
1%
#548250000000
0!
0%
#548255000000
1!
1%
#548260000000
0!
0%
#548265000000
1!
1%
#548270000000
0!
0%
#548275000000
1!
1%
#548280000000
0!
0%
#548285000000
1!
1%
#548290000000
0!
0%
#548295000000
1!
1%
#548300000000
0!
0%
#548305000000
1!
1%
#548310000000
0!
0%
#548315000000
1!
1%
#548320000000
0!
0%
#548325000000
1!
1%
#548330000000
0!
0%
#548335000000
1!
1%
#548340000000
0!
0%
#548345000000
1!
1%
#548350000000
0!
0%
#548355000000
1!
1%
#548360000000
0!
0%
#548365000000
1!
1%
#548370000000
0!
0%
#548375000000
1!
1%
#548380000000
0!
0%
#548385000000
1!
1%
#548390000000
0!
0%
#548395000000
1!
1%
#548400000000
0!
0%
#548405000000
1!
1%
#548410000000
0!
0%
#548415000000
1!
1%
#548420000000
0!
0%
#548425000000
1!
1%
#548430000000
0!
0%
#548435000000
1!
1%
#548440000000
0!
0%
#548445000000
1!
1%
#548450000000
0!
0%
#548455000000
1!
1%
#548460000000
0!
0%
#548465000000
1!
1%
#548470000000
0!
0%
#548475000000
1!
1%
#548480000000
0!
0%
#548485000000
1!
1%
#548490000000
0!
0%
#548495000000
1!
1%
#548500000000
0!
0%
#548505000000
1!
1%
#548510000000
0!
0%
#548515000000
1!
1%
#548520000000
0!
0%
#548525000000
1!
1%
#548530000000
0!
0%
#548535000000
1!
1%
#548540000000
0!
0%
#548545000000
1!
1%
#548550000000
0!
0%
#548555000000
1!
1%
#548560000000
0!
0%
#548565000000
1!
1%
#548570000000
0!
0%
#548575000000
1!
1%
#548580000000
0!
0%
#548585000000
1!
1%
#548590000000
0!
0%
#548595000000
1!
1%
#548600000000
0!
0%
#548605000000
1!
1%
#548610000000
0!
0%
#548615000000
1!
1%
#548620000000
0!
0%
#548625000000
1!
1%
#548630000000
0!
0%
#548635000000
1!
1%
#548640000000
0!
0%
#548645000000
1!
1%
#548650000000
0!
0%
#548655000000
1!
1%
#548660000000
0!
0%
#548665000000
1!
1%
#548670000000
0!
0%
#548675000000
1!
1%
#548680000000
0!
0%
#548685000000
1!
1%
#548690000000
0!
0%
#548695000000
1!
1%
#548700000000
0!
0%
#548705000000
1!
1%
#548710000000
0!
0%
#548715000000
1!
1%
#548720000000
0!
0%
#548725000000
1!
1%
#548730000000
0!
0%
#548735000000
1!
1%
#548740000000
0!
0%
#548745000000
1!
1%
#548750000000
0!
0%
#548755000000
1!
1%
#548760000000
0!
0%
#548765000000
1!
1%
#548770000000
0!
0%
#548775000000
1!
1%
#548780000000
0!
0%
#548785000000
1!
1%
#548790000000
0!
0%
#548795000000
1!
1%
#548800000000
0!
0%
#548805000000
1!
1%
#548810000000
0!
0%
#548815000000
1!
1%
#548820000000
0!
0%
#548825000000
1!
1%
#548830000000
0!
0%
#548835000000
1!
1%
#548840000000
0!
0%
#548845000000
1!
1%
#548850000000
0!
0%
#548855000000
1!
1%
#548860000000
0!
0%
#548865000000
1!
1%
#548870000000
0!
0%
#548875000000
1!
1%
#548880000000
0!
0%
#548885000000
1!
1%
#548890000000
0!
0%
#548895000000
1!
1%
#548900000000
0!
0%
#548905000000
1!
1%
#548910000000
0!
0%
#548915000000
1!
1%
#548920000000
0!
0%
#548925000000
1!
1%
#548930000000
0!
0%
#548935000000
1!
1%
#548940000000
0!
0%
#548945000000
1!
1%
#548950000000
0!
0%
#548955000000
1!
1%
#548960000000
0!
0%
#548965000000
1!
1%
#548970000000
0!
0%
#548975000000
1!
1%
#548980000000
0!
0%
#548985000000
1!
1%
#548990000000
0!
0%
#548995000000
1!
1%
#549000000000
0!
0%
#549005000000
1!
1%
#549010000000
0!
0%
#549015000000
1!
1%
#549020000000
0!
0%
#549025000000
1!
1%
#549030000000
0!
0%
#549035000000
1!
1%
#549040000000
0!
0%
#549045000000
1!
1%
#549050000000
0!
0%
#549055000000
1!
1%
#549060000000
0!
0%
#549065000000
1!
1%
#549070000000
0!
0%
#549075000000
1!
1%
#549080000000
0!
0%
#549085000000
1!
1%
#549090000000
0!
0%
#549095000000
1!
1%
#549100000000
0!
0%
#549105000000
1!
1%
#549110000000
0!
0%
#549115000000
1!
1%
#549120000000
0!
0%
#549125000000
1!
1%
#549130000000
0!
0%
#549135000000
1!
1%
#549140000000
0!
0%
#549145000000
1!
1%
#549150000000
0!
0%
#549155000000
1!
1%
#549160000000
0!
0%
#549165000000
1!
1%
#549170000000
0!
0%
#549175000000
1!
1%
#549180000000
0!
0%
#549185000000
1!
1%
#549190000000
0!
0%
#549195000000
1!
1%
#549200000000
0!
0%
#549205000000
1!
1%
#549210000000
0!
0%
#549215000000
1!
1%
#549220000000
0!
0%
#549225000000
1!
1%
#549230000000
0!
0%
#549235000000
1!
1%
#549240000000
0!
0%
#549245000000
1!
1%
#549250000000
0!
0%
#549255000000
1!
1%
#549260000000
0!
0%
#549265000000
1!
1%
#549270000000
0!
0%
#549275000000
1!
1%
#549280000000
0!
0%
#549285000000
1!
1%
#549290000000
0!
0%
#549295000000
1!
1%
#549300000000
0!
0%
#549305000000
1!
1%
#549310000000
0!
0%
#549315000000
1!
1%
#549320000000
0!
0%
#549325000000
1!
1%
#549330000000
0!
0%
#549335000000
1!
1%
#549340000000
0!
0%
#549345000000
1!
1%
#549350000000
0!
0%
#549355000000
1!
1%
#549360000000
0!
0%
#549365000000
1!
1%
#549370000000
0!
0%
#549375000000
1!
1%
#549380000000
0!
0%
#549385000000
1!
1%
#549390000000
0!
0%
#549395000000
1!
1%
#549400000000
0!
0%
#549405000000
1!
1%
#549410000000
0!
0%
#549415000000
1!
1%
#549420000000
0!
0%
#549425000000
1!
1%
#549430000000
0!
0%
#549435000000
1!
1%
#549440000000
0!
0%
#549445000000
1!
1%
#549450000000
0!
0%
#549455000000
1!
1%
#549460000000
0!
0%
#549465000000
1!
1%
#549470000000
0!
0%
#549475000000
1!
1%
#549480000000
0!
0%
#549485000000
1!
1%
#549490000000
0!
0%
#549495000000
1!
1%
#549500000000
0!
0%
#549505000000
1!
1%
#549510000000
0!
0%
#549515000000
1!
1%
#549520000000
0!
0%
#549525000000
1!
1%
#549530000000
0!
0%
#549535000000
1!
1%
#549540000000
0!
0%
#549545000000
1!
1%
#549550000000
0!
0%
#549555000000
1!
1%
#549560000000
0!
0%
#549565000000
1!
1%
#549570000000
0!
0%
#549575000000
1!
1%
#549580000000
0!
0%
#549585000000
1!
1%
#549590000000
0!
0%
#549595000000
1!
1%
#549600000000
0!
0%
#549605000000
1!
1%
#549610000000
0!
0%
#549615000000
1!
1%
#549620000000
0!
0%
#549625000000
1!
1%
#549630000000
0!
0%
#549635000000
1!
1%
#549640000000
0!
0%
#549645000000
1!
1%
#549650000000
0!
0%
#549655000000
1!
1%
#549660000000
0!
0%
#549665000000
1!
1%
#549670000000
0!
0%
#549675000000
1!
1%
#549680000000
0!
0%
#549685000000
1!
1%
#549690000000
0!
0%
#549695000000
1!
1%
#549700000000
0!
0%
#549705000000
1!
1%
#549710000000
0!
0%
#549715000000
1!
1%
#549720000000
0!
0%
#549725000000
1!
1%
#549730000000
0!
0%
#549735000000
1!
1%
#549740000000
0!
0%
#549745000000
1!
1%
#549750000000
0!
0%
#549755000000
1!
1%
#549760000000
0!
0%
#549765000000
1!
1%
#549770000000
0!
0%
#549775000000
1!
1%
#549780000000
0!
0%
#549785000000
1!
1%
#549790000000
0!
0%
#549795000000
1!
1%
#549800000000
0!
0%
#549805000000
1!
1%
#549810000000
0!
0%
#549815000000
1!
1%
#549820000000
0!
0%
#549825000000
1!
1%
#549830000000
0!
0%
#549835000000
1!
1%
#549840000000
0!
0%
#549845000000
1!
1%
#549850000000
0!
0%
#549855000000
1!
1%
#549860000000
0!
0%
#549865000000
1!
1%
#549870000000
0!
0%
#549875000000
1!
1%
#549880000000
0!
0%
#549885000000
1!
1%
#549890000000
0!
0%
#549895000000
1!
1%
#549900000000
0!
0%
#549905000000
1!
1%
#549910000000
0!
0%
#549915000000
1!
1%
#549920000000
0!
0%
#549925000000
1!
1%
#549930000000
0!
0%
#549935000000
1!
1%
#549940000000
0!
0%
#549945000000
1!
1%
#549950000000
0!
0%
#549955000000
1!
1%
#549960000000
0!
0%
#549965000000
1!
1%
#549970000000
0!
0%
#549975000000
1!
1%
#549980000000
0!
0%
#549985000000
1!
1%
#549990000000
0!
0%
#549995000000
1!
1%
#550000000000
0!
0%
#550005000000
1!
1%
#550010000000
0!
0%
#550015000000
1!
1%
#550020000000
0!
0%
#550025000000
1!
1%
#550030000000
0!
0%
#550035000000
1!
1%
#550040000000
0!
0%
#550045000000
1!
1%
#550050000000
0!
0%
#550055000000
1!
1%
#550060000000
0!
0%
#550065000000
1!
1%
#550070000000
0!
0%
#550075000000
1!
1%
#550080000000
0!
0%
#550085000000
1!
1%
#550090000000
0!
0%
#550095000000
1!
1%
#550100000000
0!
0%
#550105000000
1!
1%
#550110000000
0!
0%
#550115000000
1!
1%
#550120000000
0!
0%
#550125000000
1!
1%
#550130000000
0!
0%
#550135000000
1!
1%
#550140000000
0!
0%
#550145000000
1!
1%
#550150000000
0!
0%
#550155000000
1!
1%
#550160000000
0!
0%
#550165000000
1!
1%
#550170000000
0!
0%
#550175000000
1!
1%
#550180000000
0!
0%
#550185000000
1!
1%
#550190000000
0!
0%
#550195000000
1!
1%
#550200000000
0!
0%
#550205000000
1!
1%
#550210000000
0!
0%
#550215000000
1!
1%
#550220000000
0!
0%
#550225000000
1!
1%
#550230000000
0!
0%
#550235000000
1!
1%
#550240000000
0!
0%
#550245000000
1!
1%
#550250000000
0!
0%
#550255000000
1!
1%
#550260000000
0!
0%
#550265000000
1!
1%
#550270000000
0!
0%
#550275000000
1!
1%
#550280000000
0!
0%
#550285000000
1!
1%
#550290000000
0!
0%
#550295000000
1!
1%
#550300000000
0!
0%
#550305000000
1!
1%
#550310000000
0!
0%
#550315000000
1!
1%
#550320000000
0!
0%
#550325000000
1!
1%
#550330000000
0!
0%
#550335000000
1!
1%
#550340000000
0!
0%
#550345000000
1!
1%
#550350000000
0!
0%
#550355000000
1!
1%
#550360000000
0!
0%
#550365000000
1!
1%
#550370000000
0!
0%
#550375000000
1!
1%
#550380000000
0!
0%
#550385000000
1!
1%
#550390000000
0!
0%
#550395000000
1!
1%
#550400000000
0!
0%
#550405000000
1!
1%
#550410000000
0!
0%
#550415000000
1!
1%
#550420000000
0!
0%
#550425000000
1!
1%
#550430000000
0!
0%
#550435000000
1!
1%
#550440000000
0!
0%
#550445000000
1!
1%
#550450000000
0!
0%
#550455000000
1!
1%
#550460000000
0!
0%
#550465000000
1!
1%
#550470000000
0!
0%
#550475000000
1!
1%
#550480000000
0!
0%
#550485000000
1!
1%
#550490000000
0!
0%
#550495000000
1!
1%
#550500000000
0!
0%
#550505000000
1!
1%
#550510000000
0!
0%
#550515000000
1!
1%
#550520000000
0!
0%
#550525000000
1!
1%
#550530000000
0!
0%
#550535000000
1!
1%
#550540000000
0!
0%
#550545000000
1!
1%
#550550000000
0!
0%
#550555000000
1!
1%
#550560000000
0!
0%
#550565000000
1!
1%
#550570000000
0!
0%
#550575000000
1!
1%
#550580000000
0!
0%
#550585000000
1!
1%
#550590000000
0!
0%
#550595000000
1!
1%
#550600000000
0!
0%
#550605000000
1!
1%
#550610000000
0!
0%
#550615000000
1!
1%
#550620000000
0!
0%
#550625000000
1!
1%
#550630000000
0!
0%
#550635000000
1!
1%
#550640000000
0!
0%
#550645000000
1!
1%
#550650000000
0!
0%
#550655000000
1!
1%
#550660000000
0!
0%
#550665000000
1!
1%
#550670000000
0!
0%
#550675000000
1!
1%
#550680000000
0!
0%
#550685000000
1!
1%
#550690000000
0!
0%
#550695000000
1!
1%
#550700000000
0!
0%
#550705000000
1!
1%
#550710000000
0!
0%
#550715000000
1!
1%
#550720000000
0!
0%
#550725000000
1!
1%
#550730000000
0!
0%
#550735000000
1!
1%
#550740000000
0!
0%
#550745000000
1!
1%
#550750000000
0!
0%
#550755000000
1!
1%
#550760000000
0!
0%
#550765000000
1!
1%
#550770000000
0!
0%
#550775000000
1!
1%
#550780000000
0!
0%
#550785000000
1!
1%
#550790000000
0!
0%
#550795000000
1!
1%
#550800000000
0!
0%
#550805000000
1!
1%
#550810000000
0!
0%
#550815000000
1!
1%
#550820000000
0!
0%
#550825000000
1!
1%
#550830000000
0!
0%
#550835000000
1!
1%
#550840000000
0!
0%
#550845000000
1!
1%
#550850000000
0!
0%
#550855000000
1!
1%
#550860000000
0!
0%
#550865000000
1!
1%
#550870000000
0!
0%
#550875000000
1!
1%
#550880000000
0!
0%
#550885000000
1!
1%
#550890000000
0!
0%
#550895000000
1!
1%
#550900000000
0!
0%
#550905000000
1!
1%
#550910000000
0!
0%
#550915000000
1!
1%
#550920000000
0!
0%
#550925000000
1!
1%
#550930000000
0!
0%
#550935000000
1!
1%
#550940000000
0!
0%
#550945000000
1!
1%
#550950000000
0!
0%
#550955000000
1!
1%
#550960000000
0!
0%
#550965000000
1!
1%
#550970000000
0!
0%
#550975000000
1!
1%
#550980000000
0!
0%
#550985000000
1!
1%
#550990000000
0!
0%
#550995000000
1!
1%
#551000000000
0!
0%
#551005000000
1!
1%
#551010000000
0!
0%
#551015000000
1!
1%
#551020000000
0!
0%
#551025000000
1!
1%
#551030000000
0!
0%
#551035000000
1!
1%
#551040000000
0!
0%
#551045000000
1!
1%
#551050000000
0!
0%
#551055000000
1!
1%
#551060000000
0!
0%
#551065000000
1!
1%
#551070000000
0!
0%
#551075000000
1!
1%
#551080000000
0!
0%
#551085000000
1!
1%
#551090000000
0!
0%
#551095000000
1!
1%
#551100000000
0!
0%
#551105000000
1!
1%
#551110000000
0!
0%
#551115000000
1!
1%
#551120000000
0!
0%
#551125000000
1!
1%
#551130000000
0!
0%
#551135000000
1!
1%
#551140000000
0!
0%
#551145000000
1!
1%
#551150000000
0!
0%
#551155000000
1!
1%
#551160000000
0!
0%
#551165000000
1!
1%
#551170000000
0!
0%
#551175000000
1!
1%
#551180000000
0!
0%
#551185000000
1!
1%
#551190000000
0!
0%
#551195000000
1!
1%
#551200000000
0!
0%
#551205000000
1!
1%
#551210000000
0!
0%
#551215000000
1!
1%
#551220000000
0!
0%
#551225000000
1!
1%
#551230000000
0!
0%
#551235000000
1!
1%
#551240000000
0!
0%
#551245000000
1!
1%
#551250000000
0!
0%
#551255000000
1!
1%
#551260000000
0!
0%
#551265000000
1!
1%
#551270000000
0!
0%
#551275000000
1!
1%
#551280000000
0!
0%
#551285000000
1!
1%
#551290000000
0!
0%
#551295000000
1!
1%
#551300000000
0!
0%
#551305000000
1!
1%
#551310000000
0!
0%
#551315000000
1!
1%
#551320000000
0!
0%
#551325000000
1!
1%
#551330000000
0!
0%
#551335000000
1!
1%
#551340000000
0!
0%
#551345000000
1!
1%
#551350000000
0!
0%
#551355000000
1!
1%
#551360000000
0!
0%
#551365000000
1!
1%
#551370000000
0!
0%
#551375000000
1!
1%
#551380000000
0!
0%
#551385000000
1!
1%
#551390000000
0!
0%
#551395000000
1!
1%
#551400000000
0!
0%
#551405000000
1!
1%
#551410000000
0!
0%
#551415000000
1!
1%
#551420000000
0!
0%
#551425000000
1!
1%
#551430000000
0!
0%
#551435000000
1!
1%
#551440000000
0!
0%
#551445000000
1!
1%
#551450000000
0!
0%
#551455000000
1!
1%
#551460000000
0!
0%
#551465000000
1!
1%
#551470000000
0!
0%
#551475000000
1!
1%
#551480000000
0!
0%
#551485000000
1!
1%
#551490000000
0!
0%
#551495000000
1!
1%
#551500000000
0!
0%
#551505000000
1!
1%
#551510000000
0!
0%
#551515000000
1!
1%
#551520000000
0!
0%
#551525000000
1!
1%
#551530000000
0!
0%
#551535000000
1!
1%
#551540000000
0!
0%
#551545000000
1!
1%
#551550000000
0!
0%
#551555000000
1!
1%
#551560000000
0!
0%
#551565000000
1!
1%
#551570000000
0!
0%
#551575000000
1!
1%
#551580000000
0!
0%
#551585000000
1!
1%
#551590000000
0!
0%
#551595000000
1!
1%
#551600000000
0!
0%
#551605000000
1!
1%
#551610000000
0!
0%
#551615000000
1!
1%
#551620000000
0!
0%
#551625000000
1!
1%
#551630000000
0!
0%
#551635000000
1!
1%
#551640000000
0!
0%
#551645000000
1!
1%
#551650000000
0!
0%
#551655000000
1!
1%
#551660000000
0!
0%
#551665000000
1!
1%
#551670000000
0!
0%
#551675000000
1!
1%
#551680000000
0!
0%
#551685000000
1!
1%
#551690000000
0!
0%
#551695000000
1!
1%
#551700000000
0!
0%
#551705000000
1!
1%
#551710000000
0!
0%
#551715000000
1!
1%
#551720000000
0!
0%
#551725000000
1!
1%
#551730000000
0!
0%
#551735000000
1!
1%
#551740000000
0!
0%
#551745000000
1!
1%
#551750000000
0!
0%
#551755000000
1!
1%
#551760000000
0!
0%
#551765000000
1!
1%
#551770000000
0!
0%
#551775000000
1!
1%
#551780000000
0!
0%
#551785000000
1!
1%
#551790000000
0!
0%
#551795000000
1!
1%
#551800000000
0!
0%
#551805000000
1!
1%
#551810000000
0!
0%
#551815000000
1!
1%
#551820000000
0!
0%
#551825000000
1!
1%
#551830000000
0!
0%
#551835000000
1!
1%
#551840000000
0!
0%
#551845000000
1!
1%
#551850000000
0!
0%
#551855000000
1!
1%
#551860000000
0!
0%
#551865000000
1!
1%
#551870000000
0!
0%
#551875000000
1!
1%
#551880000000
0!
0%
#551885000000
1!
1%
#551890000000
0!
0%
#551895000000
1!
1%
#551900000000
0!
0%
#551905000000
1!
1%
#551910000000
0!
0%
#551915000000
1!
1%
#551920000000
0!
0%
#551925000000
1!
1%
#551930000000
0!
0%
#551935000000
1!
1%
#551940000000
0!
0%
#551945000000
1!
1%
#551950000000
0!
0%
#551955000000
1!
1%
#551960000000
0!
0%
#551965000000
1!
1%
#551970000000
0!
0%
#551975000000
1!
1%
#551980000000
0!
0%
#551985000000
1!
1%
#551990000000
0!
0%
#551995000000
1!
1%
#552000000000
0!
0%
#552005000000
1!
1%
#552010000000
0!
0%
#552015000000
1!
1%
#552020000000
0!
0%
#552025000000
1!
1%
#552030000000
0!
0%
#552035000000
1!
1%
#552040000000
0!
0%
#552045000000
1!
1%
#552050000000
0!
0%
#552055000000
1!
1%
#552060000000
0!
0%
#552065000000
1!
1%
#552070000000
0!
0%
#552075000000
1!
1%
#552080000000
0!
0%
#552085000000
1!
1%
#552090000000
0!
0%
#552095000000
1!
1%
#552100000000
0!
0%
#552105000000
1!
1%
#552110000000
0!
0%
#552115000000
1!
1%
#552120000000
0!
0%
#552125000000
1!
1%
#552130000000
0!
0%
#552135000000
1!
1%
#552140000000
0!
0%
#552145000000
1!
1%
#552150000000
0!
0%
#552155000000
1!
1%
#552160000000
0!
0%
#552165000000
1!
1%
#552170000000
0!
0%
#552175000000
1!
1%
#552180000000
0!
0%
#552185000000
1!
1%
#552190000000
0!
0%
#552195000000
1!
1%
#552200000000
0!
0%
#552205000000
1!
1%
#552210000000
0!
0%
#552215000000
1!
1%
#552220000000
0!
0%
#552225000000
1!
1%
#552230000000
0!
0%
#552235000000
1!
1%
#552240000000
0!
0%
#552245000000
1!
1%
#552250000000
0!
0%
#552255000000
1!
1%
#552260000000
0!
0%
#552265000000
1!
1%
#552270000000
0!
0%
#552275000000
1!
1%
#552280000000
0!
0%
#552285000000
1!
1%
#552290000000
0!
0%
#552295000000
1!
1%
#552300000000
0!
0%
#552305000000
1!
1%
#552310000000
0!
0%
#552315000000
1!
1%
#552320000000
0!
0%
#552325000000
1!
1%
#552330000000
0!
0%
#552335000000
1!
1%
#552340000000
0!
0%
#552345000000
1!
1%
#552350000000
0!
0%
#552355000000
1!
1%
#552360000000
0!
0%
#552365000000
1!
1%
#552370000000
0!
0%
#552375000000
1!
1%
#552380000000
0!
0%
#552385000000
1!
1%
#552390000000
0!
0%
#552395000000
1!
1%
#552400000000
0!
0%
#552405000000
1!
1%
#552410000000
0!
0%
#552415000000
1!
1%
#552420000000
0!
0%
#552425000000
1!
1%
#552430000000
0!
0%
#552435000000
1!
1%
#552440000000
0!
0%
#552445000000
1!
1%
#552450000000
0!
0%
#552455000000
1!
1%
#552460000000
0!
0%
#552465000000
1!
1%
#552470000000
0!
0%
#552475000000
1!
1%
#552480000000
0!
0%
#552485000000
1!
1%
#552490000000
0!
0%
#552495000000
1!
1%
#552500000000
0!
0%
#552505000000
1!
1%
#552510000000
0!
0%
#552515000000
1!
1%
#552520000000
0!
0%
#552525000000
1!
1%
#552530000000
0!
0%
#552535000000
1!
1%
#552540000000
0!
0%
#552545000000
1!
1%
#552550000000
0!
0%
#552555000000
1!
1%
#552560000000
0!
0%
#552565000000
1!
1%
#552570000000
0!
0%
#552575000000
1!
1%
#552580000000
0!
0%
#552585000000
1!
1%
#552590000000
0!
0%
#552595000000
1!
1%
#552600000000
0!
0%
#552605000000
1!
1%
#552610000000
0!
0%
#552615000000
1!
1%
#552620000000
0!
0%
#552625000000
1!
1%
#552630000000
0!
0%
#552635000000
1!
1%
#552640000000
0!
0%
#552645000000
1!
1%
#552650000000
0!
0%
#552655000000
1!
1%
#552660000000
0!
0%
#552665000000
1!
1%
#552670000000
0!
0%
#552675000000
1!
1%
#552680000000
0!
0%
#552685000000
1!
1%
#552690000000
0!
0%
#552695000000
1!
1%
#552700000000
0!
0%
#552705000000
1!
1%
#552710000000
0!
0%
#552715000000
1!
1%
#552720000000
0!
0%
#552725000000
1!
1%
#552730000000
0!
0%
#552735000000
1!
1%
#552740000000
0!
0%
#552745000000
1!
1%
#552750000000
0!
0%
#552755000000
1!
1%
#552760000000
0!
0%
#552765000000
1!
1%
#552770000000
0!
0%
#552775000000
1!
1%
#552780000000
0!
0%
#552785000000
1!
1%
#552790000000
0!
0%
#552795000000
1!
1%
#552800000000
0!
0%
#552805000000
1!
1%
#552810000000
0!
0%
#552815000000
1!
1%
#552820000000
0!
0%
#552825000000
1!
1%
#552830000000
0!
0%
#552835000000
1!
1%
#552840000000
0!
0%
#552845000000
1!
1%
#552850000000
0!
0%
#552855000000
1!
1%
#552860000000
0!
0%
#552865000000
1!
1%
#552870000000
0!
0%
#552875000000
1!
1%
#552880000000
0!
0%
#552885000000
1!
1%
#552890000000
0!
0%
#552895000000
1!
1%
#552900000000
0!
0%
#552905000000
1!
1%
#552910000000
0!
0%
#552915000000
1!
1%
#552920000000
0!
0%
#552925000000
1!
1%
#552930000000
0!
0%
#552935000000
1!
1%
#552940000000
0!
0%
#552945000000
1!
1%
#552950000000
0!
0%
#552955000000
1!
1%
#552960000000
0!
0%
#552965000000
1!
1%
#552970000000
0!
0%
#552975000000
1!
1%
#552980000000
0!
0%
#552985000000
1!
1%
#552990000000
0!
0%
#552995000000
1!
1%
#553000000000
0!
0%
#553005000000
1!
1%
#553010000000
0!
0%
#553015000000
1!
1%
#553020000000
0!
0%
#553025000000
1!
1%
#553030000000
0!
0%
#553035000000
1!
1%
#553040000000
0!
0%
#553045000000
1!
1%
#553050000000
0!
0%
#553055000000
1!
1%
#553060000000
0!
0%
#553065000000
1!
1%
#553070000000
0!
0%
#553075000000
1!
1%
#553080000000
0!
0%
#553085000000
1!
1%
#553090000000
0!
0%
#553095000000
1!
1%
#553100000000
0!
0%
#553105000000
1!
1%
#553110000000
0!
0%
#553115000000
1!
1%
#553120000000
0!
0%
#553125000000
1!
1%
#553130000000
0!
0%
#553135000000
1!
1%
#553140000000
0!
0%
#553145000000
1!
1%
#553150000000
0!
0%
#553155000000
1!
1%
#553160000000
0!
0%
#553165000000
1!
1%
#553170000000
0!
0%
#553175000000
1!
1%
#553180000000
0!
0%
#553185000000
1!
1%
#553190000000
0!
0%
#553195000000
1!
1%
#553200000000
0!
0%
#553205000000
1!
1%
#553210000000
0!
0%
#553215000000
1!
1%
#553220000000
0!
0%
#553225000000
1!
1%
#553230000000
0!
0%
#553235000000
1!
1%
#553240000000
0!
0%
#553245000000
1!
1%
#553250000000
0!
0%
#553255000000
1!
1%
#553260000000
0!
0%
#553265000000
1!
1%
#553270000000
0!
0%
#553275000000
1!
1%
#553280000000
0!
0%
#553285000000
1!
1%
#553290000000
0!
0%
#553295000000
1!
1%
#553300000000
0!
0%
#553305000000
1!
1%
#553310000000
0!
0%
#553315000000
1!
1%
#553320000000
0!
0%
#553325000000
1!
1%
#553330000000
0!
0%
#553335000000
1!
1%
#553340000000
0!
0%
#553345000000
1!
1%
#553350000000
0!
0%
#553355000000
1!
1%
#553360000000
0!
0%
#553365000000
1!
1%
#553370000000
0!
0%
#553375000000
1!
1%
#553380000000
0!
0%
#553385000000
1!
1%
#553390000000
0!
0%
#553395000000
1!
1%
#553400000000
0!
0%
#553405000000
1!
1%
#553410000000
0!
0%
#553415000000
1!
1%
#553420000000
0!
0%
#553425000000
1!
1%
#553430000000
0!
0%
#553435000000
1!
1%
#553440000000
0!
0%
#553445000000
1!
1%
#553450000000
0!
0%
#553455000000
1!
1%
#553460000000
0!
0%
#553465000000
1!
1%
#553470000000
0!
0%
#553475000000
1!
1%
#553480000000
0!
0%
#553485000000
1!
1%
#553490000000
0!
0%
#553495000000
1!
1%
#553500000000
0!
0%
#553505000000
1!
1%
#553510000000
0!
0%
#553515000000
1!
1%
#553520000000
0!
0%
#553525000000
1!
1%
#553530000000
0!
0%
#553535000000
1!
1%
#553540000000
0!
0%
#553545000000
1!
1%
#553550000000
0!
0%
#553555000000
1!
1%
#553560000000
0!
0%
#553565000000
1!
1%
#553570000000
0!
0%
#553575000000
1!
1%
#553580000000
0!
0%
#553585000000
1!
1%
#553590000000
0!
0%
#553595000000
1!
1%
#553600000000
0!
0%
#553605000000
1!
1%
#553610000000
0!
0%
#553615000000
1!
1%
#553620000000
0!
0%
#553625000000
1!
1%
#553630000000
0!
0%
#553635000000
1!
1%
#553640000000
0!
0%
#553645000000
1!
1%
#553650000000
0!
0%
#553655000000
1!
1%
#553660000000
0!
0%
#553665000000
1!
1%
#553670000000
0!
0%
#553675000000
1!
1%
#553680000000
0!
0%
#553685000000
1!
1%
#553690000000
0!
0%
#553695000000
1!
1%
#553700000000
0!
0%
#553705000000
1!
1%
#553710000000
0!
0%
#553715000000
1!
1%
#553720000000
0!
0%
#553725000000
1!
1%
#553730000000
0!
0%
#553735000000
1!
1%
#553740000000
0!
0%
#553745000000
1!
1%
#553750000000
0!
0%
#553755000000
1!
1%
#553760000000
0!
0%
#553765000000
1!
1%
#553770000000
0!
0%
#553775000000
1!
1%
#553780000000
0!
0%
#553785000000
1!
1%
#553790000000
0!
0%
#553795000000
1!
1%
#553800000000
0!
0%
#553805000000
1!
1%
#553810000000
0!
0%
#553815000000
1!
1%
#553820000000
0!
0%
#553825000000
1!
1%
#553830000000
0!
0%
#553835000000
1!
1%
#553840000000
0!
0%
#553845000000
1!
1%
#553850000000
0!
0%
#553855000000
1!
1%
#553860000000
0!
0%
#553865000000
1!
1%
#553870000000
0!
0%
#553875000000
1!
1%
#553880000000
0!
0%
#553885000000
1!
1%
#553890000000
0!
0%
#553895000000
1!
1%
#553900000000
0!
0%
#553905000000
1!
1%
#553910000000
0!
0%
#553915000000
1!
1%
#553920000000
0!
0%
#553925000000
1!
1%
#553930000000
0!
0%
#553935000000
1!
1%
#553940000000
0!
0%
#553945000000
1!
1%
#553950000000
0!
0%
#553955000000
1!
1%
#553960000000
0!
0%
#553965000000
1!
1%
#553970000000
0!
0%
#553975000000
1!
1%
#553980000000
0!
0%
#553985000000
1!
1%
#553990000000
0!
0%
#553995000000
1!
1%
#554000000000
0!
0%
#554005000000
1!
1%
#554010000000
0!
0%
#554015000000
1!
1%
#554020000000
0!
0%
#554025000000
1!
1%
#554030000000
0!
0%
#554035000000
1!
1%
#554040000000
0!
0%
#554045000000
1!
1%
#554050000000
0!
0%
#554055000000
1!
1%
#554060000000
0!
0%
#554065000000
1!
1%
#554070000000
0!
0%
#554075000000
1!
1%
#554080000000
0!
0%
#554085000000
1!
1%
#554090000000
0!
0%
#554095000000
1!
1%
#554100000000
0!
0%
#554105000000
1!
1%
#554110000000
0!
0%
#554115000000
1!
1%
#554120000000
0!
0%
#554125000000
1!
1%
#554130000000
0!
0%
#554135000000
1!
1%
#554140000000
0!
0%
#554145000000
1!
1%
#554150000000
0!
0%
#554155000000
1!
1%
#554160000000
0!
0%
#554165000000
1!
1%
#554170000000
0!
0%
#554175000000
1!
1%
#554180000000
0!
0%
#554185000000
1!
1%
#554190000000
0!
0%
#554195000000
1!
1%
#554200000000
0!
0%
#554205000000
1!
1%
#554210000000
0!
0%
#554215000000
1!
1%
#554220000000
0!
0%
#554225000000
1!
1%
#554230000000
0!
0%
#554235000000
1!
1%
#554240000000
0!
0%
#554245000000
1!
1%
#554250000000
0!
0%
#554255000000
1!
1%
#554260000000
0!
0%
#554265000000
1!
1%
#554270000000
0!
0%
#554275000000
1!
1%
#554280000000
0!
0%
#554285000000
1!
1%
#554290000000
0!
0%
#554295000000
1!
1%
#554300000000
0!
0%
#554305000000
1!
1%
#554310000000
0!
0%
#554315000000
1!
1%
#554320000000
0!
0%
#554325000000
1!
1%
#554330000000
0!
0%
#554335000000
1!
1%
#554340000000
0!
0%
#554345000000
1!
1%
#554350000000
0!
0%
#554355000000
1!
1%
#554360000000
0!
0%
#554365000000
1!
1%
#554370000000
0!
0%
#554375000000
1!
1%
#554380000000
0!
0%
#554385000000
1!
1%
#554390000000
0!
0%
#554395000000
1!
1%
#554400000000
0!
0%
#554405000000
1!
1%
#554410000000
0!
0%
#554415000000
1!
1%
#554420000000
0!
0%
#554425000000
1!
1%
#554430000000
0!
0%
#554435000000
1!
1%
#554440000000
0!
0%
#554445000000
1!
1%
#554450000000
0!
0%
#554455000000
1!
1%
#554460000000
0!
0%
#554465000000
1!
1%
#554470000000
0!
0%
#554475000000
1!
1%
#554480000000
0!
0%
#554485000000
1!
1%
#554490000000
0!
0%
#554495000000
1!
1%
#554500000000
0!
0%
#554505000000
1!
1%
#554510000000
0!
0%
#554515000000
1!
1%
#554520000000
0!
0%
#554525000000
1!
1%
#554530000000
0!
0%
#554535000000
1!
1%
#554540000000
0!
0%
#554545000000
1!
1%
#554550000000
0!
0%
#554555000000
1!
1%
#554560000000
0!
0%
#554565000000
1!
1%
#554570000000
0!
0%
#554575000000
1!
1%
#554580000000
0!
0%
#554585000000
1!
1%
#554590000000
0!
0%
#554595000000
1!
1%
#554600000000
0!
0%
#554605000000
1!
1%
#554610000000
0!
0%
#554615000000
1!
1%
#554620000000
0!
0%
#554625000000
1!
1%
#554630000000
0!
0%
#554635000000
1!
1%
#554640000000
0!
0%
#554645000000
1!
1%
#554650000000
0!
0%
#554655000000
1!
1%
#554660000000
0!
0%
#554665000000
1!
1%
#554670000000
0!
0%
#554675000000
1!
1%
#554680000000
0!
0%
#554685000000
1!
1%
#554690000000
0!
0%
#554695000000
1!
1%
#554700000000
0!
0%
#554705000000
1!
1%
#554710000000
0!
0%
#554715000000
1!
1%
#554720000000
0!
0%
#554725000000
1!
1%
#554730000000
0!
0%
#554735000000
1!
1%
#554740000000
0!
0%
#554745000000
1!
1%
#554750000000
0!
0%
#554755000000
1!
1%
#554760000000
0!
0%
#554765000000
1!
1%
#554770000000
0!
0%
#554775000000
1!
1%
#554780000000
0!
0%
#554785000000
1!
1%
#554790000000
0!
0%
#554795000000
1!
1%
#554800000000
0!
0%
#554805000000
1!
1%
#554810000000
0!
0%
#554815000000
1!
1%
#554820000000
0!
0%
#554825000000
1!
1%
#554830000000
0!
0%
#554835000000
1!
1%
#554840000000
0!
0%
#554845000000
1!
1%
#554850000000
0!
0%
#554855000000
1!
1%
#554860000000
0!
0%
#554865000000
1!
1%
#554870000000
0!
0%
#554875000000
1!
1%
#554880000000
0!
0%
#554885000000
1!
1%
#554890000000
0!
0%
#554895000000
1!
1%
#554900000000
0!
0%
#554905000000
1!
1%
#554910000000
0!
0%
#554915000000
1!
1%
#554920000000
0!
0%
#554925000000
1!
1%
#554930000000
0!
0%
#554935000000
1!
1%
#554940000000
0!
0%
#554945000000
1!
1%
#554950000000
0!
0%
#554955000000
1!
1%
#554960000000
0!
0%
#554965000000
1!
1%
#554970000000
0!
0%
#554975000000
1!
1%
#554980000000
0!
0%
#554985000000
1!
1%
#554990000000
0!
0%
#554995000000
1!
1%
#555000000000
0!
0%
#555005000000
1!
1%
#555010000000
0!
0%
#555015000000
1!
1%
#555020000000
0!
0%
#555025000000
1!
1%
#555030000000
0!
0%
#555035000000
1!
1%
#555040000000
0!
0%
#555045000000
1!
1%
#555050000000
0!
0%
#555055000000
1!
1%
#555060000000
0!
0%
#555065000000
1!
1%
#555070000000
0!
0%
#555075000000
1!
1%
#555080000000
0!
0%
#555085000000
1!
1%
#555090000000
0!
0%
#555095000000
1!
1%
#555100000000
0!
0%
#555105000000
1!
1%
#555110000000
0!
0%
#555115000000
1!
1%
#555120000000
0!
0%
#555125000000
1!
1%
#555130000000
0!
0%
#555135000000
1!
1%
#555140000000
0!
0%
#555145000000
1!
1%
#555150000000
0!
0%
#555155000000
1!
1%
#555160000000
0!
0%
#555165000000
1!
1%
#555170000000
0!
0%
#555175000000
1!
1%
#555180000000
0!
0%
#555185000000
1!
1%
#555190000000
0!
0%
#555195000000
1!
1%
#555200000000
0!
0%
#555205000000
1!
1%
#555210000000
0!
0%
#555215000000
1!
1%
#555220000000
0!
0%
#555225000000
1!
1%
#555230000000
0!
0%
#555235000000
1!
1%
#555240000000
0!
0%
#555245000000
1!
1%
#555250000000
0!
0%
#555255000000
1!
1%
#555260000000
0!
0%
#555265000000
1!
1%
#555270000000
0!
0%
#555275000000
1!
1%
#555280000000
0!
0%
#555285000000
1!
1%
#555290000000
0!
0%
#555295000000
1!
1%
#555300000000
0!
0%
#555305000000
1!
1%
#555310000000
0!
0%
#555315000000
1!
1%
#555320000000
0!
0%
#555325000000
1!
1%
#555330000000
0!
0%
#555335000000
1!
1%
#555340000000
0!
0%
#555345000000
1!
1%
#555350000000
0!
0%
#555355000000
1!
1%
#555360000000
0!
0%
#555365000000
1!
1%
#555370000000
0!
0%
#555375000000
1!
1%
#555380000000
0!
0%
#555385000000
1!
1%
#555390000000
0!
0%
#555395000000
1!
1%
#555400000000
0!
0%
#555405000000
1!
1%
#555410000000
0!
0%
#555415000000
1!
1%
#555420000000
0!
0%
#555425000000
1!
1%
#555430000000
0!
0%
#555435000000
1!
1%
#555440000000
0!
0%
#555445000000
1!
1%
#555450000000
0!
0%
#555455000000
1!
1%
#555460000000
0!
0%
#555465000000
1!
1%
#555470000000
0!
0%
#555475000000
1!
1%
#555480000000
0!
0%
#555485000000
1!
1%
#555490000000
0!
0%
#555495000000
1!
1%
#555500000000
0!
0%
#555505000000
1!
1%
#555510000000
0!
0%
#555515000000
1!
1%
#555520000000
0!
0%
#555525000000
1!
1%
#555530000000
0!
0%
#555535000000
1!
1%
#555540000000
0!
0%
#555545000000
1!
1%
#555550000000
0!
0%
#555555000000
1!
1%
#555560000000
0!
0%
#555565000000
1!
1%
#555570000000
0!
0%
#555575000000
1!
1%
#555580000000
0!
0%
#555585000000
1!
1%
#555590000000
0!
0%
#555595000000
1!
1%
#555600000000
0!
0%
#555605000000
1!
1%
#555610000000
0!
0%
#555615000000
1!
1%
#555620000000
0!
0%
#555625000000
1!
1%
#555630000000
0!
0%
#555635000000
1!
1%
#555640000000
0!
0%
#555645000000
1!
1%
#555650000000
0!
0%
#555655000000
1!
1%
#555660000000
0!
0%
#555665000000
1!
1%
#555670000000
0!
0%
#555675000000
1!
1%
#555680000000
0!
0%
#555685000000
1!
1%
#555690000000
0!
0%
#555695000000
1!
1%
#555700000000
0!
0%
#555705000000
1!
1%
#555710000000
0!
0%
#555715000000
1!
1%
#555720000000
0!
0%
#555725000000
1!
1%
#555730000000
0!
0%
#555735000000
1!
1%
#555740000000
0!
0%
#555745000000
1!
1%
#555750000000
0!
0%
#555755000000
1!
1%
#555760000000
0!
0%
#555765000000
1!
1%
#555770000000
0!
0%
#555775000000
1!
1%
#555780000000
0!
0%
#555785000000
1!
1%
#555790000000
0!
0%
#555795000000
1!
1%
#555800000000
0!
0%
#555805000000
1!
1%
#555810000000
0!
0%
#555815000000
1!
1%
#555820000000
0!
0%
#555825000000
1!
1%
#555830000000
0!
0%
#555835000000
1!
1%
#555840000000
0!
0%
#555845000000
1!
1%
#555850000000
0!
0%
#555855000000
1!
1%
#555860000000
0!
0%
#555865000000
1!
1%
#555870000000
0!
0%
#555875000000
1!
1%
#555880000000
0!
0%
#555885000000
1!
1%
#555890000000
0!
0%
#555895000000
1!
1%
#555900000000
0!
0%
#555905000000
1!
1%
#555910000000
0!
0%
#555915000000
1!
1%
#555920000000
0!
0%
#555925000000
1!
1%
#555930000000
0!
0%
#555935000000
1!
1%
#555940000000
0!
0%
#555945000000
1!
1%
#555950000000
0!
0%
#555955000000
1!
1%
#555960000000
0!
0%
#555965000000
1!
1%
#555970000000
0!
0%
#555975000000
1!
1%
#555980000000
0!
0%
#555985000000
1!
1%
#555990000000
0!
0%
#555995000000
1!
1%
#556000000000
0!
0%
#556005000000
1!
1%
#556010000000
0!
0%
#556015000000
1!
1%
#556020000000
0!
0%
#556025000000
1!
1%
#556030000000
0!
0%
#556035000000
1!
1%
#556040000000
0!
0%
#556045000000
1!
1%
#556050000000
0!
0%
#556055000000
1!
1%
#556060000000
0!
0%
#556065000000
1!
1%
#556070000000
0!
0%
#556075000000
1!
1%
#556080000000
0!
0%
#556085000000
1!
1%
#556090000000
0!
0%
#556095000000
1!
1%
#556100000000
0!
0%
#556105000000
1!
1%
#556110000000
0!
0%
#556115000000
1!
1%
#556120000000
0!
0%
#556125000000
1!
1%
#556130000000
0!
0%
#556135000000
1!
1%
#556140000000
0!
0%
#556145000000
1!
1%
#556150000000
0!
0%
#556155000000
1!
1%
#556160000000
0!
0%
#556165000000
1!
1%
#556170000000
0!
0%
#556175000000
1!
1%
#556180000000
0!
0%
#556185000000
1!
1%
#556190000000
0!
0%
#556195000000
1!
1%
#556200000000
0!
0%
#556205000000
1!
1%
#556210000000
0!
0%
#556215000000
1!
1%
#556220000000
0!
0%
#556225000000
1!
1%
#556230000000
0!
0%
#556235000000
1!
1%
#556240000000
0!
0%
#556245000000
1!
1%
#556250000000
0!
0%
#556255000000
1!
1%
#556260000000
0!
0%
#556265000000
1!
1%
#556270000000
0!
0%
#556275000000
1!
1%
#556280000000
0!
0%
#556285000000
1!
1%
#556290000000
0!
0%
#556295000000
1!
1%
#556300000000
0!
0%
#556305000000
1!
1%
#556310000000
0!
0%
#556315000000
1!
1%
#556320000000
0!
0%
#556325000000
1!
1%
#556330000000
0!
0%
#556335000000
1!
1%
#556340000000
0!
0%
#556345000000
1!
1%
#556350000000
0!
0%
#556355000000
1!
1%
#556360000000
0!
0%
#556365000000
1!
1%
#556370000000
0!
0%
#556375000000
1!
1%
#556380000000
0!
0%
#556385000000
1!
1%
#556390000000
0!
0%
#556395000000
1!
1%
#556400000000
0!
0%
#556405000000
1!
1%
#556410000000
0!
0%
#556415000000
1!
1%
#556420000000
0!
0%
#556425000000
1!
1%
#556430000000
0!
0%
#556435000000
1!
1%
#556440000000
0!
0%
#556445000000
1!
1%
#556450000000
0!
0%
#556455000000
1!
1%
#556460000000
0!
0%
#556465000000
1!
1%
#556470000000
0!
0%
#556475000000
1!
1%
#556480000000
0!
0%
#556485000000
1!
1%
#556490000000
0!
0%
#556495000000
1!
1%
#556500000000
0!
0%
#556505000000
1!
1%
#556510000000
0!
0%
#556515000000
1!
1%
#556520000000
0!
0%
#556525000000
1!
1%
#556530000000
0!
0%
#556535000000
1!
1%
#556540000000
0!
0%
#556545000000
1!
1%
#556550000000
0!
0%
#556555000000
1!
1%
#556560000000
0!
0%
#556565000000
1!
1%
#556570000000
0!
0%
#556575000000
1!
1%
#556580000000
0!
0%
#556585000000
1!
1%
#556590000000
0!
0%
#556595000000
1!
1%
#556600000000
0!
0%
#556605000000
1!
1%
#556610000000
0!
0%
#556615000000
1!
1%
#556620000000
0!
0%
#556625000000
1!
1%
#556630000000
0!
0%
#556635000000
1!
1%
#556640000000
0!
0%
#556645000000
1!
1%
#556650000000
0!
0%
#556655000000
1!
1%
#556660000000
0!
0%
#556665000000
1!
1%
#556670000000
0!
0%
#556675000000
1!
1%
#556680000000
0!
0%
#556685000000
1!
1%
#556690000000
0!
0%
#556695000000
1!
1%
#556700000000
0!
0%
#556705000000
1!
1%
#556710000000
0!
0%
#556715000000
1!
1%
#556720000000
0!
0%
#556725000000
1!
1%
#556730000000
0!
0%
#556735000000
1!
1%
#556740000000
0!
0%
#556745000000
1!
1%
#556750000000
0!
0%
#556755000000
1!
1%
#556760000000
0!
0%
#556765000000
1!
1%
#556770000000
0!
0%
#556775000000
1!
1%
#556780000000
0!
0%
#556785000000
1!
1%
#556790000000
0!
0%
#556795000000
1!
1%
#556800000000
0!
0%
#556805000000
1!
1%
#556810000000
0!
0%
#556815000000
1!
1%
#556820000000
0!
0%
#556825000000
1!
1%
#556830000000
0!
0%
#556835000000
1!
1%
#556840000000
0!
0%
#556845000000
1!
1%
#556850000000
0!
0%
#556855000000
1!
1%
#556860000000
0!
0%
#556865000000
1!
1%
#556870000000
0!
0%
#556875000000
1!
1%
#556880000000
0!
0%
#556885000000
1!
1%
#556890000000
0!
0%
#556895000000
1!
1%
#556900000000
0!
0%
#556905000000
1!
1%
#556910000000
0!
0%
#556915000000
1!
1%
#556920000000
0!
0%
#556925000000
1!
1%
#556930000000
0!
0%
#556935000000
1!
1%
#556940000000
0!
0%
#556945000000
1!
1%
#556950000000
0!
0%
#556955000000
1!
1%
#556960000000
0!
0%
#556965000000
1!
1%
#556970000000
0!
0%
#556975000000
1!
1%
#556980000000
0!
0%
#556985000000
1!
1%
#556990000000
0!
0%
#556995000000
1!
1%
#557000000000
0!
0%
#557005000000
1!
1%
#557010000000
0!
0%
#557015000000
1!
1%
#557020000000
0!
0%
#557025000000
1!
1%
#557030000000
0!
0%
#557035000000
1!
1%
#557040000000
0!
0%
#557045000000
1!
1%
#557050000000
0!
0%
#557055000000
1!
1%
#557060000000
0!
0%
#557065000000
1!
1%
#557070000000
0!
0%
#557075000000
1!
1%
#557080000000
0!
0%
#557085000000
1!
1%
#557090000000
0!
0%
#557095000000
1!
1%
#557100000000
0!
0%
#557105000000
1!
1%
#557110000000
0!
0%
#557115000000
1!
1%
#557120000000
0!
0%
#557125000000
1!
1%
#557130000000
0!
0%
#557135000000
1!
1%
#557140000000
0!
0%
#557145000000
1!
1%
#557150000000
0!
0%
#557155000000
1!
1%
#557160000000
0!
0%
#557165000000
1!
1%
#557170000000
0!
0%
#557175000000
1!
1%
#557180000000
0!
0%
#557185000000
1!
1%
#557190000000
0!
0%
#557195000000
1!
1%
#557200000000
0!
0%
#557205000000
1!
1%
#557210000000
0!
0%
#557215000000
1!
1%
#557220000000
0!
0%
#557225000000
1!
1%
#557230000000
0!
0%
#557235000000
1!
1%
#557240000000
0!
0%
#557245000000
1!
1%
#557250000000
0!
0%
#557255000000
1!
1%
#557260000000
0!
0%
#557265000000
1!
1%
#557270000000
0!
0%
#557275000000
1!
1%
#557280000000
0!
0%
#557285000000
1!
1%
#557290000000
0!
0%
#557295000000
1!
1%
#557300000000
0!
0%
#557305000000
1!
1%
#557310000000
0!
0%
#557315000000
1!
1%
#557320000000
0!
0%
#557325000000
1!
1%
#557330000000
0!
0%
#557335000000
1!
1%
#557340000000
0!
0%
#557345000000
1!
1%
#557350000000
0!
0%
#557355000000
1!
1%
#557360000000
0!
0%
#557365000000
1!
1%
#557370000000
0!
0%
#557375000000
1!
1%
#557380000000
0!
0%
#557385000000
1!
1%
#557390000000
0!
0%
#557395000000
1!
1%
#557400000000
0!
0%
#557405000000
1!
1%
#557410000000
0!
0%
#557415000000
1!
1%
#557420000000
0!
0%
#557425000000
1!
1%
#557430000000
0!
0%
#557435000000
1!
1%
#557440000000
0!
0%
#557445000000
1!
1%
#557450000000
0!
0%
#557455000000
1!
1%
#557460000000
0!
0%
#557465000000
1!
1%
#557470000000
0!
0%
#557475000000
1!
1%
#557480000000
0!
0%
#557485000000
1!
1%
#557490000000
0!
0%
#557495000000
1!
1%
#557500000000
0!
0%
#557505000000
1!
1%
#557510000000
0!
0%
#557515000000
1!
1%
#557520000000
0!
0%
#557525000000
1!
1%
#557530000000
0!
0%
#557535000000
1!
1%
#557540000000
0!
0%
#557545000000
1!
1%
#557550000000
0!
0%
#557555000000
1!
1%
#557560000000
0!
0%
#557565000000
1!
1%
#557570000000
0!
0%
#557575000000
1!
1%
#557580000000
0!
0%
#557585000000
1!
1%
#557590000000
0!
0%
#557595000000
1!
1%
#557600000000
0!
0%
#557605000000
1!
1%
#557610000000
0!
0%
#557615000000
1!
1%
#557620000000
0!
0%
#557625000000
1!
1%
#557630000000
0!
0%
#557635000000
1!
1%
#557640000000
0!
0%
#557645000000
1!
1%
#557650000000
0!
0%
#557655000000
1!
1%
#557660000000
0!
0%
#557665000000
1!
1%
#557670000000
0!
0%
#557675000000
1!
1%
#557680000000
0!
0%
#557685000000
1!
1%
#557690000000
0!
0%
#557695000000
1!
1%
#557700000000
0!
0%
#557705000000
1!
1%
#557710000000
0!
0%
#557715000000
1!
1%
#557720000000
0!
0%
#557725000000
1!
1%
#557730000000
0!
0%
#557735000000
1!
1%
#557740000000
0!
0%
#557745000000
1!
1%
#557750000000
0!
0%
#557755000000
1!
1%
#557760000000
0!
0%
#557765000000
1!
1%
#557770000000
0!
0%
#557775000000
1!
1%
#557780000000
0!
0%
#557785000000
1!
1%
#557790000000
0!
0%
#557795000000
1!
1%
#557800000000
0!
0%
#557805000000
1!
1%
#557810000000
0!
0%
#557815000000
1!
1%
#557820000000
0!
0%
#557825000000
1!
1%
#557830000000
0!
0%
#557835000000
1!
1%
#557840000000
0!
0%
#557845000000
1!
1%
#557850000000
0!
0%
#557855000000
1!
1%
#557860000000
0!
0%
#557865000000
1!
1%
#557870000000
0!
0%
#557875000000
1!
1%
#557880000000
0!
0%
#557885000000
1!
1%
#557890000000
0!
0%
#557895000000
1!
1%
#557900000000
0!
0%
#557905000000
1!
1%
#557910000000
0!
0%
#557915000000
1!
1%
#557920000000
0!
0%
#557925000000
1!
1%
#557930000000
0!
0%
#557935000000
1!
1%
#557940000000
0!
0%
#557945000000
1!
1%
#557950000000
0!
0%
#557955000000
1!
1%
#557960000000
0!
0%
#557965000000
1!
1%
#557970000000
0!
0%
#557975000000
1!
1%
#557980000000
0!
0%
#557985000000
1!
1%
#557990000000
0!
0%
#557995000000
1!
1%
#558000000000
0!
0%
#558005000000
1!
1%
#558010000000
0!
0%
#558015000000
1!
1%
#558020000000
0!
0%
#558025000000
1!
1%
#558030000000
0!
0%
#558035000000
1!
1%
#558040000000
0!
0%
#558045000000
1!
1%
#558050000000
0!
0%
#558055000000
1!
1%
#558060000000
0!
0%
#558065000000
1!
1%
#558070000000
0!
0%
#558075000000
1!
1%
#558080000000
0!
0%
#558085000000
1!
1%
#558090000000
0!
0%
#558095000000
1!
1%
#558100000000
0!
0%
#558105000000
1!
1%
#558110000000
0!
0%
#558115000000
1!
1%
#558120000000
0!
0%
#558125000000
1!
1%
#558130000000
0!
0%
#558135000000
1!
1%
#558140000000
0!
0%
#558145000000
1!
1%
#558150000000
0!
0%
#558155000000
1!
1%
#558160000000
0!
0%
#558165000000
1!
1%
#558170000000
0!
0%
#558175000000
1!
1%
#558180000000
0!
0%
#558185000000
1!
1%
#558190000000
0!
0%
#558195000000
1!
1%
#558200000000
0!
0%
#558205000000
1!
1%
#558210000000
0!
0%
#558215000000
1!
1%
#558220000000
0!
0%
#558225000000
1!
1%
#558230000000
0!
0%
#558235000000
1!
1%
#558240000000
0!
0%
#558245000000
1!
1%
#558250000000
0!
0%
#558255000000
1!
1%
#558260000000
0!
0%
#558265000000
1!
1%
#558270000000
0!
0%
#558275000000
1!
1%
#558280000000
0!
0%
#558285000000
1!
1%
#558290000000
0!
0%
#558295000000
1!
1%
#558300000000
0!
0%
#558305000000
1!
1%
#558310000000
0!
0%
#558315000000
1!
1%
#558320000000
0!
0%
#558325000000
1!
1%
#558330000000
0!
0%
#558335000000
1!
1%
#558340000000
0!
0%
#558345000000
1!
1%
#558350000000
0!
0%
#558355000000
1!
1%
#558360000000
0!
0%
#558365000000
1!
1%
#558370000000
0!
0%
#558375000000
1!
1%
#558380000000
0!
0%
#558385000000
1!
1%
#558390000000
0!
0%
#558395000000
1!
1%
#558400000000
0!
0%
#558405000000
1!
1%
#558410000000
0!
0%
#558415000000
1!
1%
#558420000000
0!
0%
#558425000000
1!
1%
#558430000000
0!
0%
#558435000000
1!
1%
#558440000000
0!
0%
#558445000000
1!
1%
#558450000000
0!
0%
#558455000000
1!
1%
#558460000000
0!
0%
#558465000000
1!
1%
#558470000000
0!
0%
#558475000000
1!
1%
#558480000000
0!
0%
#558485000000
1!
1%
#558490000000
0!
0%
#558495000000
1!
1%
#558500000000
0!
0%
#558505000000
1!
1%
#558510000000
0!
0%
#558515000000
1!
1%
#558520000000
0!
0%
#558525000000
1!
1%
#558530000000
0!
0%
#558535000000
1!
1%
#558540000000
0!
0%
#558545000000
1!
1%
#558550000000
0!
0%
#558555000000
1!
1%
#558560000000
0!
0%
#558565000000
1!
1%
#558570000000
0!
0%
#558575000000
1!
1%
#558580000000
0!
0%
#558585000000
1!
1%
#558590000000
0!
0%
#558595000000
1!
1%
#558600000000
0!
0%
#558605000000
1!
1%
#558610000000
0!
0%
#558615000000
1!
1%
#558620000000
0!
0%
#558625000000
1!
1%
#558630000000
0!
0%
#558635000000
1!
1%
#558640000000
0!
0%
#558645000000
1!
1%
#558650000000
0!
0%
#558655000000
1!
1%
#558660000000
0!
0%
#558665000000
1!
1%
#558670000000
0!
0%
#558675000000
1!
1%
#558680000000
0!
0%
#558685000000
1!
1%
#558690000000
0!
0%
#558695000000
1!
1%
#558700000000
0!
0%
#558705000000
1!
1%
#558710000000
0!
0%
#558715000000
1!
1%
#558720000000
0!
0%
#558725000000
1!
1%
#558730000000
0!
0%
#558735000000
1!
1%
#558740000000
0!
0%
#558745000000
1!
1%
#558750000000
0!
0%
#558755000000
1!
1%
#558760000000
0!
0%
#558765000000
1!
1%
#558770000000
0!
0%
#558775000000
1!
1%
#558780000000
0!
0%
#558785000000
1!
1%
#558790000000
0!
0%
#558795000000
1!
1%
#558800000000
0!
0%
#558805000000
1!
1%
#558810000000
0!
0%
#558815000000
1!
1%
#558820000000
0!
0%
#558825000000
1!
1%
#558830000000
0!
0%
#558835000000
1!
1%
#558840000000
0!
0%
#558845000000
1!
1%
#558850000000
0!
0%
#558855000000
1!
1%
#558860000000
0!
0%
#558865000000
1!
1%
#558870000000
0!
0%
#558875000000
1!
1%
#558880000000
0!
0%
#558885000000
1!
1%
#558890000000
0!
0%
#558895000000
1!
1%
#558900000000
0!
0%
#558905000000
1!
1%
#558910000000
0!
0%
#558915000000
1!
1%
#558920000000
0!
0%
#558925000000
1!
1%
#558930000000
0!
0%
#558935000000
1!
1%
#558940000000
0!
0%
#558945000000
1!
1%
#558950000000
0!
0%
#558955000000
1!
1%
#558960000000
0!
0%
#558965000000
1!
1%
#558970000000
0!
0%
#558975000000
1!
1%
#558980000000
0!
0%
#558985000000
1!
1%
#558990000000
0!
0%
#558995000000
1!
1%
#559000000000
0!
0%
#559005000000
1!
1%
#559010000000
0!
0%
#559015000000
1!
1%
#559020000000
0!
0%
#559025000000
1!
1%
#559030000000
0!
0%
#559035000000
1!
1%
#559040000000
0!
0%
#559045000000
1!
1%
#559050000000
0!
0%
#559055000000
1!
1%
#559060000000
0!
0%
#559065000000
1!
1%
#559070000000
0!
0%
#559075000000
1!
1%
#559080000000
0!
0%
#559085000000
1!
1%
#559090000000
0!
0%
#559095000000
1!
1%
#559100000000
0!
0%
#559105000000
1!
1%
#559110000000
0!
0%
#559115000000
1!
1%
#559120000000
0!
0%
#559125000000
1!
1%
#559130000000
0!
0%
#559135000000
1!
1%
#559140000000
0!
0%
#559145000000
1!
1%
#559150000000
0!
0%
#559155000000
1!
1%
#559160000000
0!
0%
#559165000000
1!
1%
#559170000000
0!
0%
#559175000000
1!
1%
#559180000000
0!
0%
#559185000000
1!
1%
#559190000000
0!
0%
#559195000000
1!
1%
#559200000000
0!
0%
#559205000000
1!
1%
#559210000000
0!
0%
#559215000000
1!
1%
#559220000000
0!
0%
#559225000000
1!
1%
#559230000000
0!
0%
#559235000000
1!
1%
#559240000000
0!
0%
#559245000000
1!
1%
#559250000000
0!
0%
#559255000000
1!
1%
#559260000000
0!
0%
#559265000000
1!
1%
#559270000000
0!
0%
#559275000000
1!
1%
#559280000000
0!
0%
#559285000000
1!
1%
#559290000000
0!
0%
#559295000000
1!
1%
#559300000000
0!
0%
#559305000000
1!
1%
#559310000000
0!
0%
#559315000000
1!
1%
#559320000000
0!
0%
#559325000000
1!
1%
#559330000000
0!
0%
#559335000000
1!
1%
#559340000000
0!
0%
#559345000000
1!
1%
#559350000000
0!
0%
#559355000000
1!
1%
#559360000000
0!
0%
#559365000000
1!
1%
#559370000000
0!
0%
#559375000000
1!
1%
#559380000000
0!
0%
#559385000000
1!
1%
#559390000000
0!
0%
#559395000000
1!
1%
#559400000000
0!
0%
#559405000000
1!
1%
#559410000000
0!
0%
#559415000000
1!
1%
#559420000000
0!
0%
#559425000000
1!
1%
#559430000000
0!
0%
#559435000000
1!
1%
#559440000000
0!
0%
#559445000000
1!
1%
#559450000000
0!
0%
#559455000000
1!
1%
#559460000000
0!
0%
#559465000000
1!
1%
#559470000000
0!
0%
#559475000000
1!
1%
#559480000000
0!
0%
#559485000000
1!
1%
#559490000000
0!
0%
#559495000000
1!
1%
#559500000000
0!
0%
#559505000000
1!
1%
#559510000000
0!
0%
#559515000000
1!
1%
#559520000000
0!
0%
#559525000000
1!
1%
#559530000000
0!
0%
#559535000000
1!
1%
#559540000000
0!
0%
#559545000000
1!
1%
#559550000000
0!
0%
#559555000000
1!
1%
#559560000000
0!
0%
#559565000000
1!
1%
#559570000000
0!
0%
#559575000000
1!
1%
#559580000000
0!
0%
#559585000000
1!
1%
#559590000000
0!
0%
#559595000000
1!
1%
#559600000000
0!
0%
#559605000000
1!
1%
#559610000000
0!
0%
#559615000000
1!
1%
#559620000000
0!
0%
#559625000000
1!
1%
#559630000000
0!
0%
#559635000000
1!
1%
#559640000000
0!
0%
#559645000000
1!
1%
#559650000000
0!
0%
#559655000000
1!
1%
#559660000000
0!
0%
#559665000000
1!
1%
#559670000000
0!
0%
#559675000000
1!
1%
#559680000000
0!
0%
#559685000000
1!
1%
#559690000000
0!
0%
#559695000000
1!
1%
#559700000000
0!
0%
#559705000000
1!
1%
#559710000000
0!
0%
#559715000000
1!
1%
#559720000000
0!
0%
#559725000000
1!
1%
#559730000000
0!
0%
#559735000000
1!
1%
#559740000000
0!
0%
#559745000000
1!
1%
#559750000000
0!
0%
#559755000000
1!
1%
#559760000000
0!
0%
#559765000000
1!
1%
#559770000000
0!
0%
#559775000000
1!
1%
#559780000000
0!
0%
#559785000000
1!
1%
#559790000000
0!
0%
#559795000000
1!
1%
#559800000000
0!
0%
#559805000000
1!
1%
#559810000000
0!
0%
#559815000000
1!
1%
#559820000000
0!
0%
#559825000000
1!
1%
#559830000000
0!
0%
#559835000000
1!
1%
#559840000000
0!
0%
#559845000000
1!
1%
#559850000000
0!
0%
#559855000000
1!
1%
#559860000000
0!
0%
#559865000000
1!
1%
#559870000000
0!
0%
#559875000000
1!
1%
#559880000000
0!
0%
#559885000000
1!
1%
#559890000000
0!
0%
#559895000000
1!
1%
#559900000000
0!
0%
#559905000000
1!
1%
#559910000000
0!
0%
#559915000000
1!
1%
#559920000000
0!
0%
#559925000000
1!
1%
#559930000000
0!
0%
#559935000000
1!
1%
#559940000000
0!
0%
#559945000000
1!
1%
#559950000000
0!
0%
#559955000000
1!
1%
#559960000000
0!
0%
#559965000000
1!
1%
#559970000000
0!
0%
#559975000000
1!
1%
#559980000000
0!
0%
#559985000000
1!
1%
#559990000000
0!
0%
#559995000000
1!
1%
#560000000000
0!
0%
#560005000000
1!
1%
#560010000000
0!
0%
#560015000000
1!
1%
#560020000000
0!
0%
#560025000000
1!
1%
#560030000000
0!
0%
#560035000000
1!
1%
#560040000000
0!
0%
#560045000000
1!
1%
#560050000000
0!
0%
#560055000000
1!
1%
#560060000000
0!
0%
#560065000000
1!
1%
#560070000000
0!
0%
#560075000000
1!
1%
#560080000000
0!
0%
#560085000000
1!
1%
#560090000000
0!
0%
#560095000000
1!
1%
#560100000000
0!
0%
#560105000000
1!
1%
#560110000000
0!
0%
#560115000000
1!
1%
#560120000000
0!
0%
#560125000000
1!
1%
#560130000000
0!
0%
#560135000000
1!
1%
#560140000000
0!
0%
#560145000000
1!
1%
#560150000000
0!
0%
#560155000000
1!
1%
#560160000000
0!
0%
#560165000000
1!
1%
#560170000000
0!
0%
#560175000000
1!
1%
#560180000000
0!
0%
#560185000000
1!
1%
#560190000000
0!
0%
#560195000000
1!
1%
#560200000000
0!
0%
#560205000000
1!
1%
#560210000000
0!
0%
#560215000000
1!
1%
#560220000000
0!
0%
#560225000000
1!
1%
#560230000000
0!
0%
#560235000000
1!
1%
#560240000000
0!
0%
#560245000000
1!
1%
#560250000000
0!
0%
#560255000000
1!
1%
#560260000000
0!
0%
#560265000000
1!
1%
#560270000000
0!
0%
#560275000000
1!
1%
#560280000000
0!
0%
#560285000000
1!
1%
#560290000000
0!
0%
#560295000000
1!
1%
#560300000000
0!
0%
#560305000000
1!
1%
#560310000000
0!
0%
#560315000000
1!
1%
#560320000000
0!
0%
#560325000000
1!
1%
#560330000000
0!
0%
#560335000000
1!
1%
#560340000000
0!
0%
#560345000000
1!
1%
#560350000000
0!
0%
#560355000000
1!
1%
#560360000000
0!
0%
#560365000000
1!
1%
#560370000000
0!
0%
#560375000000
1!
1%
#560380000000
0!
0%
#560385000000
1!
1%
#560390000000
0!
0%
#560395000000
1!
1%
#560400000000
0!
0%
#560405000000
1!
1%
#560410000000
0!
0%
#560415000000
1!
1%
#560420000000
0!
0%
#560425000000
1!
1%
#560430000000
0!
0%
#560435000000
1!
1%
#560440000000
0!
0%
#560445000000
1!
1%
#560450000000
0!
0%
#560455000000
1!
1%
#560460000000
0!
0%
#560465000000
1!
1%
#560470000000
0!
0%
#560475000000
1!
1%
#560480000000
0!
0%
#560485000000
1!
1%
#560490000000
0!
0%
#560495000000
1!
1%
#560500000000
0!
0%
#560505000000
1!
1%
#560510000000
0!
0%
#560515000000
1!
1%
#560520000000
0!
0%
#560525000000
1!
1%
#560530000000
0!
0%
#560535000000
1!
1%
#560540000000
0!
0%
#560545000000
1!
1%
#560550000000
0!
0%
#560555000000
1!
1%
#560560000000
0!
0%
#560565000000
1!
1%
#560570000000
0!
0%
#560575000000
1!
1%
#560580000000
0!
0%
#560585000000
1!
1%
#560590000000
0!
0%
#560595000000
1!
1%
#560600000000
0!
0%
#560605000000
1!
1%
#560610000000
0!
0%
#560615000000
1!
1%
#560620000000
0!
0%
#560625000000
1!
1%
#560630000000
0!
0%
#560635000000
1!
1%
#560640000000
0!
0%
#560645000000
1!
1%
#560650000000
0!
0%
#560655000000
1!
1%
#560660000000
0!
0%
#560665000000
1!
1%
#560670000000
0!
0%
#560675000000
1!
1%
#560680000000
0!
0%
#560685000000
1!
1%
#560690000000
0!
0%
#560695000000
1!
1%
#560700000000
0!
0%
#560705000000
1!
1%
#560710000000
0!
0%
#560715000000
1!
1%
#560720000000
0!
0%
#560725000000
1!
1%
#560730000000
0!
0%
#560735000000
1!
1%
#560740000000
0!
0%
#560745000000
1!
1%
#560750000000
0!
0%
#560755000000
1!
1%
#560760000000
0!
0%
#560765000000
1!
1%
#560770000000
0!
0%
#560775000000
1!
1%
#560780000000
0!
0%
#560785000000
1!
1%
#560790000000
0!
0%
#560795000000
1!
1%
#560800000000
0!
0%
#560805000000
1!
1%
#560810000000
0!
0%
#560815000000
1!
1%
#560820000000
0!
0%
#560825000000
1!
1%
#560830000000
0!
0%
#560835000000
1!
1%
#560840000000
0!
0%
#560845000000
1!
1%
#560850000000
0!
0%
#560855000000
1!
1%
#560860000000
0!
0%
#560865000000
1!
1%
#560870000000
0!
0%
#560875000000
1!
1%
#560880000000
0!
0%
#560885000000
1!
1%
#560890000000
0!
0%
#560895000000
1!
1%
#560900000000
0!
0%
#560905000000
1!
1%
#560910000000
0!
0%
#560915000000
1!
1%
#560920000000
0!
0%
#560925000000
1!
1%
#560930000000
0!
0%
#560935000000
1!
1%
#560940000000
0!
0%
#560945000000
1!
1%
#560950000000
0!
0%
#560955000000
1!
1%
#560960000000
0!
0%
#560965000000
1!
1%
#560970000000
0!
0%
#560975000000
1!
1%
#560980000000
0!
0%
#560985000000
1!
1%
#560990000000
0!
0%
#560995000000
1!
1%
#561000000000
0!
0%
#561005000000
1!
1%
#561010000000
0!
0%
#561015000000
1!
1%
#561020000000
0!
0%
#561025000000
1!
1%
#561030000000
0!
0%
#561035000000
1!
1%
#561040000000
0!
0%
#561045000000
1!
1%
#561050000000
0!
0%
#561055000000
1!
1%
#561060000000
0!
0%
#561065000000
1!
1%
#561070000000
0!
0%
#561075000000
1!
1%
#561080000000
0!
0%
#561085000000
1!
1%
#561090000000
0!
0%
#561095000000
1!
1%
#561100000000
0!
0%
#561105000000
1!
1%
#561110000000
0!
0%
#561115000000
1!
1%
#561120000000
0!
0%
#561125000000
1!
1%
#561130000000
0!
0%
#561135000000
1!
1%
#561140000000
0!
0%
#561145000000
1!
1%
#561150000000
0!
0%
#561155000000
1!
1%
#561160000000
0!
0%
#561165000000
1!
1%
#561170000000
0!
0%
#561175000000
1!
1%
#561180000000
0!
0%
#561185000000
1!
1%
#561190000000
0!
0%
#561195000000
1!
1%
#561200000000
0!
0%
#561205000000
1!
1%
#561210000000
0!
0%
#561215000000
1!
1%
#561220000000
0!
0%
#561225000000
1!
1%
#561230000000
0!
0%
#561235000000
1!
1%
#561240000000
0!
0%
#561245000000
1!
1%
#561250000000
0!
0%
#561255000000
1!
1%
#561260000000
0!
0%
#561265000000
1!
1%
#561270000000
0!
0%
#561275000000
1!
1%
#561280000000
0!
0%
#561285000000
1!
1%
#561290000000
0!
0%
#561295000000
1!
1%
#561300000000
0!
0%
#561305000000
1!
1%
#561310000000
0!
0%
#561315000000
1!
1%
#561320000000
0!
0%
#561325000000
1!
1%
#561330000000
0!
0%
#561335000000
1!
1%
#561340000000
0!
0%
#561345000000
1!
1%
#561350000000
0!
0%
#561355000000
1!
1%
#561360000000
0!
0%
#561365000000
1!
1%
#561370000000
0!
0%
#561375000000
1!
1%
#561380000000
0!
0%
#561385000000
1!
1%
#561390000000
0!
0%
#561395000000
1!
1%
#561400000000
0!
0%
#561405000000
1!
1%
#561410000000
0!
0%
#561415000000
1!
1%
#561420000000
0!
0%
#561425000000
1!
1%
#561430000000
0!
0%
#561435000000
1!
1%
#561440000000
0!
0%
#561445000000
1!
1%
#561450000000
0!
0%
#561455000000
1!
1%
#561460000000
0!
0%
#561465000000
1!
1%
#561470000000
0!
0%
#561475000000
1!
1%
#561480000000
0!
0%
#561485000000
1!
1%
#561490000000
0!
0%
#561495000000
1!
1%
#561500000000
0!
0%
#561505000000
1!
1%
#561510000000
0!
0%
#561515000000
1!
1%
#561520000000
0!
0%
#561525000000
1!
1%
#561530000000
0!
0%
#561535000000
1!
1%
#561540000000
0!
0%
#561545000000
1!
1%
#561550000000
0!
0%
#561555000000
1!
1%
#561560000000
0!
0%
#561565000000
1!
1%
#561570000000
0!
0%
#561575000000
1!
1%
#561580000000
0!
0%
#561585000000
1!
1%
#561590000000
0!
0%
#561595000000
1!
1%
#561600000000
0!
0%
#561605000000
1!
1%
#561610000000
0!
0%
#561615000000
1!
1%
#561620000000
0!
0%
#561625000000
1!
1%
#561630000000
0!
0%
#561635000000
1!
1%
#561640000000
0!
0%
#561645000000
1!
1%
#561650000000
0!
0%
#561655000000
1!
1%
#561660000000
0!
0%
#561665000000
1!
1%
#561670000000
0!
0%
#561675000000
1!
1%
#561680000000
0!
0%
#561685000000
1!
1%
#561690000000
0!
0%
#561695000000
1!
1%
#561700000000
0!
0%
#561705000000
1!
1%
#561710000000
0!
0%
#561715000000
1!
1%
#561720000000
0!
0%
#561725000000
1!
1%
#561730000000
0!
0%
#561735000000
1!
1%
#561740000000
0!
0%
#561745000000
1!
1%
#561750000000
0!
0%
#561755000000
1!
1%
#561760000000
0!
0%
#561765000000
1!
1%
#561770000000
0!
0%
#561775000000
1!
1%
#561780000000
0!
0%
#561785000000
1!
1%
#561790000000
0!
0%
#561795000000
1!
1%
#561800000000
0!
0%
#561805000000
1!
1%
#561810000000
0!
0%
#561815000000
1!
1%
#561820000000
0!
0%
#561825000000
1!
1%
#561830000000
0!
0%
#561835000000
1!
1%
#561840000000
0!
0%
#561845000000
1!
1%
#561850000000
0!
0%
#561855000000
1!
1%
#561860000000
0!
0%
#561865000000
1!
1%
#561870000000
0!
0%
#561875000000
1!
1%
#561880000000
0!
0%
#561885000000
1!
1%
#561890000000
0!
0%
#561895000000
1!
1%
#561900000000
0!
0%
#561905000000
1!
1%
#561910000000
0!
0%
#561915000000
1!
1%
#561920000000
0!
0%
#561925000000
1!
1%
#561930000000
0!
0%
#561935000000
1!
1%
#561940000000
0!
0%
#561945000000
1!
1%
#561950000000
0!
0%
#561955000000
1!
1%
#561960000000
0!
0%
#561965000000
1!
1%
#561970000000
0!
0%
#561975000000
1!
1%
#561980000000
0!
0%
#561985000000
1!
1%
#561990000000
0!
0%
#561995000000
1!
1%
#562000000000
0!
0%
#562005000000
1!
1%
#562010000000
0!
0%
#562015000000
1!
1%
#562020000000
0!
0%
#562025000000
1!
1%
#562030000000
0!
0%
#562035000000
1!
1%
#562040000000
0!
0%
#562045000000
1!
1%
#562050000000
0!
0%
#562055000000
1!
1%
#562060000000
0!
0%
#562065000000
1!
1%
#562070000000
0!
0%
#562075000000
1!
1%
#562080000000
0!
0%
#562085000000
1!
1%
#562090000000
0!
0%
#562095000000
1!
1%
#562100000000
0!
0%
#562105000000
1!
1%
#562110000000
0!
0%
#562115000000
1!
1%
#562120000000
0!
0%
#562125000000
1!
1%
#562130000000
0!
0%
#562135000000
1!
1%
#562140000000
0!
0%
#562145000000
1!
1%
#562150000000
0!
0%
#562155000000
1!
1%
#562160000000
0!
0%
#562165000000
1!
1%
#562170000000
0!
0%
#562175000000
1!
1%
#562180000000
0!
0%
#562185000000
1!
1%
#562190000000
0!
0%
#562195000000
1!
1%
#562200000000
0!
0%
#562205000000
1!
1%
#562210000000
0!
0%
#562215000000
1!
1%
#562220000000
0!
0%
#562225000000
1!
1%
#562230000000
0!
0%
#562235000000
1!
1%
#562240000000
0!
0%
#562245000000
1!
1%
#562250000000
0!
0%
#562255000000
1!
1%
#562260000000
0!
0%
#562265000000
1!
1%
#562270000000
0!
0%
#562275000000
1!
1%
#562280000000
0!
0%
#562285000000
1!
1%
#562290000000
0!
0%
#562295000000
1!
1%
#562300000000
0!
0%
#562305000000
1!
1%
#562310000000
0!
0%
#562315000000
1!
1%
#562320000000
0!
0%
#562325000000
1!
1%
#562330000000
0!
0%
#562335000000
1!
1%
#562340000000
0!
0%
#562345000000
1!
1%
#562350000000
0!
0%
#562355000000
1!
1%
#562360000000
0!
0%
#562365000000
1!
1%
#562370000000
0!
0%
#562375000000
1!
1%
#562380000000
0!
0%
#562385000000
1!
1%
#562390000000
0!
0%
#562395000000
1!
1%
#562400000000
0!
0%
#562405000000
1!
1%
#562410000000
0!
0%
#562415000000
1!
1%
#562420000000
0!
0%
#562425000000
1!
1%
#562430000000
0!
0%
#562435000000
1!
1%
#562440000000
0!
0%
#562445000000
1!
1%
#562450000000
0!
0%
#562455000000
1!
1%
#562460000000
0!
0%
#562465000000
1!
1%
#562470000000
0!
0%
#562475000000
1!
1%
#562480000000
0!
0%
#562485000000
1!
1%
#562490000000
0!
0%
#562495000000
1!
1%
#562500000000
0!
0%
#562505000000
1!
1%
#562510000000
0!
0%
#562515000000
1!
1%
#562520000000
0!
0%
#562525000000
1!
1%
#562530000000
0!
0%
#562535000000
1!
1%
#562540000000
0!
0%
#562545000000
1!
1%
#562550000000
0!
0%
#562555000000
1!
1%
#562560000000
0!
0%
#562565000000
1!
1%
#562570000000
0!
0%
#562575000000
1!
1%
#562580000000
0!
0%
#562585000000
1!
1%
#562590000000
0!
0%
#562595000000
1!
1%
#562600000000
0!
0%
#562605000000
1!
1%
#562610000000
0!
0%
#562615000000
1!
1%
#562620000000
0!
0%
#562625000000
1!
1%
#562630000000
0!
0%
#562635000000
1!
1%
#562640000000
0!
0%
#562645000000
1!
1%
#562650000000
0!
0%
#562655000000
1!
1%
#562660000000
0!
0%
#562665000000
1!
1%
#562670000000
0!
0%
#562675000000
1!
1%
#562680000000
0!
0%
#562685000000
1!
1%
#562690000000
0!
0%
#562695000000
1!
1%
#562700000000
0!
0%
#562705000000
1!
1%
#562710000000
0!
0%
#562715000000
1!
1%
#562720000000
0!
0%
#562725000000
1!
1%
#562730000000
0!
0%
#562735000000
1!
1%
#562740000000
0!
0%
#562745000000
1!
1%
#562750000000
0!
0%
#562755000000
1!
1%
#562760000000
0!
0%
#562765000000
1!
1%
#562770000000
0!
0%
#562775000000
1!
1%
#562780000000
0!
0%
#562785000000
1!
1%
#562790000000
0!
0%
#562795000000
1!
1%
#562800000000
0!
0%
#562805000000
1!
1%
#562810000000
0!
0%
#562815000000
1!
1%
#562820000000
0!
0%
#562825000000
1!
1%
#562830000000
0!
0%
#562835000000
1!
1%
#562840000000
0!
0%
#562845000000
1!
1%
#562850000000
0!
0%
#562855000000
1!
1%
#562860000000
0!
0%
#562865000000
1!
1%
#562870000000
0!
0%
#562875000000
1!
1%
#562880000000
0!
0%
#562885000000
1!
1%
#562890000000
0!
0%
#562895000000
1!
1%
#562900000000
0!
0%
#562905000000
1!
1%
#562910000000
0!
0%
#562915000000
1!
1%
#562920000000
0!
0%
#562925000000
1!
1%
#562930000000
0!
0%
#562935000000
1!
1%
#562940000000
0!
0%
#562945000000
1!
1%
#562950000000
0!
0%
#562955000000
1!
1%
#562960000000
0!
0%
#562965000000
1!
1%
#562970000000
0!
0%
#562975000000
1!
1%
#562980000000
0!
0%
#562985000000
1!
1%
#562990000000
0!
0%
#562995000000
1!
1%
#563000000000
0!
0%
#563005000000
1!
1%
#563010000000
0!
0%
#563015000000
1!
1%
#563020000000
0!
0%
#563025000000
1!
1%
#563030000000
0!
0%
#563035000000
1!
1%
#563040000000
0!
0%
#563045000000
1!
1%
#563050000000
0!
0%
#563055000000
1!
1%
#563060000000
0!
0%
#563065000000
1!
1%
#563070000000
0!
0%
#563075000000
1!
1%
#563080000000
0!
0%
#563085000000
1!
1%
#563090000000
0!
0%
#563095000000
1!
1%
#563100000000
0!
0%
#563105000000
1!
1%
#563110000000
0!
0%
#563115000000
1!
1%
#563120000000
0!
0%
#563125000000
1!
1%
#563130000000
0!
0%
#563135000000
1!
1%
#563140000000
0!
0%
#563145000000
1!
1%
#563150000000
0!
0%
#563155000000
1!
1%
#563160000000
0!
0%
#563165000000
1!
1%
#563170000000
0!
0%
#563175000000
1!
1%
#563180000000
0!
0%
#563185000000
1!
1%
#563190000000
0!
0%
#563195000000
1!
1%
#563200000000
0!
0%
#563205000000
1!
1%
#563210000000
0!
0%
#563215000000
1!
1%
#563220000000
0!
0%
#563225000000
1!
1%
#563230000000
0!
0%
#563235000000
1!
1%
#563240000000
0!
0%
#563245000000
1!
1%
#563250000000
0!
0%
#563255000000
1!
1%
#563260000000
0!
0%
#563265000000
1!
1%
#563270000000
0!
0%
#563275000000
1!
1%
#563280000000
0!
0%
#563285000000
1!
1%
#563290000000
0!
0%
#563295000000
1!
1%
#563300000000
0!
0%
#563305000000
1!
1%
#563310000000
0!
0%
#563315000000
1!
1%
#563320000000
0!
0%
#563325000000
1!
1%
#563330000000
0!
0%
#563335000000
1!
1%
#563340000000
0!
0%
#563345000000
1!
1%
#563350000000
0!
0%
#563355000000
1!
1%
#563360000000
0!
0%
#563365000000
1!
1%
#563370000000
0!
0%
#563375000000
1!
1%
#563380000000
0!
0%
#563385000000
1!
1%
#563390000000
0!
0%
#563395000000
1!
1%
#563400000000
0!
0%
#563405000000
1!
1%
#563410000000
0!
0%
#563415000000
1!
1%
#563420000000
0!
0%
#563425000000
1!
1%
#563430000000
0!
0%
#563435000000
1!
1%
#563440000000
0!
0%
#563445000000
1!
1%
#563450000000
0!
0%
#563455000000
1!
1%
#563460000000
0!
0%
#563465000000
1!
1%
#563470000000
0!
0%
#563475000000
1!
1%
#563480000000
0!
0%
#563485000000
1!
1%
#563490000000
0!
0%
#563495000000
1!
1%
#563500000000
0!
0%
#563505000000
1!
1%
#563510000000
0!
0%
#563515000000
1!
1%
#563520000000
0!
0%
#563525000000
1!
1%
#563530000000
0!
0%
#563535000000
1!
1%
#563540000000
0!
0%
#563545000000
1!
1%
#563550000000
0!
0%
#563555000000
1!
1%
#563560000000
0!
0%
#563565000000
1!
1%
#563570000000
0!
0%
#563575000000
1!
1%
#563580000000
0!
0%
#563585000000
1!
1%
#563590000000
0!
0%
#563595000000
1!
1%
#563600000000
0!
0%
#563605000000
1!
1%
#563610000000
0!
0%
#563615000000
1!
1%
#563620000000
0!
0%
#563625000000
1!
1%
#563630000000
0!
0%
#563635000000
1!
1%
#563640000000
0!
0%
#563645000000
1!
1%
#563650000000
0!
0%
#563655000000
1!
1%
#563660000000
0!
0%
#563665000000
1!
1%
#563670000000
0!
0%
#563675000000
1!
1%
#563680000000
0!
0%
#563685000000
1!
1%
#563690000000
0!
0%
#563695000000
1!
1%
#563700000000
0!
0%
#563705000000
1!
1%
#563710000000
0!
0%
#563715000000
1!
1%
#563720000000
0!
0%
#563725000000
1!
1%
#563730000000
0!
0%
#563735000000
1!
1%
#563740000000
0!
0%
#563745000000
1!
1%
#563750000000
0!
0%
#563755000000
1!
1%
#563760000000
0!
0%
#563765000000
1!
1%
#563770000000
0!
0%
#563775000000
1!
1%
#563780000000
0!
0%
#563785000000
1!
1%
#563790000000
0!
0%
#563795000000
1!
1%
#563800000000
0!
0%
#563805000000
1!
1%
#563810000000
0!
0%
#563815000000
1!
1%
#563820000000
0!
0%
#563825000000
1!
1%
#563830000000
0!
0%
#563835000000
1!
1%
#563840000000
0!
0%
#563845000000
1!
1%
#563850000000
0!
0%
#563855000000
1!
1%
#563860000000
0!
0%
#563865000000
1!
1%
#563870000000
0!
0%
#563875000000
1!
1%
#563880000000
0!
0%
#563885000000
1!
1%
#563890000000
0!
0%
#563895000000
1!
1%
#563900000000
0!
0%
#563905000000
1!
1%
#563910000000
0!
0%
#563915000000
1!
1%
#563920000000
0!
0%
#563925000000
1!
1%
#563930000000
0!
0%
#563935000000
1!
1%
#563940000000
0!
0%
#563945000000
1!
1%
#563950000000
0!
0%
#563955000000
1!
1%
#563960000000
0!
0%
#563965000000
1!
1%
#563970000000
0!
0%
#563975000000
1!
1%
#563980000000
0!
0%
#563985000000
1!
1%
#563990000000
0!
0%
#563995000000
1!
1%
#564000000000
0!
0%
#564005000000
1!
1%
#564010000000
0!
0%
#564015000000
1!
1%
#564020000000
0!
0%
#564025000000
1!
1%
#564030000000
0!
0%
#564035000000
1!
1%
#564040000000
0!
0%
#564045000000
1!
1%
#564050000000
0!
0%
#564055000000
1!
1%
#564060000000
0!
0%
#564065000000
1!
1%
#564070000000
0!
0%
#564075000000
1!
1%
#564080000000
0!
0%
#564085000000
1!
1%
#564090000000
0!
0%
#564095000000
1!
1%
#564100000000
0!
0%
#564105000000
1!
1%
#564110000000
0!
0%
#564115000000
1!
1%
#564120000000
0!
0%
#564125000000
1!
1%
#564130000000
0!
0%
#564135000000
1!
1%
#564140000000
0!
0%
#564145000000
1!
1%
#564150000000
0!
0%
#564155000000
1!
1%
#564160000000
0!
0%
#564165000000
1!
1%
#564170000000
0!
0%
#564175000000
1!
1%
#564180000000
0!
0%
#564185000000
1!
1%
#564190000000
0!
0%
#564195000000
1!
1%
#564200000000
0!
0%
#564205000000
1!
1%
#564210000000
0!
0%
#564215000000
1!
1%
#564220000000
0!
0%
#564225000000
1!
1%
#564230000000
0!
0%
#564235000000
1!
1%
#564240000000
0!
0%
#564245000000
1!
1%
#564250000000
0!
0%
#564255000000
1!
1%
#564260000000
0!
0%
#564265000000
1!
1%
#564270000000
0!
0%
#564275000000
1!
1%
#564280000000
0!
0%
#564285000000
1!
1%
#564290000000
0!
0%
#564295000000
1!
1%
#564300000000
0!
0%
#564305000000
1!
1%
#564310000000
0!
0%
#564315000000
1!
1%
#564320000000
0!
0%
#564325000000
1!
1%
#564330000000
0!
0%
#564335000000
1!
1%
#564340000000
0!
0%
#564345000000
1!
1%
#564350000000
0!
0%
#564355000000
1!
1%
#564360000000
0!
0%
#564365000000
1!
1%
#564370000000
0!
0%
#564375000000
1!
1%
#564380000000
0!
0%
#564385000000
1!
1%
#564390000000
0!
0%
#564395000000
1!
1%
#564400000000
0!
0%
#564405000000
1!
1%
#564410000000
0!
0%
#564415000000
1!
1%
#564420000000
0!
0%
#564425000000
1!
1%
#564430000000
0!
0%
#564435000000
1!
1%
#564440000000
0!
0%
#564445000000
1!
1%
#564450000000
0!
0%
#564455000000
1!
1%
#564460000000
0!
0%
#564465000000
1!
1%
#564470000000
0!
0%
#564475000000
1!
1%
#564480000000
0!
0%
#564485000000
1!
1%
#564490000000
0!
0%
#564495000000
1!
1%
#564500000000
0!
0%
#564505000000
1!
1%
#564510000000
0!
0%
#564515000000
1!
1%
#564520000000
0!
0%
#564525000000
1!
1%
#564530000000
0!
0%
#564535000000
1!
1%
#564540000000
0!
0%
#564545000000
1!
1%
#564550000000
0!
0%
#564555000000
1!
1%
#564560000000
0!
0%
#564565000000
1!
1%
#564570000000
0!
0%
#564575000000
1!
1%
#564580000000
0!
0%
#564585000000
1!
1%
#564590000000
0!
0%
#564595000000
1!
1%
#564600000000
0!
0%
#564605000000
1!
1%
#564610000000
0!
0%
#564615000000
1!
1%
#564620000000
0!
0%
#564625000000
1!
1%
#564630000000
0!
0%
#564635000000
1!
1%
#564640000000
0!
0%
#564645000000
1!
1%
#564650000000
0!
0%
#564655000000
1!
1%
#564660000000
0!
0%
#564665000000
1!
1%
#564670000000
0!
0%
#564675000000
1!
1%
#564680000000
0!
0%
#564685000000
1!
1%
#564690000000
0!
0%
#564695000000
1!
1%
#564700000000
0!
0%
#564705000000
1!
1%
#564710000000
0!
0%
#564715000000
1!
1%
#564720000000
0!
0%
#564725000000
1!
1%
#564730000000
0!
0%
#564735000000
1!
1%
#564740000000
0!
0%
#564745000000
1!
1%
#564750000000
0!
0%
#564755000000
1!
1%
#564760000000
0!
0%
#564765000000
1!
1%
#564770000000
0!
0%
#564775000000
1!
1%
#564780000000
0!
0%
#564785000000
1!
1%
#564790000000
0!
0%
#564795000000
1!
1%
#564800000000
0!
0%
#564805000000
1!
1%
#564810000000
0!
0%
#564815000000
1!
1%
#564820000000
0!
0%
#564825000000
1!
1%
#564830000000
0!
0%
#564835000000
1!
1%
#564840000000
0!
0%
#564845000000
1!
1%
#564850000000
0!
0%
#564855000000
1!
1%
#564860000000
0!
0%
#564865000000
1!
1%
#564870000000
0!
0%
#564875000000
1!
1%
#564880000000
0!
0%
#564885000000
1!
1%
#564890000000
0!
0%
#564895000000
1!
1%
#564900000000
0!
0%
#564905000000
1!
1%
#564910000000
0!
0%
#564915000000
1!
1%
#564920000000
0!
0%
#564925000000
1!
1%
#564930000000
0!
0%
#564935000000
1!
1%
#564940000000
0!
0%
#564945000000
1!
1%
#564950000000
0!
0%
#564955000000
1!
1%
#564960000000
0!
0%
#564965000000
1!
1%
#564970000000
0!
0%
#564975000000
1!
1%
#564980000000
0!
0%
#564985000000
1!
1%
#564990000000
0!
0%
#564995000000
1!
1%
#565000000000
0!
0%
#565005000000
1!
1%
#565010000000
0!
0%
#565015000000
1!
1%
#565020000000
0!
0%
#565025000000
1!
1%
#565030000000
0!
0%
#565035000000
1!
1%
#565040000000
0!
0%
#565045000000
1!
1%
#565050000000
0!
0%
#565055000000
1!
1%
#565060000000
0!
0%
#565065000000
1!
1%
#565070000000
0!
0%
#565075000000
1!
1%
#565080000000
0!
0%
#565085000000
1!
1%
#565090000000
0!
0%
#565095000000
1!
1%
#565100000000
0!
0%
#565105000000
1!
1%
#565110000000
0!
0%
#565115000000
1!
1%
#565120000000
0!
0%
#565125000000
1!
1%
#565130000000
0!
0%
#565135000000
1!
1%
#565140000000
0!
0%
#565145000000
1!
1%
#565150000000
0!
0%
#565155000000
1!
1%
#565160000000
0!
0%
#565165000000
1!
1%
#565170000000
0!
0%
#565175000000
1!
1%
#565180000000
0!
0%
#565185000000
1!
1%
#565190000000
0!
0%
#565195000000
1!
1%
#565200000000
0!
0%
#565205000000
1!
1%
#565210000000
0!
0%
#565215000000
1!
1%
#565220000000
0!
0%
#565225000000
1!
1%
#565230000000
0!
0%
#565235000000
1!
1%
#565240000000
0!
0%
#565245000000
1!
1%
#565250000000
0!
0%
#565255000000
1!
1%
#565260000000
0!
0%
#565265000000
1!
1%
#565270000000
0!
0%
#565275000000
1!
1%
#565280000000
0!
0%
#565285000000
1!
1%
#565290000000
0!
0%
#565295000000
1!
1%
#565300000000
0!
0%
#565305000000
1!
1%
#565310000000
0!
0%
#565315000000
1!
1%
#565320000000
0!
0%
#565325000000
1!
1%
#565330000000
0!
0%
#565335000000
1!
1%
#565340000000
0!
0%
#565345000000
1!
1%
#565350000000
0!
0%
#565355000000
1!
1%
#565360000000
0!
0%
#565365000000
1!
1%
#565370000000
0!
0%
#565375000000
1!
1%
#565380000000
0!
0%
#565385000000
1!
1%
#565390000000
0!
0%
#565395000000
1!
1%
#565400000000
0!
0%
#565405000000
1!
1%
#565410000000
0!
0%
#565415000000
1!
1%
#565420000000
0!
0%
#565425000000
1!
1%
#565430000000
0!
0%
#565435000000
1!
1%
#565440000000
0!
0%
#565445000000
1!
1%
#565450000000
0!
0%
#565455000000
1!
1%
#565460000000
0!
0%
#565465000000
1!
1%
#565470000000
0!
0%
#565475000000
1!
1%
#565480000000
0!
0%
#565485000000
1!
1%
#565490000000
0!
0%
#565495000000
1!
1%
#565500000000
0!
0%
#565505000000
1!
1%
#565510000000
0!
0%
#565515000000
1!
1%
#565520000000
0!
0%
#565525000000
1!
1%
#565530000000
0!
0%
#565535000000
1!
1%
#565540000000
0!
0%
#565545000000
1!
1%
#565550000000
0!
0%
#565555000000
1!
1%
#565560000000
0!
0%
#565565000000
1!
1%
#565570000000
0!
0%
#565575000000
1!
1%
#565580000000
0!
0%
#565585000000
1!
1%
#565590000000
0!
0%
#565595000000
1!
1%
#565600000000
0!
0%
#565605000000
1!
1%
#565610000000
0!
0%
#565615000000
1!
1%
#565620000000
0!
0%
#565625000000
1!
1%
#565630000000
0!
0%
#565635000000
1!
1%
#565640000000
0!
0%
#565645000000
1!
1%
#565650000000
0!
0%
#565655000000
1!
1%
#565660000000
0!
0%
#565665000000
1!
1%
#565670000000
0!
0%
#565675000000
1!
1%
#565680000000
0!
0%
#565685000000
1!
1%
#565690000000
0!
0%
#565695000000
1!
1%
#565700000000
0!
0%
#565705000000
1!
1%
#565710000000
0!
0%
#565715000000
1!
1%
#565720000000
0!
0%
#565725000000
1!
1%
#565730000000
0!
0%
#565735000000
1!
1%
#565740000000
0!
0%
#565745000000
1!
1%
#565750000000
0!
0%
#565755000000
1!
1%
#565760000000
0!
0%
#565765000000
1!
1%
#565770000000
0!
0%
#565775000000
1!
1%
#565780000000
0!
0%
#565785000000
1!
1%
#565790000000
0!
0%
#565795000000
1!
1%
#565800000000
0!
0%
#565805000000
1!
1%
#565810000000
0!
0%
#565815000000
1!
1%
#565820000000
0!
0%
#565825000000
1!
1%
#565830000000
0!
0%
#565835000000
1!
1%
#565840000000
0!
0%
#565845000000
1!
1%
#565850000000
0!
0%
#565855000000
1!
1%
#565860000000
0!
0%
#565865000000
1!
1%
#565870000000
0!
0%
#565875000000
1!
1%
#565880000000
0!
0%
#565885000000
1!
1%
#565890000000
0!
0%
#565895000000
1!
1%
#565900000000
0!
0%
#565905000000
1!
1%
#565910000000
0!
0%
#565915000000
1!
1%
#565920000000
0!
0%
#565925000000
1!
1%
#565930000000
0!
0%
#565935000000
1!
1%
#565940000000
0!
0%
#565945000000
1!
1%
#565950000000
0!
0%
#565955000000
1!
1%
#565960000000
0!
0%
#565965000000
1!
1%
#565970000000
0!
0%
#565975000000
1!
1%
#565980000000
0!
0%
#565985000000
1!
1%
#565990000000
0!
0%
#565995000000
1!
1%
#566000000000
0!
0%
#566005000000
1!
1%
#566010000000
0!
0%
#566015000000
1!
1%
#566020000000
0!
0%
#566025000000
1!
1%
#566030000000
0!
0%
#566035000000
1!
1%
#566040000000
0!
0%
#566045000000
1!
1%
#566050000000
0!
0%
#566055000000
1!
1%
#566060000000
0!
0%
#566065000000
1!
1%
#566070000000
0!
0%
#566075000000
1!
1%
#566080000000
0!
0%
#566085000000
1!
1%
#566090000000
0!
0%
#566095000000
1!
1%
#566100000000
0!
0%
#566105000000
1!
1%
#566110000000
0!
0%
#566115000000
1!
1%
#566120000000
0!
0%
#566125000000
1!
1%
#566130000000
0!
0%
#566135000000
1!
1%
#566140000000
0!
0%
#566145000000
1!
1%
#566150000000
0!
0%
#566155000000
1!
1%
#566160000000
0!
0%
#566165000000
1!
1%
#566170000000
0!
0%
#566175000000
1!
1%
#566180000000
0!
0%
#566185000000
1!
1%
#566190000000
0!
0%
#566195000000
1!
1%
#566200000000
0!
0%
#566205000000
1!
1%
#566210000000
0!
0%
#566215000000
1!
1%
#566220000000
0!
0%
#566225000000
1!
1%
#566230000000
0!
0%
#566235000000
1!
1%
#566240000000
0!
0%
#566245000000
1!
1%
#566250000000
0!
0%
#566255000000
1!
1%
#566260000000
0!
0%
#566265000000
1!
1%
#566270000000
0!
0%
#566275000000
1!
1%
#566280000000
0!
0%
#566285000000
1!
1%
#566290000000
0!
0%
#566295000000
1!
1%
#566300000000
0!
0%
#566305000000
1!
1%
#566310000000
0!
0%
#566315000000
1!
1%
#566320000000
0!
0%
#566325000000
1!
1%
#566330000000
0!
0%
#566335000000
1!
1%
#566340000000
0!
0%
#566345000000
1!
1%
#566350000000
0!
0%
#566355000000
1!
1%
#566360000000
0!
0%
#566365000000
1!
1%
#566370000000
0!
0%
#566375000000
1!
1%
#566380000000
0!
0%
#566385000000
1!
1%
#566390000000
0!
0%
#566395000000
1!
1%
#566400000000
0!
0%
#566405000000
1!
1%
#566410000000
0!
0%
#566415000000
1!
1%
#566420000000
0!
0%
#566425000000
1!
1%
#566430000000
0!
0%
#566435000000
1!
1%
#566440000000
0!
0%
#566445000000
1!
1%
#566450000000
0!
0%
#566455000000
1!
1%
#566460000000
0!
0%
#566465000000
1!
1%
#566470000000
0!
0%
#566475000000
1!
1%
#566480000000
0!
0%
#566485000000
1!
1%
#566490000000
0!
0%
#566495000000
1!
1%
#566500000000
0!
0%
#566505000000
1!
1%
#566510000000
0!
0%
#566515000000
1!
1%
#566520000000
0!
0%
#566525000000
1!
1%
#566530000000
0!
0%
#566535000000
1!
1%
#566540000000
0!
0%
#566545000000
1!
1%
#566550000000
0!
0%
#566555000000
1!
1%
#566560000000
0!
0%
#566565000000
1!
1%
#566570000000
0!
0%
#566575000000
1!
1%
#566580000000
0!
0%
#566585000000
1!
1%
#566590000000
0!
0%
#566595000000
1!
1%
#566600000000
0!
0%
#566605000000
1!
1%
#566610000000
0!
0%
#566615000000
1!
1%
#566620000000
0!
0%
#566625000000
1!
1%
#566630000000
0!
0%
#566635000000
1!
1%
#566640000000
0!
0%
#566645000000
1!
1%
#566650000000
0!
0%
#566655000000
1!
1%
#566660000000
0!
0%
#566665000000
1!
1%
#566670000000
0!
0%
#566675000000
1!
1%
#566680000000
0!
0%
#566685000000
1!
1%
#566690000000
0!
0%
#566695000000
1!
1%
#566700000000
0!
0%
#566705000000
1!
1%
#566710000000
0!
0%
#566715000000
1!
1%
#566720000000
0!
0%
#566725000000
1!
1%
#566730000000
0!
0%
#566735000000
1!
1%
#566740000000
0!
0%
#566745000000
1!
1%
#566750000000
0!
0%
#566755000000
1!
1%
#566760000000
0!
0%
#566765000000
1!
1%
#566770000000
0!
0%
#566775000000
1!
1%
#566780000000
0!
0%
#566785000000
1!
1%
#566790000000
0!
0%
#566795000000
1!
1%
#566800000000
0!
0%
#566805000000
1!
1%
#566810000000
0!
0%
#566815000000
1!
1%
#566820000000
0!
0%
#566825000000
1!
1%
#566830000000
0!
0%
#566835000000
1!
1%
#566840000000
0!
0%
#566845000000
1!
1%
#566850000000
0!
0%
#566855000000
1!
1%
#566860000000
0!
0%
#566865000000
1!
1%
#566870000000
0!
0%
#566875000000
1!
1%
#566880000000
0!
0%
#566885000000
1!
1%
#566890000000
0!
0%
#566895000000
1!
1%
#566900000000
0!
0%
#566905000000
1!
1%
#566910000000
0!
0%
#566915000000
1!
1%
#566920000000
0!
0%
#566925000000
1!
1%
#566930000000
0!
0%
#566935000000
1!
1%
#566940000000
0!
0%
#566945000000
1!
1%
#566950000000
0!
0%
#566955000000
1!
1%
#566960000000
0!
0%
#566965000000
1!
1%
#566970000000
0!
0%
#566975000000
1!
1%
#566980000000
0!
0%
#566985000000
1!
1%
#566990000000
0!
0%
#566995000000
1!
1%
#567000000000
0!
0%
#567005000000
1!
1%
#567010000000
0!
0%
#567015000000
1!
1%
#567020000000
0!
0%
#567025000000
1!
1%
#567030000000
0!
0%
#567035000000
1!
1%
#567040000000
0!
0%
#567045000000
1!
1%
#567050000000
0!
0%
#567055000000
1!
1%
#567060000000
0!
0%
#567065000000
1!
1%
#567070000000
0!
0%
#567075000000
1!
1%
#567080000000
0!
0%
#567085000000
1!
1%
#567090000000
0!
0%
#567095000000
1!
1%
#567100000000
0!
0%
#567105000000
1!
1%
#567110000000
0!
0%
#567115000000
1!
1%
#567120000000
0!
0%
#567125000000
1!
1%
#567130000000
0!
0%
#567135000000
1!
1%
#567140000000
0!
0%
#567145000000
1!
1%
#567150000000
0!
0%
#567155000000
1!
1%
#567160000000
0!
0%
#567165000000
1!
1%
#567170000000
0!
0%
#567175000000
1!
1%
#567180000000
0!
0%
#567185000000
1!
1%
#567190000000
0!
0%
#567195000000
1!
1%
#567200000000
0!
0%
#567205000000
1!
1%
#567210000000
0!
0%
#567215000000
1!
1%
#567220000000
0!
0%
#567225000000
1!
1%
#567230000000
0!
0%
#567235000000
1!
1%
#567240000000
0!
0%
#567245000000
1!
1%
#567250000000
0!
0%
#567255000000
1!
1%
#567260000000
0!
0%
#567265000000
1!
1%
#567270000000
0!
0%
#567275000000
1!
1%
#567280000000
0!
0%
#567285000000
1!
1%
#567290000000
0!
0%
#567295000000
1!
1%
#567300000000
0!
0%
#567305000000
1!
1%
#567310000000
0!
0%
#567315000000
1!
1%
#567320000000
0!
0%
#567325000000
1!
1%
#567330000000
0!
0%
#567335000000
1!
1%
#567340000000
0!
0%
#567345000000
1!
1%
#567350000000
0!
0%
#567355000000
1!
1%
#567360000000
0!
0%
#567365000000
1!
1%
#567370000000
0!
0%
#567375000000
1!
1%
#567380000000
0!
0%
#567385000000
1!
1%
#567390000000
0!
0%
#567395000000
1!
1%
#567400000000
0!
0%
#567405000000
1!
1%
#567410000000
0!
0%
#567415000000
1!
1%
#567420000000
0!
0%
#567425000000
1!
1%
#567430000000
0!
0%
#567435000000
1!
1%
#567440000000
0!
0%
#567445000000
1!
1%
#567450000000
0!
0%
#567455000000
1!
1%
#567460000000
0!
0%
#567465000000
1!
1%
#567470000000
0!
0%
#567475000000
1!
1%
#567480000000
0!
0%
#567485000000
1!
1%
#567490000000
0!
0%
#567495000000
1!
1%
#567500000000
0!
0%
#567505000000
1!
1%
#567510000000
0!
0%
#567515000000
1!
1%
#567520000000
0!
0%
#567525000000
1!
1%
#567530000000
0!
0%
#567535000000
1!
1%
#567540000000
0!
0%
#567545000000
1!
1%
#567550000000
0!
0%
#567555000000
1!
1%
#567560000000
0!
0%
#567565000000
1!
1%
#567570000000
0!
0%
#567575000000
1!
1%
#567580000000
0!
0%
#567585000000
1!
1%
#567590000000
0!
0%
#567595000000
1!
1%
#567600000000
0!
0%
#567605000000
1!
1%
#567610000000
0!
0%
#567615000000
1!
1%
#567620000000
0!
0%
#567625000000
1!
1%
#567630000000
0!
0%
#567635000000
1!
1%
#567640000000
0!
0%
#567645000000
1!
1%
#567650000000
0!
0%
#567655000000
1!
1%
#567660000000
0!
0%
#567665000000
1!
1%
#567670000000
0!
0%
#567675000000
1!
1%
#567680000000
0!
0%
#567685000000
1!
1%
#567690000000
0!
0%
#567695000000
1!
1%
#567700000000
0!
0%
#567705000000
1!
1%
#567710000000
0!
0%
#567715000000
1!
1%
#567720000000
0!
0%
#567725000000
1!
1%
#567730000000
0!
0%
#567735000000
1!
1%
#567740000000
0!
0%
#567745000000
1!
1%
#567750000000
0!
0%
#567755000000
1!
1%
#567760000000
0!
0%
#567765000000
1!
1%
#567770000000
0!
0%
#567775000000
1!
1%
#567780000000
0!
0%
#567785000000
1!
1%
#567790000000
0!
0%
#567795000000
1!
1%
#567800000000
0!
0%
#567805000000
1!
1%
#567810000000
0!
0%
#567815000000
1!
1%
#567820000000
0!
0%
#567825000000
1!
1%
#567830000000
0!
0%
#567835000000
1!
1%
#567840000000
0!
0%
#567845000000
1!
1%
#567850000000
0!
0%
#567855000000
1!
1%
#567860000000
0!
0%
#567865000000
1!
1%
#567870000000
0!
0%
#567875000000
1!
1%
#567880000000
0!
0%
#567885000000
1!
1%
#567890000000
0!
0%
#567895000000
1!
1%
#567900000000
0!
0%
#567905000000
1!
1%
#567910000000
0!
0%
#567915000000
1!
1%
#567920000000
0!
0%
#567925000000
1!
1%
#567930000000
0!
0%
#567935000000
1!
1%
#567940000000
0!
0%
#567945000000
1!
1%
#567950000000
0!
0%
#567955000000
1!
1%
#567960000000
0!
0%
#567965000000
1!
1%
#567970000000
0!
0%
#567975000000
1!
1%
#567980000000
0!
0%
#567985000000
1!
1%
#567990000000
0!
0%
#567995000000
1!
1%
#568000000000
0!
0%
#568005000000
1!
1%
#568010000000
0!
0%
#568015000000
1!
1%
#568020000000
0!
0%
#568025000000
1!
1%
#568030000000
0!
0%
#568035000000
1!
1%
#568040000000
0!
0%
#568045000000
1!
1%
#568050000000
0!
0%
#568055000000
1!
1%
#568060000000
0!
0%
#568065000000
1!
1%
#568070000000
0!
0%
#568075000000
1!
1%
#568080000000
0!
0%
#568085000000
1!
1%
#568090000000
0!
0%
#568095000000
1!
1%
#568100000000
0!
0%
#568105000000
1!
1%
#568110000000
0!
0%
#568115000000
1!
1%
#568120000000
0!
0%
#568125000000
1!
1%
#568130000000
0!
0%
#568135000000
1!
1%
#568140000000
0!
0%
#568145000000
1!
1%
#568150000000
0!
0%
#568155000000
1!
1%
#568160000000
0!
0%
#568165000000
1!
1%
#568170000000
0!
0%
#568175000000
1!
1%
#568180000000
0!
0%
#568185000000
1!
1%
#568190000000
0!
0%
#568195000000
1!
1%
#568200000000
0!
0%
#568205000000
1!
1%
#568210000000
0!
0%
#568215000000
1!
1%
#568220000000
0!
0%
#568225000000
1!
1%
#568230000000
0!
0%
#568235000000
1!
1%
#568240000000
0!
0%
#568245000000
1!
1%
#568250000000
0!
0%
#568255000000
1!
1%
#568260000000
0!
0%
#568265000000
1!
1%
#568270000000
0!
0%
#568275000000
1!
1%
#568280000000
0!
0%
#568285000000
1!
1%
#568290000000
0!
0%
#568295000000
1!
1%
#568300000000
0!
0%
#568305000000
1!
1%
#568310000000
0!
0%
#568315000000
1!
1%
#568320000000
0!
0%
#568325000000
1!
1%
#568330000000
0!
0%
#568335000000
1!
1%
#568340000000
0!
0%
#568345000000
1!
1%
#568350000000
0!
0%
#568355000000
1!
1%
#568360000000
0!
0%
#568365000000
1!
1%
#568370000000
0!
0%
#568375000000
1!
1%
#568380000000
0!
0%
#568385000000
1!
1%
#568390000000
0!
0%
#568395000000
1!
1%
#568400000000
0!
0%
#568405000000
1!
1%
#568410000000
0!
0%
#568415000000
1!
1%
#568420000000
0!
0%
#568425000000
1!
1%
#568430000000
0!
0%
#568435000000
1!
1%
#568440000000
0!
0%
#568445000000
1!
1%
#568450000000
0!
0%
#568455000000
1!
1%
#568460000000
0!
0%
#568465000000
1!
1%
#568470000000
0!
0%
#568475000000
1!
1%
#568480000000
0!
0%
#568485000000
1!
1%
#568490000000
0!
0%
#568495000000
1!
1%
#568500000000
0!
0%
#568505000000
1!
1%
#568510000000
0!
0%
#568515000000
1!
1%
#568520000000
0!
0%
#568525000000
1!
1%
#568530000000
0!
0%
#568535000000
1!
1%
#568540000000
0!
0%
#568545000000
1!
1%
#568550000000
0!
0%
#568555000000
1!
1%
#568560000000
0!
0%
#568565000000
1!
1%
#568570000000
0!
0%
#568575000000
1!
1%
#568580000000
0!
0%
#568585000000
1!
1%
#568590000000
0!
0%
#568595000000
1!
1%
#568600000000
0!
0%
#568605000000
1!
1%
#568610000000
0!
0%
#568615000000
1!
1%
#568620000000
0!
0%
#568625000000
1!
1%
#568630000000
0!
0%
#568635000000
1!
1%
#568640000000
0!
0%
#568645000000
1!
1%
#568650000000
0!
0%
#568655000000
1!
1%
#568660000000
0!
0%
#568665000000
1!
1%
#568670000000
0!
0%
#568675000000
1!
1%
#568680000000
0!
0%
#568685000000
1!
1%
#568690000000
0!
0%
#568695000000
1!
1%
#568700000000
0!
0%
#568705000000
1!
1%
#568710000000
0!
0%
#568715000000
1!
1%
#568720000000
0!
0%
#568725000000
1!
1%
#568730000000
0!
0%
#568735000000
1!
1%
#568740000000
0!
0%
#568745000000
1!
1%
#568750000000
0!
0%
#568755000000
1!
1%
#568760000000
0!
0%
#568765000000
1!
1%
#568770000000
0!
0%
#568775000000
1!
1%
#568780000000
0!
0%
#568785000000
1!
1%
#568790000000
0!
0%
#568795000000
1!
1%
#568800000000
0!
0%
#568805000000
1!
1%
#568810000000
0!
0%
#568815000000
1!
1%
#568820000000
0!
0%
#568825000000
1!
1%
#568830000000
0!
0%
#568835000000
1!
1%
#568840000000
0!
0%
#568845000000
1!
1%
#568850000000
0!
0%
#568855000000
1!
1%
#568860000000
0!
0%
#568865000000
1!
1%
#568870000000
0!
0%
#568875000000
1!
1%
#568880000000
0!
0%
#568885000000
1!
1%
#568890000000
0!
0%
#568895000000
1!
1%
#568900000000
0!
0%
#568905000000
1!
1%
#568910000000
0!
0%
#568915000000
1!
1%
#568920000000
0!
0%
#568925000000
1!
1%
#568930000000
0!
0%
#568935000000
1!
1%
#568940000000
0!
0%
#568945000000
1!
1%
#568950000000
0!
0%
#568955000000
1!
1%
#568960000000
0!
0%
#568965000000
1!
1%
#568970000000
0!
0%
#568975000000
1!
1%
#568980000000
0!
0%
#568985000000
1!
1%
#568990000000
0!
0%
#568995000000
1!
1%
#569000000000
0!
0%
#569005000000
1!
1%
#569010000000
0!
0%
#569015000000
1!
1%
#569020000000
0!
0%
#569025000000
1!
1%
#569030000000
0!
0%
#569035000000
1!
1%
#569040000000
0!
0%
#569045000000
1!
1%
#569050000000
0!
0%
#569055000000
1!
1%
#569060000000
0!
0%
#569065000000
1!
1%
#569070000000
0!
0%
#569075000000
1!
1%
#569080000000
0!
0%
#569085000000
1!
1%
#569090000000
0!
0%
#569095000000
1!
1%
#569100000000
0!
0%
#569105000000
1!
1%
#569110000000
0!
0%
#569115000000
1!
1%
#569120000000
0!
0%
#569125000000
1!
1%
#569130000000
0!
0%
#569135000000
1!
1%
#569140000000
0!
0%
#569145000000
1!
1%
#569150000000
0!
0%
#569155000000
1!
1%
#569160000000
0!
0%
#569165000000
1!
1%
#569170000000
0!
0%
#569175000000
1!
1%
#569180000000
0!
0%
#569185000000
1!
1%
#569190000000
0!
0%
#569195000000
1!
1%
#569200000000
0!
0%
#569205000000
1!
1%
#569210000000
0!
0%
#569215000000
1!
1%
#569220000000
0!
0%
#569225000000
1!
1%
#569230000000
0!
0%
#569235000000
1!
1%
#569240000000
0!
0%
#569245000000
1!
1%
#569250000000
0!
0%
#569255000000
1!
1%
#569260000000
0!
0%
#569265000000
1!
1%
#569270000000
0!
0%
#569275000000
1!
1%
#569280000000
0!
0%
#569285000000
1!
1%
#569290000000
0!
0%
#569295000000
1!
1%
#569300000000
0!
0%
#569305000000
1!
1%
#569310000000
0!
0%
#569315000000
1!
1%
#569320000000
0!
0%
#569325000000
1!
1%
#569330000000
0!
0%
#569335000000
1!
1%
#569340000000
0!
0%
#569345000000
1!
1%
#569350000000
0!
0%
#569355000000
1!
1%
#569360000000
0!
0%
#569365000000
1!
1%
#569370000000
0!
0%
#569375000000
1!
1%
#569380000000
0!
0%
#569385000000
1!
1%
#569390000000
0!
0%
#569395000000
1!
1%
#569400000000
0!
0%
#569405000000
1!
1%
#569410000000
0!
0%
#569415000000
1!
1%
#569420000000
0!
0%
#569425000000
1!
1%
#569430000000
0!
0%
#569435000000
1!
1%
#569440000000
0!
0%
#569445000000
1!
1%
#569450000000
0!
0%
#569455000000
1!
1%
#569460000000
0!
0%
#569465000000
1!
1%
#569470000000
0!
0%
#569475000000
1!
1%
#569480000000
0!
0%
#569485000000
1!
1%
#569490000000
0!
0%
#569495000000
1!
1%
#569500000000
0!
0%
#569505000000
1!
1%
#569510000000
0!
0%
#569515000000
1!
1%
#569520000000
0!
0%
#569525000000
1!
1%
#569530000000
0!
0%
#569535000000
1!
1%
#569540000000
0!
0%
#569545000000
1!
1%
#569550000000
0!
0%
#569555000000
1!
1%
#569560000000
0!
0%
#569565000000
1!
1%
#569570000000
0!
0%
#569575000000
1!
1%
#569580000000
0!
0%
#569585000000
1!
1%
#569590000000
0!
0%
#569595000000
1!
1%
#569600000000
0!
0%
#569605000000
1!
1%
#569610000000
0!
0%
#569615000000
1!
1%
#569620000000
0!
0%
#569625000000
1!
1%
#569630000000
0!
0%
#569635000000
1!
1%
#569640000000
0!
0%
#569645000000
1!
1%
#569650000000
0!
0%
#569655000000
1!
1%
#569660000000
0!
0%
#569665000000
1!
1%
#569670000000
0!
0%
#569675000000
1!
1%
#569680000000
0!
0%
#569685000000
1!
1%
#569690000000
0!
0%
#569695000000
1!
1%
#569700000000
0!
0%
#569705000000
1!
1%
#569710000000
0!
0%
#569715000000
1!
1%
#569720000000
0!
0%
#569725000000
1!
1%
#569730000000
0!
0%
#569735000000
1!
1%
#569740000000
0!
0%
#569745000000
1!
1%
#569750000000
0!
0%
#569755000000
1!
1%
#569760000000
0!
0%
#569765000000
1!
1%
#569770000000
0!
0%
#569775000000
1!
1%
#569780000000
0!
0%
#569785000000
1!
1%
#569790000000
0!
0%
#569795000000
1!
1%
#569800000000
0!
0%
#569805000000
1!
1%
#569810000000
0!
0%
#569815000000
1!
1%
#569820000000
0!
0%
#569825000000
1!
1%
#569830000000
0!
0%
#569835000000
1!
1%
#569840000000
0!
0%
#569845000000
1!
1%
#569850000000
0!
0%
#569855000000
1!
1%
#569860000000
0!
0%
#569865000000
1!
1%
#569870000000
0!
0%
#569875000000
1!
1%
#569880000000
0!
0%
#569885000000
1!
1%
#569890000000
0!
0%
#569895000000
1!
1%
#569900000000
0!
0%
#569905000000
1!
1%
#569910000000
0!
0%
#569915000000
1!
1%
#569920000000
0!
0%
#569925000000
1!
1%
#569930000000
0!
0%
#569935000000
1!
1%
#569940000000
0!
0%
#569945000000
1!
1%
#569950000000
0!
0%
#569955000000
1!
1%
#569960000000
0!
0%
#569965000000
1!
1%
#569970000000
0!
0%
#569975000000
1!
1%
#569980000000
0!
0%
#569985000000
1!
1%
#569990000000
0!
0%
#569995000000
1!
1%
#570000000000
0!
0%
#570005000000
1!
1%
#570010000000
0!
0%
#570015000000
1!
1%
#570020000000
0!
0%
#570025000000
1!
1%
#570030000000
0!
0%
#570035000000
1!
1%
#570040000000
0!
0%
#570045000000
1!
1%
#570050000000
0!
0%
#570055000000
1!
1%
#570060000000
0!
0%
#570065000000
1!
1%
#570070000000
0!
0%
#570075000000
1!
1%
#570080000000
0!
0%
#570085000000
1!
1%
#570090000000
0!
0%
#570095000000
1!
1%
#570100000000
0!
0%
#570105000000
1!
1%
#570110000000
0!
0%
#570115000000
1!
1%
#570120000000
0!
0%
#570125000000
1!
1%
#570130000000
0!
0%
#570135000000
1!
1%
#570140000000
0!
0%
#570145000000
1!
1%
#570150000000
0!
0%
#570155000000
1!
1%
#570160000000
0!
0%
#570165000000
1!
1%
#570170000000
0!
0%
#570175000000
1!
1%
#570180000000
0!
0%
#570185000000
1!
1%
#570190000000
0!
0%
#570195000000
1!
1%
#570200000000
0!
0%
#570205000000
1!
1%
#570210000000
0!
0%
#570215000000
1!
1%
#570220000000
0!
0%
#570225000000
1!
1%
#570230000000
0!
0%
#570235000000
1!
1%
#570240000000
0!
0%
#570245000000
1!
1%
#570250000000
0!
0%
#570255000000
1!
1%
#570260000000
0!
0%
#570265000000
1!
1%
#570270000000
0!
0%
#570275000000
1!
1%
#570280000000
0!
0%
#570285000000
1!
1%
#570290000000
0!
0%
#570295000000
1!
1%
#570300000000
0!
0%
#570305000000
1!
1%
#570310000000
0!
0%
#570315000000
1!
1%
#570320000000
0!
0%
#570325000000
1!
1%
#570330000000
0!
0%
#570335000000
1!
1%
#570340000000
0!
0%
#570345000000
1!
1%
#570350000000
0!
0%
#570355000000
1!
1%
#570360000000
0!
0%
#570365000000
1!
1%
#570370000000
0!
0%
#570375000000
1!
1%
#570380000000
0!
0%
#570385000000
1!
1%
#570390000000
0!
0%
#570395000000
1!
1%
#570400000000
0!
0%
#570405000000
1!
1%
#570410000000
0!
0%
#570415000000
1!
1%
#570420000000
0!
0%
#570425000000
1!
1%
#570430000000
0!
0%
#570435000000
1!
1%
#570440000000
0!
0%
#570445000000
1!
1%
#570450000000
0!
0%
#570455000000
1!
1%
#570460000000
0!
0%
#570465000000
1!
1%
#570470000000
0!
0%
#570475000000
1!
1%
#570480000000
0!
0%
#570485000000
1!
1%
#570490000000
0!
0%
#570495000000
1!
1%
#570500000000
0!
0%
#570505000000
1!
1%
#570510000000
0!
0%
#570515000000
1!
1%
#570520000000
0!
0%
#570525000000
1!
1%
#570530000000
0!
0%
#570535000000
1!
1%
#570540000000
0!
0%
#570545000000
1!
1%
#570550000000
0!
0%
#570555000000
1!
1%
#570560000000
0!
0%
#570565000000
1!
1%
#570570000000
0!
0%
#570575000000
1!
1%
#570580000000
0!
0%
#570585000000
1!
1%
#570590000000
0!
0%
#570595000000
1!
1%
#570600000000
0!
0%
#570605000000
1!
1%
#570610000000
0!
0%
#570615000000
1!
1%
#570620000000
0!
0%
#570625000000
1!
1%
#570630000000
0!
0%
#570635000000
1!
1%
#570640000000
0!
0%
#570645000000
1!
1%
#570650000000
0!
0%
#570655000000
1!
1%
#570660000000
0!
0%
#570665000000
1!
1%
#570670000000
0!
0%
#570675000000
1!
1%
#570680000000
0!
0%
#570685000000
1!
1%
#570690000000
0!
0%
#570695000000
1!
1%
#570700000000
0!
0%
#570705000000
1!
1%
#570710000000
0!
0%
#570715000000
1!
1%
#570720000000
0!
0%
#570725000000
1!
1%
#570730000000
0!
0%
#570735000000
1!
1%
#570740000000
0!
0%
#570745000000
1!
1%
#570750000000
0!
0%
#570755000000
1!
1%
#570760000000
0!
0%
#570765000000
1!
1%
#570770000000
0!
0%
#570775000000
1!
1%
#570780000000
0!
0%
#570785000000
1!
1%
#570790000000
0!
0%
#570795000000
1!
1%
#570800000000
0!
0%
#570805000000
1!
1%
#570810000000
0!
0%
#570815000000
1!
1%
#570820000000
0!
0%
#570825000000
1!
1%
#570830000000
0!
0%
#570835000000
1!
1%
#570840000000
0!
0%
#570845000000
1!
1%
#570850000000
0!
0%
#570855000000
1!
1%
#570860000000
0!
0%
#570865000000
1!
1%
#570870000000
0!
0%
#570875000000
1!
1%
#570880000000
0!
0%
#570885000000
1!
1%
#570890000000
0!
0%
#570895000000
1!
1%
#570900000000
0!
0%
#570905000000
1!
1%
#570910000000
0!
0%
#570915000000
1!
1%
#570920000000
0!
0%
#570925000000
1!
1%
#570930000000
0!
0%
#570935000000
1!
1%
#570940000000
0!
0%
#570945000000
1!
1%
#570950000000
0!
0%
#570955000000
1!
1%
#570960000000
0!
0%
#570965000000
1!
1%
#570970000000
0!
0%
#570975000000
1!
1%
#570980000000
0!
0%
#570985000000
1!
1%
#570990000000
0!
0%
#570995000000
1!
1%
#571000000000
0!
0%
#571005000000
1!
1%
#571010000000
0!
0%
#571015000000
1!
1%
#571020000000
0!
0%
#571025000000
1!
1%
#571030000000
0!
0%
#571035000000
1!
1%
#571040000000
0!
0%
#571045000000
1!
1%
#571050000000
0!
0%
#571055000000
1!
1%
#571060000000
0!
0%
#571065000000
1!
1%
#571070000000
0!
0%
#571075000000
1!
1%
#571080000000
0!
0%
#571085000000
1!
1%
#571090000000
0!
0%
#571095000000
1!
1%
#571100000000
0!
0%
#571105000000
1!
1%
#571110000000
0!
0%
#571115000000
1!
1%
#571120000000
0!
0%
#571125000000
1!
1%
#571130000000
0!
0%
#571135000000
1!
1%
#571140000000
0!
0%
#571145000000
1!
1%
#571150000000
0!
0%
#571155000000
1!
1%
#571160000000
0!
0%
#571165000000
1!
1%
#571170000000
0!
0%
#571175000000
1!
1%
#571180000000
0!
0%
#571185000000
1!
1%
#571190000000
0!
0%
#571195000000
1!
1%
#571200000000
0!
0%
#571205000000
1!
1%
#571210000000
0!
0%
#571215000000
1!
1%
#571220000000
0!
0%
#571225000000
1!
1%
#571230000000
0!
0%
#571235000000
1!
1%
#571240000000
0!
0%
#571245000000
1!
1%
#571250000000
0!
0%
#571255000000
1!
1%
#571260000000
0!
0%
#571265000000
1!
1%
#571270000000
0!
0%
#571275000000
1!
1%
#571280000000
0!
0%
#571285000000
1!
1%
#571290000000
0!
0%
#571295000000
1!
1%
#571300000000
0!
0%
#571305000000
1!
1%
#571310000000
0!
0%
#571315000000
1!
1%
#571320000000
0!
0%
#571325000000
1!
1%
#571330000000
0!
0%
#571335000000
1!
1%
#571340000000
0!
0%
#571345000000
1!
1%
#571350000000
0!
0%
#571355000000
1!
1%
#571360000000
0!
0%
#571365000000
1!
1%
#571370000000
0!
0%
#571375000000
1!
1%
#571380000000
0!
0%
#571385000000
1!
1%
#571390000000
0!
0%
#571395000000
1!
1%
#571400000000
0!
0%
#571405000000
1!
1%
#571410000000
0!
0%
#571415000000
1!
1%
#571420000000
0!
0%
#571425000000
1!
1%
#571430000000
0!
0%
#571435000000
1!
1%
#571440000000
0!
0%
#571445000000
1!
1%
#571450000000
0!
0%
#571455000000
1!
1%
#571460000000
0!
0%
#571465000000
1!
1%
#571470000000
0!
0%
#571475000000
1!
1%
#571480000000
0!
0%
#571485000000
1!
1%
#571490000000
0!
0%
#571495000000
1!
1%
#571500000000
0!
0%
#571505000000
1!
1%
#571510000000
0!
0%
#571515000000
1!
1%
#571520000000
0!
0%
#571525000000
1!
1%
#571530000000
0!
0%
#571535000000
1!
1%
#571540000000
0!
0%
#571545000000
1!
1%
#571550000000
0!
0%
#571555000000
1!
1%
#571560000000
0!
0%
#571565000000
1!
1%
#571570000000
0!
0%
#571575000000
1!
1%
#571580000000
0!
0%
#571585000000
1!
1%
#571590000000
0!
0%
#571595000000
1!
1%
#571600000000
0!
0%
#571605000000
1!
1%
#571610000000
0!
0%
#571615000000
1!
1%
#571620000000
0!
0%
#571625000000
1!
1%
#571630000000
0!
0%
#571635000000
1!
1%
#571640000000
0!
0%
#571645000000
1!
1%
#571650000000
0!
0%
#571655000000
1!
1%
#571660000000
0!
0%
#571665000000
1!
1%
#571670000000
0!
0%
#571675000000
1!
1%
#571680000000
0!
0%
#571685000000
1!
1%
#571690000000
0!
0%
#571695000000
1!
1%
#571700000000
0!
0%
#571705000000
1!
1%
#571710000000
0!
0%
#571715000000
1!
1%
#571720000000
0!
0%
#571725000000
1!
1%
#571730000000
0!
0%
#571735000000
1!
1%
#571740000000
0!
0%
#571745000000
1!
1%
#571750000000
0!
0%
#571755000000
1!
1%
#571760000000
0!
0%
#571765000000
1!
1%
#571770000000
0!
0%
#571775000000
1!
1%
#571780000000
0!
0%
#571785000000
1!
1%
#571790000000
0!
0%
#571795000000
1!
1%
#571800000000
0!
0%
#571805000000
1!
1%
#571810000000
0!
0%
#571815000000
1!
1%
#571820000000
0!
0%
#571825000000
1!
1%
#571830000000
0!
0%
#571835000000
1!
1%
#571840000000
0!
0%
#571845000000
1!
1%
#571850000000
0!
0%
#571855000000
1!
1%
#571860000000
0!
0%
#571865000000
1!
1%
#571870000000
0!
0%
#571875000000
1!
1%
#571880000000
0!
0%
#571885000000
1!
1%
#571890000000
0!
0%
#571895000000
1!
1%
#571900000000
0!
0%
#571905000000
1!
1%
#571910000000
0!
0%
#571915000000
1!
1%
#571920000000
0!
0%
#571925000000
1!
1%
#571930000000
0!
0%
#571935000000
1!
1%
#571940000000
0!
0%
#571945000000
1!
1%
#571950000000
0!
0%
#571955000000
1!
1%
#571960000000
0!
0%
#571965000000
1!
1%
#571970000000
0!
0%
#571975000000
1!
1%
#571980000000
0!
0%
#571985000000
1!
1%
#571990000000
0!
0%
#571995000000
1!
1%
#572000000000
0!
0%
#572005000000
1!
1%
#572010000000
0!
0%
#572015000000
1!
1%
#572020000000
0!
0%
#572025000000
1!
1%
#572030000000
0!
0%
#572035000000
1!
1%
#572040000000
0!
0%
#572045000000
1!
1%
#572050000000
0!
0%
#572055000000
1!
1%
#572060000000
0!
0%
#572065000000
1!
1%
#572070000000
0!
0%
#572075000000
1!
1%
#572080000000
0!
0%
#572085000000
1!
1%
#572090000000
0!
0%
#572095000000
1!
1%
#572100000000
0!
0%
#572105000000
1!
1%
#572110000000
0!
0%
#572115000000
1!
1%
#572120000000
0!
0%
#572125000000
1!
1%
#572130000000
0!
0%
#572135000000
1!
1%
#572140000000
0!
0%
#572145000000
1!
1%
#572150000000
0!
0%
#572155000000
1!
1%
#572160000000
0!
0%
#572165000000
1!
1%
#572170000000
0!
0%
#572175000000
1!
1%
#572180000000
0!
0%
#572185000000
1!
1%
#572190000000
0!
0%
#572195000000
1!
1%
#572200000000
0!
0%
#572205000000
1!
1%
#572210000000
0!
0%
#572215000000
1!
1%
#572220000000
0!
0%
#572225000000
1!
1%
#572230000000
0!
0%
#572235000000
1!
1%
#572240000000
0!
0%
#572245000000
1!
1%
#572250000000
0!
0%
#572255000000
1!
1%
#572260000000
0!
0%
#572265000000
1!
1%
#572270000000
0!
0%
#572275000000
1!
1%
#572280000000
0!
0%
#572285000000
1!
1%
#572290000000
0!
0%
#572295000000
1!
1%
#572300000000
0!
0%
#572305000000
1!
1%
#572310000000
0!
0%
#572315000000
1!
1%
#572320000000
0!
0%
#572325000000
1!
1%
#572330000000
0!
0%
#572335000000
1!
1%
#572340000000
0!
0%
#572345000000
1!
1%
#572350000000
0!
0%
#572355000000
1!
1%
#572360000000
0!
0%
#572365000000
1!
1%
#572370000000
0!
0%
#572375000000
1!
1%
#572380000000
0!
0%
#572385000000
1!
1%
#572390000000
0!
0%
#572395000000
1!
1%
#572400000000
0!
0%
#572405000000
1!
1%
#572410000000
0!
0%
#572415000000
1!
1%
#572420000000
0!
0%
#572425000000
1!
1%
#572430000000
0!
0%
#572435000000
1!
1%
#572440000000
0!
0%
#572445000000
1!
1%
#572450000000
0!
0%
#572455000000
1!
1%
#572460000000
0!
0%
#572465000000
1!
1%
#572470000000
0!
0%
#572475000000
1!
1%
#572480000000
0!
0%
#572485000000
1!
1%
#572490000000
0!
0%
#572495000000
1!
1%
#572500000000
0!
0%
#572505000000
1!
1%
#572510000000
0!
0%
#572515000000
1!
1%
#572520000000
0!
0%
#572525000000
1!
1%
#572530000000
0!
0%
#572535000000
1!
1%
#572540000000
0!
0%
#572545000000
1!
1%
#572550000000
0!
0%
#572555000000
1!
1%
#572560000000
0!
0%
#572565000000
1!
1%
#572570000000
0!
0%
#572575000000
1!
1%
#572580000000
0!
0%
#572585000000
1!
1%
#572590000000
0!
0%
#572595000000
1!
1%
#572600000000
0!
0%
#572605000000
1!
1%
#572610000000
0!
0%
#572615000000
1!
1%
#572620000000
0!
0%
#572625000000
1!
1%
#572630000000
0!
0%
#572635000000
1!
1%
#572640000000
0!
0%
#572645000000
1!
1%
#572650000000
0!
0%
#572655000000
1!
1%
#572660000000
0!
0%
#572665000000
1!
1%
#572670000000
0!
0%
#572675000000
1!
1%
#572680000000
0!
0%
#572685000000
1!
1%
#572690000000
0!
0%
#572695000000
1!
1%
#572700000000
0!
0%
#572705000000
1!
1%
#572710000000
0!
0%
#572715000000
1!
1%
#572720000000
0!
0%
#572725000000
1!
1%
#572730000000
0!
0%
#572735000000
1!
1%
#572740000000
0!
0%
#572745000000
1!
1%
#572750000000
0!
0%
#572755000000
1!
1%
#572760000000
0!
0%
#572765000000
1!
1%
#572770000000
0!
0%
#572775000000
1!
1%
#572780000000
0!
0%
#572785000000
1!
1%
#572790000000
0!
0%
#572795000000
1!
1%
#572800000000
0!
0%
#572805000000
1!
1%
#572810000000
0!
0%
#572815000000
1!
1%
#572820000000
0!
0%
#572825000000
1!
1%
#572830000000
0!
0%
#572835000000
1!
1%
#572840000000
0!
0%
#572845000000
1!
1%
#572850000000
0!
0%
#572855000000
1!
1%
#572860000000
0!
0%
#572865000000
1!
1%
#572870000000
0!
0%
#572875000000
1!
1%
#572880000000
0!
0%
#572885000000
1!
1%
#572890000000
0!
0%
#572895000000
1!
1%
#572900000000
0!
0%
#572905000000
1!
1%
#572910000000
0!
0%
#572915000000
1!
1%
#572920000000
0!
0%
#572925000000
1!
1%
#572930000000
0!
0%
#572935000000
1!
1%
#572940000000
0!
0%
#572945000000
1!
1%
#572950000000
0!
0%
#572955000000
1!
1%
#572960000000
0!
0%
#572965000000
1!
1%
#572970000000
0!
0%
#572975000000
1!
1%
#572980000000
0!
0%
#572985000000
1!
1%
#572990000000
0!
0%
#572995000000
1!
1%
#573000000000
0!
0%
#573005000000
1!
1%
#573010000000
0!
0%
#573015000000
1!
1%
#573020000000
0!
0%
#573025000000
1!
1%
#573030000000
0!
0%
#573035000000
1!
1%
#573040000000
0!
0%
#573045000000
1!
1%
#573050000000
0!
0%
#573055000000
1!
1%
#573060000000
0!
0%
#573065000000
1!
1%
#573070000000
0!
0%
#573075000000
1!
1%
#573080000000
0!
0%
#573085000000
1!
1%
#573090000000
0!
0%
#573095000000
1!
1%
#573100000000
0!
0%
#573105000000
1!
1%
#573110000000
0!
0%
#573115000000
1!
1%
#573120000000
0!
0%
#573125000000
1!
1%
#573130000000
0!
0%
#573135000000
1!
1%
#573140000000
0!
0%
#573145000000
1!
1%
#573150000000
0!
0%
#573155000000
1!
1%
#573160000000
0!
0%
#573165000000
1!
1%
#573170000000
0!
0%
#573175000000
1!
1%
#573180000000
0!
0%
#573185000000
1!
1%
#573190000000
0!
0%
#573195000000
1!
1%
#573200000000
0!
0%
#573205000000
1!
1%
#573210000000
0!
0%
#573215000000
1!
1%
#573220000000
0!
0%
#573225000000
1!
1%
#573230000000
0!
0%
#573235000000
1!
1%
#573240000000
0!
0%
#573245000000
1!
1%
#573250000000
0!
0%
#573255000000
1!
1%
#573260000000
0!
0%
#573265000000
1!
1%
#573270000000
0!
0%
#573275000000
1!
1%
#573280000000
0!
0%
#573285000000
1!
1%
#573290000000
0!
0%
#573295000000
1!
1%
#573300000000
0!
0%
#573305000000
1!
1%
#573310000000
0!
0%
#573315000000
1!
1%
#573320000000
0!
0%
#573325000000
1!
1%
#573330000000
0!
0%
#573335000000
1!
1%
#573340000000
0!
0%
#573345000000
1!
1%
#573350000000
0!
0%
#573355000000
1!
1%
#573360000000
0!
0%
#573365000000
1!
1%
#573370000000
0!
0%
#573375000000
1!
1%
#573380000000
0!
0%
#573385000000
1!
1%
#573390000000
0!
0%
#573395000000
1!
1%
#573400000000
0!
0%
#573405000000
1!
1%
#573410000000
0!
0%
#573415000000
1!
1%
#573420000000
0!
0%
#573425000000
1!
1%
#573430000000
0!
0%
#573435000000
1!
1%
#573440000000
0!
0%
#573445000000
1!
1%
#573450000000
0!
0%
#573455000000
1!
1%
#573460000000
0!
0%
#573465000000
1!
1%
#573470000000
0!
0%
#573475000000
1!
1%
#573480000000
0!
0%
#573485000000
1!
1%
#573490000000
0!
0%
#573495000000
1!
1%
#573500000000
0!
0%
#573505000000
1!
1%
#573510000000
0!
0%
#573515000000
1!
1%
#573520000000
0!
0%
#573525000000
1!
1%
#573530000000
0!
0%
#573535000000
1!
1%
#573540000000
0!
0%
#573545000000
1!
1%
#573550000000
0!
0%
#573555000000
1!
1%
#573560000000
0!
0%
#573565000000
1!
1%
#573570000000
0!
0%
#573575000000
1!
1%
#573580000000
0!
0%
#573585000000
1!
1%
#573590000000
0!
0%
#573595000000
1!
1%
#573600000000
0!
0%
#573605000000
1!
1%
#573610000000
0!
0%
#573615000000
1!
1%
#573620000000
0!
0%
#573625000000
1!
1%
#573630000000
0!
0%
#573635000000
1!
1%
#573640000000
0!
0%
#573645000000
1!
1%
#573650000000
0!
0%
#573655000000
1!
1%
#573660000000
0!
0%
#573665000000
1!
1%
#573670000000
0!
0%
#573675000000
1!
1%
#573680000000
0!
0%
#573685000000
1!
1%
#573690000000
0!
0%
#573695000000
1!
1%
#573700000000
0!
0%
#573705000000
1!
1%
#573710000000
0!
0%
#573715000000
1!
1%
#573720000000
0!
0%
#573725000000
1!
1%
#573730000000
0!
0%
#573735000000
1!
1%
#573740000000
0!
0%
#573745000000
1!
1%
#573750000000
0!
0%
#573755000000
1!
1%
#573760000000
0!
0%
#573765000000
1!
1%
#573770000000
0!
0%
#573775000000
1!
1%
#573780000000
0!
0%
#573785000000
1!
1%
#573790000000
0!
0%
#573795000000
1!
1%
#573800000000
0!
0%
#573805000000
1!
1%
#573810000000
0!
0%
#573815000000
1!
1%
#573820000000
0!
0%
#573825000000
1!
1%
#573830000000
0!
0%
#573835000000
1!
1%
#573840000000
0!
0%
#573845000000
1!
1%
#573850000000
0!
0%
#573855000000
1!
1%
#573860000000
0!
0%
#573865000000
1!
1%
#573870000000
0!
0%
#573875000000
1!
1%
#573880000000
0!
0%
#573885000000
1!
1%
#573890000000
0!
0%
#573895000000
1!
1%
#573900000000
0!
0%
#573905000000
1!
1%
#573910000000
0!
0%
#573915000000
1!
1%
#573920000000
0!
0%
#573925000000
1!
1%
#573930000000
0!
0%
#573935000000
1!
1%
#573940000000
0!
0%
#573945000000
1!
1%
#573950000000
0!
0%
#573955000000
1!
1%
#573960000000
0!
0%
#573965000000
1!
1%
#573970000000
0!
0%
#573975000000
1!
1%
#573980000000
0!
0%
#573985000000
1!
1%
#573990000000
0!
0%
#573995000000
1!
1%
#574000000000
0!
0%
#574005000000
1!
1%
#574010000000
0!
0%
#574015000000
1!
1%
#574020000000
0!
0%
#574025000000
1!
1%
#574030000000
0!
0%
#574035000000
1!
1%
#574040000000
0!
0%
#574045000000
1!
1%
#574050000000
0!
0%
#574055000000
1!
1%
#574060000000
0!
0%
#574065000000
1!
1%
#574070000000
0!
0%
#574075000000
1!
1%
#574080000000
0!
0%
#574085000000
1!
1%
#574090000000
0!
0%
#574095000000
1!
1%
#574100000000
0!
0%
#574105000000
1!
1%
#574110000000
0!
0%
#574115000000
1!
1%
#574120000000
0!
0%
#574125000000
1!
1%
#574130000000
0!
0%
#574135000000
1!
1%
#574140000000
0!
0%
#574145000000
1!
1%
#574150000000
0!
0%
#574155000000
1!
1%
#574160000000
0!
0%
#574165000000
1!
1%
#574170000000
0!
0%
#574175000000
1!
1%
#574180000000
0!
0%
#574185000000
1!
1%
#574190000000
0!
0%
#574195000000
1!
1%
#574200000000
0!
0%
#574205000000
1!
1%
#574210000000
0!
0%
#574215000000
1!
1%
#574220000000
0!
0%
#574225000000
1!
1%
#574230000000
0!
0%
#574235000000
1!
1%
#574240000000
0!
0%
#574245000000
1!
1%
#574250000000
0!
0%
#574255000000
1!
1%
#574260000000
0!
0%
#574265000000
1!
1%
#574270000000
0!
0%
#574275000000
1!
1%
#574280000000
0!
0%
#574285000000
1!
1%
#574290000000
0!
0%
#574295000000
1!
1%
#574300000000
0!
0%
#574305000000
1!
1%
#574310000000
0!
0%
#574315000000
1!
1%
#574320000000
0!
0%
#574325000000
1!
1%
#574330000000
0!
0%
#574335000000
1!
1%
#574340000000
0!
0%
#574345000000
1!
1%
#574350000000
0!
0%
#574355000000
1!
1%
#574360000000
0!
0%
#574365000000
1!
1%
#574370000000
0!
0%
#574375000000
1!
1%
#574380000000
0!
0%
#574385000000
1!
1%
#574390000000
0!
0%
#574395000000
1!
1%
#574400000000
0!
0%
#574405000000
1!
1%
#574410000000
0!
0%
#574415000000
1!
1%
#574420000000
0!
0%
#574425000000
1!
1%
#574430000000
0!
0%
#574435000000
1!
1%
#574440000000
0!
0%
#574445000000
1!
1%
#574450000000
0!
0%
#574455000000
1!
1%
#574460000000
0!
0%
#574465000000
1!
1%
#574470000000
0!
0%
#574475000000
1!
1%
#574480000000
0!
0%
#574485000000
1!
1%
#574490000000
0!
0%
#574495000000
1!
1%
#574500000000
0!
0%
#574505000000
1!
1%
#574510000000
0!
0%
#574515000000
1!
1%
#574520000000
0!
0%
#574525000000
1!
1%
#574530000000
0!
0%
#574535000000
1!
1%
#574540000000
0!
0%
#574545000000
1!
1%
#574550000000
0!
0%
#574555000000
1!
1%
#574560000000
0!
0%
#574565000000
1!
1%
#574570000000
0!
0%
#574575000000
1!
1%
#574580000000
0!
0%
#574585000000
1!
1%
#574590000000
0!
0%
#574595000000
1!
1%
#574600000000
0!
0%
#574605000000
1!
1%
#574610000000
0!
0%
#574615000000
1!
1%
#574620000000
0!
0%
#574625000000
1!
1%
#574630000000
0!
0%
#574635000000
1!
1%
#574640000000
0!
0%
#574645000000
1!
1%
#574650000000
0!
0%
#574655000000
1!
1%
#574660000000
0!
0%
#574665000000
1!
1%
#574670000000
0!
0%
#574675000000
1!
1%
#574680000000
0!
0%
#574685000000
1!
1%
#574690000000
0!
0%
#574695000000
1!
1%
#574700000000
0!
0%
#574705000000
1!
1%
#574710000000
0!
0%
#574715000000
1!
1%
#574720000000
0!
0%
#574725000000
1!
1%
#574730000000
0!
0%
#574735000000
1!
1%
#574740000000
0!
0%
#574745000000
1!
1%
#574750000000
0!
0%
#574755000000
1!
1%
#574760000000
0!
0%
#574765000000
1!
1%
#574770000000
0!
0%
#574775000000
1!
1%
#574780000000
0!
0%
#574785000000
1!
1%
#574790000000
0!
0%
#574795000000
1!
1%
#574800000000
0!
0%
#574805000000
1!
1%
#574810000000
0!
0%
#574815000000
1!
1%
#574820000000
0!
0%
#574825000000
1!
1%
#574830000000
0!
0%
#574835000000
1!
1%
#574840000000
0!
0%
#574845000000
1!
1%
#574850000000
0!
0%
#574855000000
1!
1%
#574860000000
0!
0%
#574865000000
1!
1%
#574870000000
0!
0%
#574875000000
1!
1%
#574880000000
0!
0%
#574885000000
1!
1%
#574890000000
0!
0%
#574895000000
1!
1%
#574900000000
0!
0%
#574905000000
1!
1%
#574910000000
0!
0%
#574915000000
1!
1%
#574920000000
0!
0%
#574925000000
1!
1%
#574930000000
0!
0%
#574935000000
1!
1%
#574940000000
0!
0%
#574945000000
1!
1%
#574950000000
0!
0%
#574955000000
1!
1%
#574960000000
0!
0%
#574965000000
1!
1%
#574970000000
0!
0%
#574975000000
1!
1%
#574980000000
0!
0%
#574985000000
1!
1%
#574990000000
0!
0%
#574995000000
1!
1%
#575000000000
0!
0%
#575005000000
1!
1%
#575010000000
0!
0%
#575015000000
1!
1%
#575020000000
0!
0%
#575025000000
1!
1%
#575030000000
0!
0%
#575035000000
1!
1%
#575040000000
0!
0%
#575045000000
1!
1%
#575050000000
0!
0%
#575055000000
1!
1%
#575060000000
0!
0%
#575065000000
1!
1%
#575070000000
0!
0%
#575075000000
1!
1%
#575080000000
0!
0%
#575085000000
1!
1%
#575090000000
0!
0%
#575095000000
1!
1%
#575100000000
0!
0%
#575105000000
1!
1%
#575110000000
0!
0%
#575115000000
1!
1%
#575120000000
0!
0%
#575125000000
1!
1%
#575130000000
0!
0%
#575135000000
1!
1%
#575140000000
0!
0%
#575145000000
1!
1%
#575150000000
0!
0%
#575155000000
1!
1%
#575160000000
0!
0%
#575165000000
1!
1%
#575170000000
0!
0%
#575175000000
1!
1%
#575180000000
0!
0%
#575185000000
1!
1%
#575190000000
0!
0%
#575195000000
1!
1%
#575200000000
0!
0%
#575205000000
1!
1%
#575210000000
0!
0%
#575215000000
1!
1%
#575220000000
0!
0%
#575225000000
1!
1%
#575230000000
0!
0%
#575235000000
1!
1%
#575240000000
0!
0%
#575245000000
1!
1%
#575250000000
0!
0%
#575255000000
1!
1%
#575260000000
0!
0%
#575265000000
1!
1%
#575270000000
0!
0%
#575275000000
1!
1%
#575280000000
0!
0%
#575285000000
1!
1%
#575290000000
0!
0%
#575295000000
1!
1%
#575300000000
0!
0%
#575305000000
1!
1%
#575310000000
0!
0%
#575315000000
1!
1%
#575320000000
0!
0%
#575325000000
1!
1%
#575330000000
0!
0%
#575335000000
1!
1%
#575340000000
0!
0%
#575345000000
1!
1%
#575350000000
0!
0%
#575355000000
1!
1%
#575360000000
0!
0%
#575365000000
1!
1%
#575370000000
0!
0%
#575375000000
1!
1%
#575380000000
0!
0%
#575385000000
1!
1%
#575390000000
0!
0%
#575395000000
1!
1%
#575400000000
0!
0%
#575405000000
1!
1%
#575410000000
0!
0%
#575415000000
1!
1%
#575420000000
0!
0%
#575425000000
1!
1%
#575430000000
0!
0%
#575435000000
1!
1%
#575440000000
0!
0%
#575445000000
1!
1%
#575450000000
0!
0%
#575455000000
1!
1%
#575460000000
0!
0%
#575465000000
1!
1%
#575470000000
0!
0%
#575475000000
1!
1%
#575480000000
0!
0%
#575485000000
1!
1%
#575490000000
0!
0%
#575495000000
1!
1%
#575500000000
0!
0%
#575505000000
1!
1%
#575510000000
0!
0%
#575515000000
1!
1%
#575520000000
0!
0%
#575525000000
1!
1%
#575530000000
0!
0%
#575535000000
1!
1%
#575540000000
0!
0%
#575545000000
1!
1%
#575550000000
0!
0%
#575555000000
1!
1%
#575560000000
0!
0%
#575565000000
1!
1%
#575570000000
0!
0%
#575575000000
1!
1%
#575580000000
0!
0%
#575585000000
1!
1%
#575590000000
0!
0%
#575595000000
1!
1%
#575600000000
0!
0%
#575605000000
1!
1%
#575610000000
0!
0%
#575615000000
1!
1%
#575620000000
0!
0%
#575625000000
1!
1%
#575630000000
0!
0%
#575635000000
1!
1%
#575640000000
0!
0%
#575645000000
1!
1%
#575650000000
0!
0%
#575655000000
1!
1%
#575660000000
0!
0%
#575665000000
1!
1%
#575670000000
0!
0%
#575675000000
1!
1%
#575680000000
0!
0%
#575685000000
1!
1%
#575690000000
0!
0%
#575695000000
1!
1%
#575700000000
0!
0%
#575705000000
1!
1%
#575710000000
0!
0%
#575715000000
1!
1%
#575720000000
0!
0%
#575725000000
1!
1%
#575730000000
0!
0%
#575735000000
1!
1%
#575740000000
0!
0%
#575745000000
1!
1%
#575750000000
0!
0%
#575755000000
1!
1%
#575760000000
0!
0%
#575765000000
1!
1%
#575770000000
0!
0%
#575775000000
1!
1%
#575780000000
0!
0%
#575785000000
1!
1%
#575790000000
0!
0%
#575795000000
1!
1%
#575800000000
0!
0%
#575805000000
1!
1%
#575810000000
0!
0%
#575815000000
1!
1%
#575820000000
0!
0%
#575825000000
1!
1%
#575830000000
0!
0%
#575835000000
1!
1%
#575840000000
0!
0%
#575845000000
1!
1%
#575850000000
0!
0%
#575855000000
1!
1%
#575860000000
0!
0%
#575865000000
1!
1%
#575870000000
0!
0%
#575875000000
1!
1%
#575880000000
0!
0%
#575885000000
1!
1%
#575890000000
0!
0%
#575895000000
1!
1%
#575900000000
0!
0%
#575905000000
1!
1%
#575910000000
0!
0%
#575915000000
1!
1%
#575920000000
0!
0%
#575925000000
1!
1%
#575930000000
0!
0%
#575935000000
1!
1%
#575940000000
0!
0%
#575945000000
1!
1%
#575950000000
0!
0%
#575955000000
1!
1%
#575960000000
0!
0%
#575965000000
1!
1%
#575970000000
0!
0%
#575975000000
1!
1%
#575980000000
0!
0%
#575985000000
1!
1%
#575990000000
0!
0%
#575995000000
1!
1%
#576000000000
0!
0%
#576005000000
1!
1%
#576010000000
0!
0%
#576015000000
1!
1%
#576020000000
0!
0%
#576025000000
1!
1%
#576030000000
0!
0%
#576035000000
1!
1%
#576040000000
0!
0%
#576045000000
1!
1%
#576050000000
0!
0%
#576055000000
1!
1%
#576060000000
0!
0%
#576065000000
1!
1%
#576070000000
0!
0%
#576075000000
1!
1%
#576080000000
0!
0%
#576085000000
1!
1%
#576090000000
0!
0%
#576095000000
1!
1%
#576100000000
0!
0%
#576105000000
1!
1%
#576110000000
0!
0%
#576115000000
1!
1%
#576120000000
0!
0%
#576125000000
1!
1%
#576130000000
0!
0%
#576135000000
1!
1%
#576140000000
0!
0%
#576145000000
1!
1%
#576150000000
0!
0%
#576155000000
1!
1%
#576160000000
0!
0%
#576165000000
1!
1%
#576170000000
0!
0%
#576175000000
1!
1%
#576180000000
0!
0%
#576185000000
1!
1%
#576190000000
0!
0%
#576195000000
1!
1%
#576200000000
0!
0%
#576205000000
1!
1%
#576210000000
0!
0%
#576215000000
1!
1%
#576220000000
0!
0%
#576225000000
1!
1%
#576230000000
0!
0%
#576235000000
1!
1%
#576240000000
0!
0%
#576245000000
1!
1%
#576250000000
0!
0%
#576255000000
1!
1%
#576260000000
0!
0%
#576265000000
1!
1%
#576270000000
0!
0%
#576275000000
1!
1%
#576280000000
0!
0%
#576285000000
1!
1%
#576290000000
0!
0%
#576295000000
1!
1%
#576300000000
0!
0%
#576305000000
1!
1%
#576310000000
0!
0%
#576315000000
1!
1%
#576320000000
0!
0%
#576325000000
1!
1%
#576330000000
0!
0%
#576335000000
1!
1%
#576340000000
0!
0%
#576345000000
1!
1%
#576350000000
0!
0%
#576355000000
1!
1%
#576360000000
0!
0%
#576365000000
1!
1%
#576370000000
0!
0%
#576375000000
1!
1%
#576380000000
0!
0%
#576385000000
1!
1%
#576390000000
0!
0%
#576395000000
1!
1%
#576400000000
0!
0%
#576405000000
1!
1%
#576410000000
0!
0%
#576415000000
1!
1%
#576420000000
0!
0%
#576425000000
1!
1%
#576430000000
0!
0%
#576435000000
1!
1%
#576440000000
0!
0%
#576445000000
1!
1%
#576450000000
0!
0%
#576455000000
1!
1%
#576460000000
0!
0%
#576465000000
1!
1%
#576470000000
0!
0%
#576475000000
1!
1%
#576480000000
0!
0%
#576485000000
1!
1%
#576490000000
0!
0%
#576495000000
1!
1%
#576500000000
0!
0%
#576505000000
1!
1%
#576510000000
0!
0%
#576515000000
1!
1%
#576520000000
0!
0%
#576525000000
1!
1%
#576530000000
0!
0%
#576535000000
1!
1%
#576540000000
0!
0%
#576545000000
1!
1%
#576550000000
0!
0%
#576555000000
1!
1%
#576560000000
0!
0%
#576565000000
1!
1%
#576570000000
0!
0%
#576575000000
1!
1%
#576580000000
0!
0%
#576585000000
1!
1%
#576590000000
0!
0%
#576595000000
1!
1%
#576600000000
0!
0%
#576605000000
1!
1%
#576610000000
0!
0%
#576615000000
1!
1%
#576620000000
0!
0%
#576625000000
1!
1%
#576630000000
0!
0%
#576635000000
1!
1%
#576640000000
0!
0%
#576645000000
1!
1%
#576650000000
0!
0%
#576655000000
1!
1%
#576660000000
0!
0%
#576665000000
1!
1%
#576670000000
0!
0%
#576675000000
1!
1%
#576680000000
0!
0%
#576685000000
1!
1%
#576690000000
0!
0%
#576695000000
1!
1%
#576700000000
0!
0%
#576705000000
1!
1%
#576710000000
0!
0%
#576715000000
1!
1%
#576720000000
0!
0%
#576725000000
1!
1%
#576730000000
0!
0%
#576735000000
1!
1%
#576740000000
0!
0%
#576745000000
1!
1%
#576750000000
0!
0%
#576755000000
1!
1%
#576760000000
0!
0%
#576765000000
1!
1%
#576770000000
0!
0%
#576775000000
1!
1%
#576780000000
0!
0%
#576785000000
1!
1%
#576790000000
0!
0%
#576795000000
1!
1%
#576800000000
0!
0%
#576805000000
1!
1%
#576810000000
0!
0%
#576815000000
1!
1%
#576820000000
0!
0%
#576825000000
1!
1%
#576830000000
0!
0%
#576835000000
1!
1%
#576840000000
0!
0%
#576845000000
1!
1%
#576850000000
0!
0%
#576855000000
1!
1%
#576860000000
0!
0%
#576865000000
1!
1%
#576870000000
0!
0%
#576875000000
1!
1%
#576880000000
0!
0%
#576885000000
1!
1%
#576890000000
0!
0%
#576895000000
1!
1%
#576900000000
0!
0%
#576905000000
1!
1%
#576910000000
0!
0%
#576915000000
1!
1%
#576920000000
0!
0%
#576925000000
1!
1%
#576930000000
0!
0%
#576935000000
1!
1%
#576940000000
0!
0%
#576945000000
1!
1%
#576950000000
0!
0%
#576955000000
1!
1%
#576960000000
0!
0%
#576965000000
1!
1%
#576970000000
0!
0%
#576975000000
1!
1%
#576980000000
0!
0%
#576985000000
1!
1%
#576990000000
0!
0%
#576995000000
1!
1%
#577000000000
0!
0%
#577005000000
1!
1%
#577010000000
0!
0%
#577015000000
1!
1%
#577020000000
0!
0%
#577025000000
1!
1%
#577030000000
0!
0%
#577035000000
1!
1%
#577040000000
0!
0%
#577045000000
1!
1%
#577050000000
0!
0%
#577055000000
1!
1%
#577060000000
0!
0%
#577065000000
1!
1%
#577070000000
0!
0%
#577075000000
1!
1%
#577080000000
0!
0%
#577085000000
1!
1%
#577090000000
0!
0%
#577095000000
1!
1%
#577100000000
0!
0%
#577105000000
1!
1%
#577110000000
0!
0%
#577115000000
1!
1%
#577120000000
0!
0%
#577125000000
1!
1%
#577130000000
0!
0%
#577135000000
1!
1%
#577140000000
0!
0%
#577145000000
1!
1%
#577150000000
0!
0%
#577155000000
1!
1%
#577160000000
0!
0%
#577165000000
1!
1%
#577170000000
0!
0%
#577175000000
1!
1%
#577180000000
0!
0%
#577185000000
1!
1%
#577190000000
0!
0%
#577195000000
1!
1%
#577200000000
0!
0%
#577205000000
1!
1%
#577210000000
0!
0%
#577215000000
1!
1%
#577220000000
0!
0%
#577225000000
1!
1%
#577230000000
0!
0%
#577235000000
1!
1%
#577240000000
0!
0%
#577245000000
1!
1%
#577250000000
0!
0%
#577255000000
1!
1%
#577260000000
0!
0%
#577265000000
1!
1%
#577270000000
0!
0%
#577275000000
1!
1%
#577280000000
0!
0%
#577285000000
1!
1%
#577290000000
0!
0%
#577295000000
1!
1%
#577300000000
0!
0%
#577305000000
1!
1%
#577310000000
0!
0%
#577315000000
1!
1%
#577320000000
0!
0%
#577325000000
1!
1%
#577330000000
0!
0%
#577335000000
1!
1%
#577340000000
0!
0%
#577345000000
1!
1%
#577350000000
0!
0%
#577355000000
1!
1%
#577360000000
0!
0%
#577365000000
1!
1%
#577370000000
0!
0%
#577375000000
1!
1%
#577380000000
0!
0%
#577385000000
1!
1%
#577390000000
0!
0%
#577395000000
1!
1%
#577400000000
0!
0%
#577405000000
1!
1%
#577410000000
0!
0%
#577415000000
1!
1%
#577420000000
0!
0%
#577425000000
1!
1%
#577430000000
0!
0%
#577435000000
1!
1%
#577440000000
0!
0%
#577445000000
1!
1%
#577450000000
0!
0%
#577455000000
1!
1%
#577460000000
0!
0%
#577465000000
1!
1%
#577470000000
0!
0%
#577475000000
1!
1%
#577480000000
0!
0%
#577485000000
1!
1%
#577490000000
0!
0%
#577495000000
1!
1%
#577500000000
0!
0%
#577505000000
1!
1%
#577510000000
0!
0%
#577515000000
1!
1%
#577520000000
0!
0%
#577525000000
1!
1%
#577530000000
0!
0%
#577535000000
1!
1%
#577540000000
0!
0%
#577545000000
1!
1%
#577550000000
0!
0%
#577555000000
1!
1%
#577560000000
0!
0%
#577565000000
1!
1%
#577570000000
0!
0%
#577575000000
1!
1%
#577580000000
0!
0%
#577585000000
1!
1%
#577590000000
0!
0%
#577595000000
1!
1%
#577600000000
0!
0%
#577605000000
1!
1%
#577610000000
0!
0%
#577615000000
1!
1%
#577620000000
0!
0%
#577625000000
1!
1%
#577630000000
0!
0%
#577635000000
1!
1%
#577640000000
0!
0%
#577645000000
1!
1%
#577650000000
0!
0%
#577655000000
1!
1%
#577660000000
0!
0%
#577665000000
1!
1%
#577670000000
0!
0%
#577675000000
1!
1%
#577680000000
0!
0%
#577685000000
1!
1%
#577690000000
0!
0%
#577695000000
1!
1%
#577700000000
0!
0%
#577705000000
1!
1%
#577710000000
0!
0%
#577715000000
1!
1%
#577720000000
0!
0%
#577725000000
1!
1%
#577730000000
0!
0%
#577735000000
1!
1%
#577740000000
0!
0%
#577745000000
1!
1%
#577750000000
0!
0%
#577755000000
1!
1%
#577760000000
0!
0%
#577765000000
1!
1%
#577770000000
0!
0%
#577775000000
1!
1%
#577780000000
0!
0%
#577785000000
1!
1%
#577790000000
0!
0%
#577795000000
1!
1%
#577800000000
0!
0%
#577805000000
1!
1%
#577810000000
0!
0%
#577815000000
1!
1%
#577820000000
0!
0%
#577825000000
1!
1%
#577830000000
0!
0%
#577835000000
1!
1%
#577840000000
0!
0%
#577845000000
1!
1%
#577850000000
0!
0%
#577855000000
1!
1%
#577860000000
0!
0%
#577865000000
1!
1%
#577870000000
0!
0%
#577875000000
1!
1%
#577880000000
0!
0%
#577885000000
1!
1%
#577890000000
0!
0%
#577895000000
1!
1%
#577900000000
0!
0%
#577905000000
1!
1%
#577910000000
0!
0%
#577915000000
1!
1%
#577920000000
0!
0%
#577925000000
1!
1%
#577930000000
0!
0%
#577935000000
1!
1%
#577940000000
0!
0%
#577945000000
1!
1%
#577950000000
0!
0%
#577955000000
1!
1%
#577960000000
0!
0%
#577965000000
1!
1%
#577970000000
0!
0%
#577975000000
1!
1%
#577980000000
0!
0%
#577985000000
1!
1%
#577990000000
0!
0%
#577995000000
1!
1%
#578000000000
0!
0%
#578005000000
1!
1%
#578010000000
0!
0%
#578015000000
1!
1%
#578020000000
0!
0%
#578025000000
1!
1%
#578030000000
0!
0%
#578035000000
1!
1%
#578040000000
0!
0%
#578045000000
1!
1%
#578050000000
0!
0%
#578055000000
1!
1%
#578060000000
0!
0%
#578065000000
1!
1%
#578070000000
0!
0%
#578075000000
1!
1%
#578080000000
0!
0%
#578085000000
1!
1%
#578090000000
0!
0%
#578095000000
1!
1%
#578100000000
0!
0%
#578105000000
1!
1%
#578110000000
0!
0%
#578115000000
1!
1%
#578120000000
0!
0%
#578125000000
1!
1%
#578130000000
0!
0%
#578135000000
1!
1%
#578140000000
0!
0%
#578145000000
1!
1%
#578150000000
0!
0%
#578155000000
1!
1%
#578160000000
0!
0%
#578165000000
1!
1%
#578170000000
0!
0%
#578175000000
1!
1%
#578180000000
0!
0%
#578185000000
1!
1%
#578190000000
0!
0%
#578195000000
1!
1%
#578200000000
0!
0%
#578205000000
1!
1%
#578210000000
0!
0%
#578215000000
1!
1%
#578220000000
0!
0%
#578225000000
1!
1%
#578230000000
0!
0%
#578235000000
1!
1%
#578240000000
0!
0%
#578245000000
1!
1%
#578250000000
0!
0%
#578255000000
1!
1%
#578260000000
0!
0%
#578265000000
1!
1%
#578270000000
0!
0%
#578275000000
1!
1%
#578280000000
0!
0%
#578285000000
1!
1%
#578290000000
0!
0%
#578295000000
1!
1%
#578300000000
0!
0%
#578305000000
1!
1%
#578310000000
0!
0%
#578315000000
1!
1%
#578320000000
0!
0%
#578325000000
1!
1%
#578330000000
0!
0%
#578335000000
1!
1%
#578340000000
0!
0%
#578345000000
1!
1%
#578350000000
0!
0%
#578355000000
1!
1%
#578360000000
0!
0%
#578365000000
1!
1%
#578370000000
0!
0%
#578375000000
1!
1%
#578380000000
0!
0%
#578385000000
1!
1%
#578390000000
0!
0%
#578395000000
1!
1%
#578400000000
0!
0%
#578405000000
1!
1%
#578410000000
0!
0%
#578415000000
1!
1%
#578420000000
0!
0%
#578425000000
1!
1%
#578430000000
0!
0%
#578435000000
1!
1%
#578440000000
0!
0%
#578445000000
1!
1%
#578450000000
0!
0%
#578455000000
1!
1%
#578460000000
0!
0%
#578465000000
1!
1%
#578470000000
0!
0%
#578475000000
1!
1%
#578480000000
0!
0%
#578485000000
1!
1%
#578490000000
0!
0%
#578495000000
1!
1%
#578500000000
0!
0%
#578505000000
1!
1%
#578510000000
0!
0%
#578515000000
1!
1%
#578520000000
0!
0%
#578525000000
1!
1%
#578530000000
0!
0%
#578535000000
1!
1%
#578540000000
0!
0%
#578545000000
1!
1%
#578550000000
0!
0%
#578555000000
1!
1%
#578560000000
0!
0%
#578565000000
1!
1%
#578570000000
0!
0%
#578575000000
1!
1%
#578580000000
0!
0%
#578585000000
1!
1%
#578590000000
0!
0%
#578595000000
1!
1%
#578600000000
0!
0%
#578605000000
1!
1%
#578610000000
0!
0%
#578615000000
1!
1%
#578620000000
0!
0%
#578625000000
1!
1%
#578630000000
0!
0%
#578635000000
1!
1%
#578640000000
0!
0%
#578645000000
1!
1%
#578650000000
0!
0%
#578655000000
1!
1%
#578660000000
0!
0%
#578665000000
1!
1%
#578670000000
0!
0%
#578675000000
1!
1%
#578680000000
0!
0%
#578685000000
1!
1%
#578690000000
0!
0%
#578695000000
1!
1%
#578700000000
0!
0%
#578705000000
1!
1%
#578710000000
0!
0%
#578715000000
1!
1%
#578720000000
0!
0%
#578725000000
1!
1%
#578730000000
0!
0%
#578735000000
1!
1%
#578740000000
0!
0%
#578745000000
1!
1%
#578750000000
0!
0%
#578755000000
1!
1%
#578760000000
0!
0%
#578765000000
1!
1%
#578770000000
0!
0%
#578775000000
1!
1%
#578780000000
0!
0%
#578785000000
1!
1%
#578790000000
0!
0%
#578795000000
1!
1%
#578800000000
0!
0%
#578805000000
1!
1%
#578810000000
0!
0%
#578815000000
1!
1%
#578820000000
0!
0%
#578825000000
1!
1%
#578830000000
0!
0%
#578835000000
1!
1%
#578840000000
0!
0%
#578845000000
1!
1%
#578850000000
0!
0%
#578855000000
1!
1%
#578860000000
0!
0%
#578865000000
1!
1%
#578870000000
0!
0%
#578875000000
1!
1%
#578880000000
0!
0%
#578885000000
1!
1%
#578890000000
0!
0%
#578895000000
1!
1%
#578900000000
0!
0%
#578905000000
1!
1%
#578910000000
0!
0%
#578915000000
1!
1%
#578920000000
0!
0%
#578925000000
1!
1%
#578930000000
0!
0%
#578935000000
1!
1%
#578940000000
0!
0%
#578945000000
1!
1%
#578950000000
0!
0%
#578955000000
1!
1%
#578960000000
0!
0%
#578965000000
1!
1%
#578970000000
0!
0%
#578975000000
1!
1%
#578980000000
0!
0%
#578985000000
1!
1%
#578990000000
0!
0%
#578995000000
1!
1%
#579000000000
0!
0%
#579005000000
1!
1%
#579010000000
0!
0%
#579015000000
1!
1%
#579020000000
0!
0%
#579025000000
1!
1%
#579030000000
0!
0%
#579035000000
1!
1%
#579040000000
0!
0%
#579045000000
1!
1%
#579050000000
0!
0%
#579055000000
1!
1%
#579060000000
0!
0%
#579065000000
1!
1%
#579070000000
0!
0%
#579075000000
1!
1%
#579080000000
0!
0%
#579085000000
1!
1%
#579090000000
0!
0%
#579095000000
1!
1%
#579100000000
0!
0%
#579105000000
1!
1%
#579110000000
0!
0%
#579115000000
1!
1%
#579120000000
0!
0%
#579125000000
1!
1%
#579130000000
0!
0%
#579135000000
1!
1%
#579140000000
0!
0%
#579145000000
1!
1%
#579150000000
0!
0%
#579155000000
1!
1%
#579160000000
0!
0%
#579165000000
1!
1%
#579170000000
0!
0%
#579175000000
1!
1%
#579180000000
0!
0%
#579185000000
1!
1%
#579190000000
0!
0%
#579195000000
1!
1%
#579200000000
0!
0%
#579205000000
1!
1%
#579210000000
0!
0%
#579215000000
1!
1%
#579220000000
0!
0%
#579225000000
1!
1%
#579230000000
0!
0%
#579235000000
1!
1%
#579240000000
0!
0%
#579245000000
1!
1%
#579250000000
0!
0%
#579255000000
1!
1%
#579260000000
0!
0%
#579265000000
1!
1%
#579270000000
0!
0%
#579275000000
1!
1%
#579280000000
0!
0%
#579285000000
1!
1%
#579290000000
0!
0%
#579295000000
1!
1%
#579300000000
0!
0%
#579305000000
1!
1%
#579310000000
0!
0%
#579315000000
1!
1%
#579320000000
0!
0%
#579325000000
1!
1%
#579330000000
0!
0%
#579335000000
1!
1%
#579340000000
0!
0%
#579345000000
1!
1%
#579350000000
0!
0%
#579355000000
1!
1%
#579360000000
0!
0%
#579365000000
1!
1%
#579370000000
0!
0%
#579375000000
1!
1%
#579380000000
0!
0%
#579385000000
1!
1%
#579390000000
0!
0%
#579395000000
1!
1%
#579400000000
0!
0%
#579405000000
1!
1%
#579410000000
0!
0%
#579415000000
1!
1%
#579420000000
0!
0%
#579425000000
1!
1%
#579430000000
0!
0%
#579435000000
1!
1%
#579440000000
0!
0%
#579445000000
1!
1%
#579450000000
0!
0%
#579455000000
1!
1%
#579460000000
0!
0%
#579465000000
1!
1%
#579470000000
0!
0%
#579475000000
1!
1%
#579480000000
0!
0%
#579485000000
1!
1%
#579490000000
0!
0%
#579495000000
1!
1%
#579500000000
0!
0%
#579505000000
1!
1%
#579510000000
0!
0%
#579515000000
1!
1%
#579520000000
0!
0%
#579525000000
1!
1%
#579530000000
0!
0%
#579535000000
1!
1%
#579540000000
0!
0%
#579545000000
1!
1%
#579550000000
0!
0%
#579555000000
1!
1%
#579560000000
0!
0%
#579565000000
1!
1%
#579570000000
0!
0%
#579575000000
1!
1%
#579580000000
0!
0%
#579585000000
1!
1%
#579590000000
0!
0%
#579595000000
1!
1%
#579600000000
0!
0%
#579605000000
1!
1%
#579610000000
0!
0%
#579615000000
1!
1%
#579620000000
0!
0%
#579625000000
1!
1%
#579630000000
0!
0%
#579635000000
1!
1%
#579640000000
0!
0%
#579645000000
1!
1%
#579650000000
0!
0%
#579655000000
1!
1%
#579660000000
0!
0%
#579665000000
1!
1%
#579670000000
0!
0%
#579675000000
1!
1%
#579680000000
0!
0%
#579685000000
1!
1%
#579690000000
0!
0%
#579695000000
1!
1%
#579700000000
0!
0%
#579705000000
1!
1%
#579710000000
0!
0%
#579715000000
1!
1%
#579720000000
0!
0%
#579725000000
1!
1%
#579730000000
0!
0%
#579735000000
1!
1%
#579740000000
0!
0%
#579745000000
1!
1%
#579750000000
0!
0%
#579755000000
1!
1%
#579760000000
0!
0%
#579765000000
1!
1%
#579770000000
0!
0%
#579775000000
1!
1%
#579780000000
0!
0%
#579785000000
1!
1%
#579790000000
0!
0%
#579795000000
1!
1%
#579800000000
0!
0%
#579805000000
1!
1%
#579810000000
0!
0%
#579815000000
1!
1%
#579820000000
0!
0%
#579825000000
1!
1%
#579830000000
0!
0%
#579835000000
1!
1%
#579840000000
0!
0%
#579845000000
1!
1%
#579850000000
0!
0%
#579855000000
1!
1%
#579860000000
0!
0%
#579865000000
1!
1%
#579870000000
0!
0%
#579875000000
1!
1%
#579880000000
0!
0%
#579885000000
1!
1%
#579890000000
0!
0%
#579895000000
1!
1%
#579900000000
0!
0%
#579905000000
1!
1%
#579910000000
0!
0%
#579915000000
1!
1%
#579920000000
0!
0%
#579925000000
1!
1%
#579930000000
0!
0%
#579935000000
1!
1%
#579940000000
0!
0%
#579945000000
1!
1%
#579950000000
0!
0%
#579955000000
1!
1%
#579960000000
0!
0%
#579965000000
1!
1%
#579970000000
0!
0%
#579975000000
1!
1%
#579980000000
0!
0%
#579985000000
1!
1%
#579990000000
0!
0%
#579995000000
1!
1%
#580000000000
0!
0%
#580005000000
1!
1%
#580010000000
0!
0%
#580015000000
1!
1%
#580020000000
0!
0%
#580025000000
1!
1%
#580030000000
0!
0%
#580035000000
1!
1%
#580040000000
0!
0%
#580045000000
1!
1%
#580050000000
0!
0%
#580055000000
1!
1%
#580060000000
0!
0%
#580065000000
1!
1%
#580070000000
0!
0%
#580075000000
1!
1%
#580080000000
0!
0%
#580085000000
1!
1%
#580090000000
0!
0%
#580095000000
1!
1%
#580100000000
0!
0%
#580105000000
1!
1%
#580110000000
0!
0%
#580115000000
1!
1%
#580120000000
0!
0%
#580125000000
1!
1%
#580130000000
0!
0%
#580135000000
1!
1%
#580140000000
0!
0%
#580145000000
1!
1%
#580150000000
0!
0%
#580155000000
1!
1%
#580160000000
0!
0%
#580165000000
1!
1%
#580170000000
0!
0%
#580175000000
1!
1%
#580180000000
0!
0%
#580185000000
1!
1%
#580190000000
0!
0%
#580195000000
1!
1%
#580200000000
0!
0%
#580205000000
1!
1%
#580210000000
0!
0%
#580215000000
1!
1%
#580220000000
0!
0%
#580225000000
1!
1%
#580230000000
0!
0%
#580235000000
1!
1%
#580240000000
0!
0%
#580245000000
1!
1%
#580250000000
0!
0%
#580255000000
1!
1%
#580260000000
0!
0%
#580265000000
1!
1%
#580270000000
0!
0%
#580275000000
1!
1%
#580280000000
0!
0%
#580285000000
1!
1%
#580290000000
0!
0%
#580295000000
1!
1%
#580300000000
0!
0%
#580305000000
1!
1%
#580310000000
0!
0%
#580315000000
1!
1%
#580320000000
0!
0%
#580325000000
1!
1%
#580330000000
0!
0%
#580335000000
1!
1%
#580340000000
0!
0%
#580345000000
1!
1%
#580350000000
0!
0%
#580355000000
1!
1%
#580360000000
0!
0%
#580365000000
1!
1%
#580370000000
0!
0%
#580375000000
1!
1%
#580380000000
0!
0%
#580385000000
1!
1%
#580390000000
0!
0%
#580395000000
1!
1%
#580400000000
0!
0%
#580405000000
1!
1%
#580410000000
0!
0%
#580415000000
1!
1%
#580420000000
0!
0%
#580425000000
1!
1%
#580430000000
0!
0%
#580435000000
1!
1%
#580440000000
0!
0%
#580445000000
1!
1%
#580450000000
0!
0%
#580455000000
1!
1%
#580460000000
0!
0%
#580465000000
1!
1%
#580470000000
0!
0%
#580475000000
1!
1%
#580480000000
0!
0%
#580485000000
1!
1%
#580490000000
0!
0%
#580495000000
1!
1%
#580500000000
0!
0%
#580505000000
1!
1%
#580510000000
0!
0%
#580515000000
1!
1%
#580520000000
0!
0%
#580525000000
1!
1%
#580530000000
0!
0%
#580535000000
1!
1%
#580540000000
0!
0%
#580545000000
1!
1%
#580550000000
0!
0%
#580555000000
1!
1%
#580560000000
0!
0%
#580565000000
1!
1%
#580570000000
0!
0%
#580575000000
1!
1%
#580580000000
0!
0%
#580585000000
1!
1%
#580590000000
0!
0%
#580595000000
1!
1%
#580600000000
0!
0%
#580605000000
1!
1%
#580610000000
0!
0%
#580615000000
1!
1%
#580620000000
0!
0%
#580625000000
1!
1%
#580630000000
0!
0%
#580635000000
1!
1%
#580640000000
0!
0%
#580645000000
1!
1%
#580650000000
0!
0%
#580655000000
1!
1%
#580660000000
0!
0%
#580665000000
1!
1%
#580670000000
0!
0%
#580675000000
1!
1%
#580680000000
0!
0%
#580685000000
1!
1%
#580690000000
0!
0%
#580695000000
1!
1%
#580700000000
0!
0%
#580705000000
1!
1%
#580710000000
0!
0%
#580715000000
1!
1%
#580720000000
0!
0%
#580725000000
1!
1%
#580730000000
0!
0%
#580735000000
1!
1%
#580740000000
0!
0%
#580745000000
1!
1%
#580750000000
0!
0%
#580755000000
1!
1%
#580760000000
0!
0%
#580765000000
1!
1%
#580770000000
0!
0%
#580775000000
1!
1%
#580780000000
0!
0%
#580785000000
1!
1%
#580790000000
0!
0%
#580795000000
1!
1%
#580800000000
0!
0%
#580805000000
1!
1%
#580810000000
0!
0%
#580815000000
1!
1%
#580820000000
0!
0%
#580825000000
1!
1%
#580830000000
0!
0%
#580835000000
1!
1%
#580840000000
0!
0%
#580845000000
1!
1%
#580850000000
0!
0%
#580855000000
1!
1%
#580860000000
0!
0%
#580865000000
1!
1%
#580870000000
0!
0%
#580875000000
1!
1%
#580880000000
0!
0%
#580885000000
1!
1%
#580890000000
0!
0%
#580895000000
1!
1%
#580900000000
0!
0%
#580905000000
1!
1%
#580910000000
0!
0%
#580915000000
1!
1%
#580920000000
0!
0%
#580925000000
1!
1%
#580930000000
0!
0%
#580935000000
1!
1%
#580940000000
0!
0%
#580945000000
1!
1%
#580950000000
0!
0%
#580955000000
1!
1%
#580960000000
0!
0%
#580965000000
1!
1%
#580970000000
0!
0%
#580975000000
1!
1%
#580980000000
0!
0%
#580985000000
1!
1%
#580990000000
0!
0%
#580995000000
1!
1%
#581000000000
0!
0%
#581005000000
1!
1%
#581010000000
0!
0%
#581015000000
1!
1%
#581020000000
0!
0%
#581025000000
1!
1%
#581030000000
0!
0%
#581035000000
1!
1%
#581040000000
0!
0%
#581045000000
1!
1%
#581050000000
0!
0%
#581055000000
1!
1%
#581060000000
0!
0%
#581065000000
1!
1%
#581070000000
0!
0%
#581075000000
1!
1%
#581080000000
0!
0%
#581085000000
1!
1%
#581090000000
0!
0%
#581095000000
1!
1%
#581100000000
0!
0%
#581105000000
1!
1%
#581110000000
0!
0%
#581115000000
1!
1%
#581120000000
0!
0%
#581125000000
1!
1%
#581130000000
0!
0%
#581135000000
1!
1%
#581140000000
0!
0%
#581145000000
1!
1%
#581150000000
0!
0%
#581155000000
1!
1%
#581160000000
0!
0%
#581165000000
1!
1%
#581170000000
0!
0%
#581175000000
1!
1%
#581180000000
0!
0%
#581185000000
1!
1%
#581190000000
0!
0%
#581195000000
1!
1%
#581200000000
0!
0%
#581205000000
1!
1%
#581210000000
0!
0%
#581215000000
1!
1%
#581220000000
0!
0%
#581225000000
1!
1%
#581230000000
0!
0%
#581235000000
1!
1%
#581240000000
0!
0%
#581245000000
1!
1%
#581250000000
0!
0%
#581255000000
1!
1%
#581260000000
0!
0%
#581265000000
1!
1%
#581270000000
0!
0%
#581275000000
1!
1%
#581280000000
0!
0%
#581285000000
1!
1%
#581290000000
0!
0%
#581295000000
1!
1%
#581300000000
0!
0%
#581305000000
1!
1%
#581310000000
0!
0%
#581315000000
1!
1%
#581320000000
0!
0%
#581325000000
1!
1%
#581330000000
0!
0%
#581335000000
1!
1%
#581340000000
0!
0%
#581345000000
1!
1%
#581350000000
0!
0%
#581355000000
1!
1%
#581360000000
0!
0%
#581365000000
1!
1%
#581370000000
0!
0%
#581375000000
1!
1%
#581380000000
0!
0%
#581385000000
1!
1%
#581390000000
0!
0%
#581395000000
1!
1%
#581400000000
0!
0%
#581405000000
1!
1%
#581410000000
0!
0%
#581415000000
1!
1%
#581420000000
0!
0%
#581425000000
1!
1%
#581430000000
0!
0%
#581435000000
1!
1%
#581440000000
0!
0%
#581445000000
1!
1%
#581450000000
0!
0%
#581455000000
1!
1%
#581460000000
0!
0%
#581465000000
1!
1%
#581470000000
0!
0%
#581475000000
1!
1%
#581480000000
0!
0%
#581485000000
1!
1%
#581490000000
0!
0%
#581495000000
1!
1%
#581500000000
0!
0%
#581505000000
1!
1%
#581510000000
0!
0%
#581515000000
1!
1%
#581520000000
0!
0%
#581525000000
1!
1%
#581530000000
0!
0%
#581535000000
1!
1%
#581540000000
0!
0%
#581545000000
1!
1%
#581550000000
0!
0%
#581555000000
1!
1%
#581560000000
0!
0%
#581565000000
1!
1%
#581570000000
0!
0%
#581575000000
1!
1%
#581580000000
0!
0%
#581585000000
1!
1%
#581590000000
0!
0%
#581595000000
1!
1%
#581600000000
0!
0%
#581605000000
1!
1%
#581610000000
0!
0%
#581615000000
1!
1%
#581620000000
0!
0%
#581625000000
1!
1%
#581630000000
0!
0%
#581635000000
1!
1%
#581640000000
0!
0%
#581645000000
1!
1%
#581650000000
0!
0%
#581655000000
1!
1%
#581660000000
0!
0%
#581665000000
1!
1%
#581670000000
0!
0%
#581675000000
1!
1%
#581680000000
0!
0%
#581685000000
1!
1%
#581690000000
0!
0%
#581695000000
1!
1%
#581700000000
0!
0%
#581705000000
1!
1%
#581710000000
0!
0%
#581715000000
1!
1%
#581720000000
0!
0%
#581725000000
1!
1%
#581730000000
0!
0%
#581735000000
1!
1%
#581740000000
0!
0%
#581745000000
1!
1%
#581750000000
0!
0%
#581755000000
1!
1%
#581760000000
0!
0%
#581765000000
1!
1%
#581770000000
0!
0%
#581775000000
1!
1%
#581780000000
0!
0%
#581785000000
1!
1%
#581790000000
0!
0%
#581795000000
1!
1%
#581800000000
0!
0%
#581805000000
1!
1%
#581810000000
0!
0%
#581815000000
1!
1%
#581820000000
0!
0%
#581825000000
1!
1%
#581830000000
0!
0%
#581835000000
1!
1%
#581840000000
0!
0%
#581845000000
1!
1%
#581850000000
0!
0%
#581855000000
1!
1%
#581860000000
0!
0%
#581865000000
1!
1%
#581870000000
0!
0%
#581875000000
1!
1%
#581880000000
0!
0%
#581885000000
1!
1%
#581890000000
0!
0%
#581895000000
1!
1%
#581900000000
0!
0%
#581905000000
1!
1%
#581910000000
0!
0%
#581915000000
1!
1%
#581920000000
0!
0%
#581925000000
1!
1%
#581930000000
0!
0%
#581935000000
1!
1%
#581940000000
0!
0%
#581945000000
1!
1%
#581950000000
0!
0%
#581955000000
1!
1%
#581960000000
0!
0%
#581965000000
1!
1%
#581970000000
0!
0%
#581975000000
1!
1%
#581980000000
0!
0%
#581985000000
1!
1%
#581990000000
0!
0%
#581995000000
1!
1%
#582000000000
0!
0%
#582005000000
1!
1%
#582010000000
0!
0%
#582015000000
1!
1%
#582020000000
0!
0%
#582025000000
1!
1%
#582030000000
0!
0%
#582035000000
1!
1%
#582040000000
0!
0%
#582045000000
1!
1%
#582050000000
0!
0%
#582055000000
1!
1%
#582060000000
0!
0%
#582065000000
1!
1%
#582070000000
0!
0%
#582075000000
1!
1%
#582080000000
0!
0%
#582085000000
1!
1%
#582090000000
0!
0%
#582095000000
1!
1%
#582100000000
0!
0%
#582105000000
1!
1%
#582110000000
0!
0%
#582115000000
1!
1%
#582120000000
0!
0%
#582125000000
1!
1%
#582130000000
0!
0%
#582135000000
1!
1%
#582140000000
0!
0%
#582145000000
1!
1%
#582150000000
0!
0%
#582155000000
1!
1%
#582160000000
0!
0%
#582165000000
1!
1%
#582170000000
0!
0%
#582175000000
1!
1%
#582180000000
0!
0%
#582185000000
1!
1%
#582190000000
0!
0%
#582195000000
1!
1%
#582200000000
0!
0%
#582205000000
1!
1%
#582210000000
0!
0%
#582215000000
1!
1%
#582220000000
0!
0%
#582225000000
1!
1%
#582230000000
0!
0%
#582235000000
1!
1%
#582240000000
0!
0%
#582245000000
1!
1%
#582250000000
0!
0%
#582255000000
1!
1%
#582260000000
0!
0%
#582265000000
1!
1%
#582270000000
0!
0%
#582275000000
1!
1%
#582280000000
0!
0%
#582285000000
1!
1%
#582290000000
0!
0%
#582295000000
1!
1%
#582300000000
0!
0%
#582305000000
1!
1%
#582310000000
0!
0%
#582315000000
1!
1%
#582320000000
0!
0%
#582325000000
1!
1%
#582330000000
0!
0%
#582335000000
1!
1%
#582340000000
0!
0%
#582345000000
1!
1%
#582350000000
0!
0%
#582355000000
1!
1%
#582360000000
0!
0%
#582365000000
1!
1%
#582370000000
0!
0%
#582375000000
1!
1%
#582380000000
0!
0%
#582385000000
1!
1%
#582390000000
0!
0%
#582395000000
1!
1%
#582400000000
0!
0%
#582405000000
1!
1%
#582410000000
0!
0%
#582415000000
1!
1%
#582420000000
0!
0%
#582425000000
1!
1%
#582430000000
0!
0%
#582435000000
1!
1%
#582440000000
0!
0%
#582445000000
1!
1%
#582450000000
0!
0%
#582455000000
1!
1%
#582460000000
0!
0%
#582465000000
1!
1%
#582470000000
0!
0%
#582475000000
1!
1%
#582480000000
0!
0%
#582485000000
1!
1%
#582490000000
0!
0%
#582495000000
1!
1%
#582500000000
0!
0%
#582505000000
1!
1%
#582510000000
0!
0%
#582515000000
1!
1%
#582520000000
0!
0%
#582525000000
1!
1%
#582530000000
0!
0%
#582535000000
1!
1%
#582540000000
0!
0%
#582545000000
1!
1%
#582550000000
0!
0%
#582555000000
1!
1%
#582560000000
0!
0%
#582565000000
1!
1%
#582570000000
0!
0%
#582575000000
1!
1%
#582580000000
0!
0%
#582585000000
1!
1%
#582590000000
0!
0%
#582595000000
1!
1%
#582600000000
0!
0%
#582605000000
1!
1%
#582610000000
0!
0%
#582615000000
1!
1%
#582620000000
0!
0%
#582625000000
1!
1%
#582630000000
0!
0%
#582635000000
1!
1%
#582640000000
0!
0%
#582645000000
1!
1%
#582650000000
0!
0%
#582655000000
1!
1%
#582660000000
0!
0%
#582665000000
1!
1%
#582670000000
0!
0%
#582675000000
1!
1%
#582680000000
0!
0%
#582685000000
1!
1%
#582690000000
0!
0%
#582695000000
1!
1%
#582700000000
0!
0%
#582705000000
1!
1%
#582710000000
0!
0%
#582715000000
1!
1%
#582720000000
0!
0%
#582725000000
1!
1%
#582730000000
0!
0%
#582735000000
1!
1%
#582740000000
0!
0%
#582745000000
1!
1%
#582750000000
0!
0%
#582755000000
1!
1%
#582760000000
0!
0%
#582765000000
1!
1%
#582770000000
0!
0%
#582775000000
1!
1%
#582780000000
0!
0%
#582785000000
1!
1%
#582790000000
0!
0%
#582795000000
1!
1%
#582800000000
0!
0%
#582805000000
1!
1%
#582810000000
0!
0%
#582815000000
1!
1%
#582820000000
0!
0%
#582825000000
1!
1%
#582830000000
0!
0%
#582835000000
1!
1%
#582840000000
0!
0%
#582845000000
1!
1%
#582850000000
0!
0%
#582855000000
1!
1%
#582860000000
0!
0%
#582865000000
1!
1%
#582870000000
0!
0%
#582875000000
1!
1%
#582880000000
0!
0%
#582885000000
1!
1%
#582890000000
0!
0%
#582895000000
1!
1%
#582900000000
0!
0%
#582905000000
1!
1%
#582910000000
0!
0%
#582915000000
1!
1%
#582920000000
0!
0%
#582925000000
1!
1%
#582930000000
0!
0%
#582935000000
1!
1%
#582940000000
0!
0%
#582945000000
1!
1%
#582950000000
0!
0%
#582955000000
1!
1%
#582960000000
0!
0%
#582965000000
1!
1%
#582970000000
0!
0%
#582975000000
1!
1%
#582980000000
0!
0%
#582985000000
1!
1%
#582990000000
0!
0%
#582995000000
1!
1%
#583000000000
0!
0%
#583005000000
1!
1%
#583010000000
0!
0%
#583015000000
1!
1%
#583020000000
0!
0%
#583025000000
1!
1%
#583030000000
0!
0%
#583035000000
1!
1%
#583040000000
0!
0%
#583045000000
1!
1%
#583050000000
0!
0%
#583055000000
1!
1%
#583060000000
0!
0%
#583065000000
1!
1%
#583070000000
0!
0%
#583075000000
1!
1%
#583080000000
0!
0%
#583085000000
1!
1%
#583090000000
0!
0%
#583095000000
1!
1%
#583100000000
0!
0%
#583105000000
1!
1%
#583110000000
0!
0%
#583115000000
1!
1%
#583120000000
0!
0%
#583125000000
1!
1%
#583130000000
0!
0%
#583135000000
1!
1%
#583140000000
0!
0%
#583145000000
1!
1%
#583150000000
0!
0%
#583155000000
1!
1%
#583160000000
0!
0%
#583165000000
1!
1%
#583170000000
0!
0%
#583175000000
1!
1%
#583180000000
0!
0%
#583185000000
1!
1%
#583190000000
0!
0%
#583195000000
1!
1%
#583200000000
0!
0%
#583205000000
1!
1%
#583210000000
0!
0%
#583215000000
1!
1%
#583220000000
0!
0%
#583225000000
1!
1%
#583230000000
0!
0%
#583235000000
1!
1%
#583240000000
0!
0%
#583245000000
1!
1%
#583250000000
0!
0%
#583255000000
1!
1%
#583260000000
0!
0%
#583265000000
1!
1%
#583270000000
0!
0%
#583275000000
1!
1%
#583280000000
0!
0%
#583285000000
1!
1%
#583290000000
0!
0%
#583295000000
1!
1%
#583300000000
0!
0%
#583305000000
1!
1%
#583310000000
0!
0%
#583315000000
1!
1%
#583320000000
0!
0%
#583325000000
1!
1%
#583330000000
0!
0%
#583335000000
1!
1%
#583340000000
0!
0%
#583345000000
1!
1%
#583350000000
0!
0%
#583355000000
1!
1%
#583360000000
0!
0%
#583365000000
1!
1%
#583370000000
0!
0%
#583375000000
1!
1%
#583380000000
0!
0%
#583385000000
1!
1%
#583390000000
0!
0%
#583395000000
1!
1%
#583400000000
0!
0%
#583405000000
1!
1%
#583410000000
0!
0%
#583415000000
1!
1%
#583420000000
0!
0%
#583425000000
1!
1%
#583430000000
0!
0%
#583435000000
1!
1%
#583440000000
0!
0%
#583445000000
1!
1%
#583450000000
0!
0%
#583455000000
1!
1%
#583460000000
0!
0%
#583465000000
1!
1%
#583470000000
0!
0%
#583475000000
1!
1%
#583480000000
0!
0%
#583485000000
1!
1%
#583490000000
0!
0%
#583495000000
1!
1%
#583500000000
0!
0%
#583505000000
1!
1%
#583510000000
0!
0%
#583515000000
1!
1%
#583520000000
0!
0%
#583525000000
1!
1%
#583530000000
0!
0%
#583535000000
1!
1%
#583540000000
0!
0%
#583545000000
1!
1%
#583550000000
0!
0%
#583555000000
1!
1%
#583560000000
0!
0%
#583565000000
1!
1%
#583570000000
0!
0%
#583575000000
1!
1%
#583580000000
0!
0%
#583585000000
1!
1%
#583590000000
0!
0%
#583595000000
1!
1%
#583600000000
0!
0%
#583605000000
1!
1%
#583610000000
0!
0%
#583615000000
1!
1%
#583620000000
0!
0%
#583625000000
1!
1%
#583630000000
0!
0%
#583635000000
1!
1%
#583640000000
0!
0%
#583645000000
1!
1%
#583650000000
0!
0%
#583655000000
1!
1%
#583660000000
0!
0%
#583665000000
1!
1%
#583670000000
0!
0%
#583675000000
1!
1%
#583680000000
0!
0%
#583685000000
1!
1%
#583690000000
0!
0%
#583695000000
1!
1%
#583700000000
0!
0%
#583705000000
1!
1%
#583710000000
0!
0%
#583715000000
1!
1%
#583720000000
0!
0%
#583725000000
1!
1%
#583730000000
0!
0%
#583735000000
1!
1%
#583740000000
0!
0%
#583745000000
1!
1%
#583750000000
0!
0%
#583755000000
1!
1%
#583760000000
0!
0%
#583765000000
1!
1%
#583770000000
0!
0%
#583775000000
1!
1%
#583780000000
0!
0%
#583785000000
1!
1%
#583790000000
0!
0%
#583795000000
1!
1%
#583800000000
0!
0%
#583805000000
1!
1%
#583810000000
0!
0%
#583815000000
1!
1%
#583820000000
0!
0%
#583825000000
1!
1%
#583830000000
0!
0%
#583835000000
1!
1%
#583840000000
0!
0%
#583845000000
1!
1%
#583850000000
0!
0%
#583855000000
1!
1%
#583860000000
0!
0%
#583865000000
1!
1%
#583870000000
0!
0%
#583875000000
1!
1%
#583880000000
0!
0%
#583885000000
1!
1%
#583890000000
0!
0%
#583895000000
1!
1%
#583900000000
0!
0%
#583905000000
1!
1%
#583910000000
0!
0%
#583915000000
1!
1%
#583920000000
0!
0%
#583925000000
1!
1%
#583930000000
0!
0%
#583935000000
1!
1%
#583940000000
0!
0%
#583945000000
1!
1%
#583950000000
0!
0%
#583955000000
1!
1%
#583960000000
0!
0%
#583965000000
1!
1%
#583970000000
0!
0%
#583975000000
1!
1%
#583980000000
0!
0%
#583985000000
1!
1%
#583990000000
0!
0%
#583995000000
1!
1%
#584000000000
0!
0%
#584005000000
1!
1%
#584010000000
0!
0%
#584015000000
1!
1%
#584020000000
0!
0%
#584025000000
1!
1%
#584030000000
0!
0%
#584035000000
1!
1%
#584040000000
0!
0%
#584045000000
1!
1%
#584050000000
0!
0%
#584055000000
1!
1%
#584060000000
0!
0%
#584065000000
1!
1%
#584070000000
0!
0%
#584075000000
1!
1%
#584080000000
0!
0%
#584085000000
1!
1%
#584090000000
0!
0%
#584095000000
1!
1%
#584100000000
0!
0%
#584105000000
1!
1%
#584110000000
0!
0%
#584115000000
1!
1%
#584120000000
0!
0%
#584125000000
1!
1%
#584130000000
0!
0%
#584135000000
1!
1%
#584140000000
0!
0%
#584145000000
1!
1%
#584150000000
0!
0%
#584155000000
1!
1%
#584160000000
0!
0%
#584165000000
1!
1%
#584170000000
0!
0%
#584175000000
1!
1%
#584180000000
0!
0%
#584185000000
1!
1%
#584190000000
0!
0%
#584195000000
1!
1%
#584200000000
0!
0%
#584205000000
1!
1%
#584210000000
0!
0%
#584215000000
1!
1%
#584220000000
0!
0%
#584225000000
1!
1%
#584230000000
0!
0%
#584235000000
1!
1%
#584240000000
0!
0%
#584245000000
1!
1%
#584250000000
0!
0%
#584255000000
1!
1%
#584260000000
0!
0%
#584265000000
1!
1%
#584270000000
0!
0%
#584275000000
1!
1%
#584280000000
0!
0%
#584285000000
1!
1%
#584290000000
0!
0%
#584295000000
1!
1%
#584300000000
0!
0%
#584305000000
1!
1%
#584310000000
0!
0%
#584315000000
1!
1%
#584320000000
0!
0%
#584325000000
1!
1%
#584330000000
0!
0%
#584335000000
1!
1%
#584340000000
0!
0%
#584345000000
1!
1%
#584350000000
0!
0%
#584355000000
1!
1%
#584360000000
0!
0%
#584365000000
1!
1%
#584370000000
0!
0%
#584375000000
1!
1%
#584380000000
0!
0%
#584385000000
1!
1%
#584390000000
0!
0%
#584395000000
1!
1%
#584400000000
0!
0%
#584405000000
1!
1%
#584410000000
0!
0%
#584415000000
1!
1%
#584420000000
0!
0%
#584425000000
1!
1%
#584430000000
0!
0%
#584435000000
1!
1%
#584440000000
0!
0%
#584445000000
1!
1%
#584450000000
0!
0%
#584455000000
1!
1%
#584460000000
0!
0%
#584465000000
1!
1%
#584470000000
0!
0%
#584475000000
1!
1%
#584480000000
0!
0%
#584485000000
1!
1%
#584490000000
0!
0%
#584495000000
1!
1%
#584500000000
0!
0%
#584505000000
1!
1%
#584510000000
0!
0%
#584515000000
1!
1%
#584520000000
0!
0%
#584525000000
1!
1%
#584530000000
0!
0%
#584535000000
1!
1%
#584540000000
0!
0%
#584545000000
1!
1%
#584550000000
0!
0%
#584555000000
1!
1%
#584560000000
0!
0%
#584565000000
1!
1%
#584570000000
0!
0%
#584575000000
1!
1%
#584580000000
0!
0%
#584585000000
1!
1%
#584590000000
0!
0%
#584595000000
1!
1%
#584600000000
0!
0%
#584605000000
1!
1%
#584610000000
0!
0%
#584615000000
1!
1%
#584620000000
0!
0%
#584625000000
1!
1%
#584630000000
0!
0%
#584635000000
1!
1%
#584640000000
0!
0%
#584645000000
1!
1%
#584650000000
0!
0%
#584655000000
1!
1%
#584660000000
0!
0%
#584665000000
1!
1%
#584670000000
0!
0%
#584675000000
1!
1%
#584680000000
0!
0%
#584685000000
1!
1%
#584690000000
0!
0%
#584695000000
1!
1%
#584700000000
0!
0%
#584705000000
1!
1%
#584710000000
0!
0%
#584715000000
1!
1%
#584720000000
0!
0%
#584725000000
1!
1%
#584730000000
0!
0%
#584735000000
1!
1%
#584740000000
0!
0%
#584745000000
1!
1%
#584750000000
0!
0%
#584755000000
1!
1%
#584760000000
0!
0%
#584765000000
1!
1%
#584770000000
0!
0%
#584775000000
1!
1%
#584780000000
0!
0%
#584785000000
1!
1%
#584790000000
0!
0%
#584795000000
1!
1%
#584800000000
0!
0%
#584805000000
1!
1%
#584810000000
0!
0%
#584815000000
1!
1%
#584820000000
0!
0%
#584825000000
1!
1%
#584830000000
0!
0%
#584835000000
1!
1%
#584840000000
0!
0%
#584845000000
1!
1%
#584850000000
0!
0%
#584855000000
1!
1%
#584860000000
0!
0%
#584865000000
1!
1%
#584870000000
0!
0%
#584875000000
1!
1%
#584880000000
0!
0%
#584885000000
1!
1%
#584890000000
0!
0%
#584895000000
1!
1%
#584900000000
0!
0%
#584905000000
1!
1%
#584910000000
0!
0%
#584915000000
1!
1%
#584920000000
0!
0%
#584925000000
1!
1%
#584930000000
0!
0%
#584935000000
1!
1%
#584940000000
0!
0%
#584945000000
1!
1%
#584950000000
0!
0%
#584955000000
1!
1%
#584960000000
0!
0%
#584965000000
1!
1%
#584970000000
0!
0%
#584975000000
1!
1%
#584980000000
0!
0%
#584985000000
1!
1%
#584990000000
0!
0%
#584995000000
1!
1%
#585000000000
0!
0%
#585005000000
1!
1%
#585010000000
0!
0%
#585015000000
1!
1%
#585020000000
0!
0%
#585025000000
1!
1%
#585030000000
0!
0%
#585035000000
1!
1%
#585040000000
0!
0%
#585045000000
1!
1%
#585050000000
0!
0%
#585055000000
1!
1%
#585060000000
0!
0%
#585065000000
1!
1%
#585070000000
0!
0%
#585075000000
1!
1%
#585080000000
0!
0%
#585085000000
1!
1%
#585090000000
0!
0%
#585095000000
1!
1%
#585100000000
0!
0%
#585105000000
1!
1%
#585110000000
0!
0%
#585115000000
1!
1%
#585120000000
0!
0%
#585125000000
1!
1%
#585130000000
0!
0%
#585135000000
1!
1%
#585140000000
0!
0%
#585145000000
1!
1%
#585150000000
0!
0%
#585155000000
1!
1%
#585160000000
0!
0%
#585165000000
1!
1%
#585170000000
0!
0%
#585175000000
1!
1%
#585180000000
0!
0%
#585185000000
1!
1%
#585190000000
0!
0%
#585195000000
1!
1%
#585200000000
0!
0%
#585205000000
1!
1%
#585210000000
0!
0%
#585215000000
1!
1%
#585220000000
0!
0%
#585225000000
1!
1%
#585230000000
0!
0%
#585235000000
1!
1%
#585240000000
0!
0%
#585245000000
1!
1%
#585250000000
0!
0%
#585255000000
1!
1%
#585260000000
0!
0%
#585265000000
1!
1%
#585270000000
0!
0%
#585275000000
1!
1%
#585280000000
0!
0%
#585285000000
1!
1%
#585290000000
0!
0%
#585295000000
1!
1%
#585300000000
0!
0%
#585305000000
1!
1%
#585310000000
0!
0%
#585315000000
1!
1%
#585320000000
0!
0%
#585325000000
1!
1%
#585330000000
0!
0%
#585335000000
1!
1%
#585340000000
0!
0%
#585345000000
1!
1%
#585350000000
0!
0%
#585355000000
1!
1%
#585360000000
0!
0%
#585365000000
1!
1%
#585370000000
0!
0%
#585375000000
1!
1%
#585380000000
0!
0%
#585385000000
1!
1%
#585390000000
0!
0%
#585395000000
1!
1%
#585400000000
0!
0%
#585405000000
1!
1%
#585410000000
0!
0%
#585415000000
1!
1%
#585420000000
0!
0%
#585425000000
1!
1%
#585430000000
0!
0%
#585435000000
1!
1%
#585440000000
0!
0%
#585445000000
1!
1%
#585450000000
0!
0%
#585455000000
1!
1%
#585460000000
0!
0%
#585465000000
1!
1%
#585470000000
0!
0%
#585475000000
1!
1%
#585480000000
0!
0%
#585485000000
1!
1%
#585490000000
0!
0%
#585495000000
1!
1%
#585500000000
0!
0%
#585505000000
1!
1%
#585510000000
0!
0%
#585515000000
1!
1%
#585520000000
0!
0%
#585525000000
1!
1%
#585530000000
0!
0%
#585535000000
1!
1%
#585540000000
0!
0%
#585545000000
1!
1%
#585550000000
0!
0%
#585555000000
1!
1%
#585560000000
0!
0%
#585565000000
1!
1%
#585570000000
0!
0%
#585575000000
1!
1%
#585580000000
0!
0%
#585585000000
1!
1%
#585590000000
0!
0%
#585595000000
1!
1%
#585600000000
0!
0%
#585605000000
1!
1%
#585610000000
0!
0%
#585615000000
1!
1%
#585620000000
0!
0%
#585625000000
1!
1%
#585630000000
0!
0%
#585635000000
1!
1%
#585640000000
0!
0%
#585645000000
1!
1%
#585650000000
0!
0%
#585655000000
1!
1%
#585660000000
0!
0%
#585665000000
1!
1%
#585670000000
0!
0%
#585675000000
1!
1%
#585680000000
0!
0%
#585685000000
1!
1%
#585690000000
0!
0%
#585695000000
1!
1%
#585700000000
0!
0%
#585705000000
1!
1%
#585710000000
0!
0%
#585715000000
1!
1%
#585720000000
0!
0%
#585725000000
1!
1%
#585730000000
0!
0%
#585735000000
1!
1%
#585740000000
0!
0%
#585745000000
1!
1%
#585750000000
0!
0%
#585755000000
1!
1%
#585760000000
0!
0%
#585765000000
1!
1%
#585770000000
0!
0%
#585775000000
1!
1%
#585780000000
0!
0%
#585785000000
1!
1%
#585790000000
0!
0%
#585795000000
1!
1%
#585800000000
0!
0%
#585805000000
1!
1%
#585810000000
0!
0%
#585815000000
1!
1%
#585820000000
0!
0%
#585825000000
1!
1%
#585830000000
0!
0%
#585835000000
1!
1%
#585840000000
0!
0%
#585845000000
1!
1%
#585850000000
0!
0%
#585855000000
1!
1%
#585860000000
0!
0%
#585865000000
1!
1%
#585870000000
0!
0%
#585875000000
1!
1%
#585880000000
0!
0%
#585885000000
1!
1%
#585890000000
0!
0%
#585895000000
1!
1%
#585900000000
0!
0%
#585905000000
1!
1%
#585910000000
0!
0%
#585915000000
1!
1%
#585920000000
0!
0%
#585925000000
1!
1%
#585930000000
0!
0%
#585935000000
1!
1%
#585940000000
0!
0%
#585945000000
1!
1%
#585950000000
0!
0%
#585955000000
1!
1%
#585960000000
0!
0%
#585965000000
1!
1%
#585970000000
0!
0%
#585975000000
1!
1%
#585980000000
0!
0%
#585985000000
1!
1%
#585990000000
0!
0%
#585995000000
1!
1%
#586000000000
0!
0%
#586005000000
1!
1%
#586010000000
0!
0%
#586015000000
1!
1%
#586020000000
0!
0%
#586025000000
1!
1%
#586030000000
0!
0%
#586035000000
1!
1%
#586040000000
0!
0%
#586045000000
1!
1%
#586050000000
0!
0%
#586055000000
1!
1%
#586060000000
0!
0%
#586065000000
1!
1%
#586070000000
0!
0%
#586075000000
1!
1%
#586080000000
0!
0%
#586085000000
1!
1%
#586090000000
0!
0%
#586095000000
1!
1%
#586100000000
0!
0%
#586105000000
1!
1%
#586110000000
0!
0%
#586115000000
1!
1%
#586120000000
0!
0%
#586125000000
1!
1%
#586130000000
0!
0%
#586135000000
1!
1%
#586140000000
0!
0%
#586145000000
1!
1%
#586150000000
0!
0%
#586155000000
1!
1%
#586160000000
0!
0%
#586165000000
1!
1%
#586170000000
0!
0%
#586175000000
1!
1%
#586180000000
0!
0%
#586185000000
1!
1%
#586190000000
0!
0%
#586195000000
1!
1%
#586200000000
0!
0%
#586205000000
1!
1%
#586210000000
0!
0%
#586215000000
1!
1%
#586220000000
0!
0%
#586225000000
1!
1%
#586230000000
0!
0%
#586235000000
1!
1%
#586240000000
0!
0%
#586245000000
1!
1%
#586250000000
0!
0%
#586255000000
1!
1%
#586260000000
0!
0%
#586265000000
1!
1%
#586270000000
0!
0%
#586275000000
1!
1%
#586280000000
0!
0%
#586285000000
1!
1%
#586290000000
0!
0%
#586295000000
1!
1%
#586300000000
0!
0%
#586305000000
1!
1%
#586310000000
0!
0%
#586315000000
1!
1%
#586320000000
0!
0%
#586325000000
1!
1%
#586330000000
0!
0%
#586335000000
1!
1%
#586340000000
0!
0%
#586345000000
1!
1%
#586350000000
0!
0%
#586355000000
1!
1%
#586360000000
0!
0%
#586365000000
1!
1%
#586370000000
0!
0%
#586375000000
1!
1%
#586380000000
0!
0%
#586385000000
1!
1%
#586390000000
0!
0%
#586395000000
1!
1%
#586400000000
0!
0%
#586405000000
1!
1%
#586410000000
0!
0%
#586415000000
1!
1%
#586420000000
0!
0%
#586425000000
1!
1%
#586430000000
0!
0%
#586435000000
1!
1%
#586440000000
0!
0%
#586445000000
1!
1%
#586450000000
0!
0%
#586455000000
1!
1%
#586460000000
0!
0%
#586465000000
1!
1%
#586470000000
0!
0%
#586475000000
1!
1%
#586480000000
0!
0%
#586485000000
1!
1%
#586490000000
0!
0%
#586495000000
1!
1%
#586500000000
0!
0%
#586505000000
1!
1%
#586510000000
0!
0%
#586515000000
1!
1%
#586520000000
0!
0%
#586525000000
1!
1%
#586530000000
0!
0%
#586535000000
1!
1%
#586540000000
0!
0%
#586545000000
1!
1%
#586550000000
0!
0%
#586555000000
1!
1%
#586560000000
0!
0%
#586565000000
1!
1%
#586570000000
0!
0%
#586575000000
1!
1%
#586580000000
0!
0%
#586585000000
1!
1%
#586590000000
0!
0%
#586595000000
1!
1%
#586600000000
0!
0%
#586605000000
1!
1%
#586610000000
0!
0%
#586615000000
1!
1%
#586620000000
0!
0%
#586625000000
1!
1%
#586630000000
0!
0%
#586635000000
1!
1%
#586640000000
0!
0%
#586645000000
1!
1%
#586650000000
0!
0%
#586655000000
1!
1%
#586660000000
0!
0%
#586665000000
1!
1%
#586670000000
0!
0%
#586675000000
1!
1%
#586680000000
0!
0%
#586685000000
1!
1%
#586690000000
0!
0%
#586695000000
1!
1%
#586700000000
0!
0%
#586705000000
1!
1%
#586710000000
0!
0%
#586715000000
1!
1%
#586720000000
0!
0%
#586725000000
1!
1%
#586730000000
0!
0%
#586735000000
1!
1%
#586740000000
0!
0%
#586745000000
1!
1%
#586750000000
0!
0%
#586755000000
1!
1%
#586760000000
0!
0%
#586765000000
1!
1%
#586770000000
0!
0%
#586775000000
1!
1%
#586780000000
0!
0%
#586785000000
1!
1%
#586790000000
0!
0%
#586795000000
1!
1%
#586800000000
0!
0%
#586805000000
1!
1%
#586810000000
0!
0%
#586815000000
1!
1%
#586820000000
0!
0%
#586825000000
1!
1%
#586830000000
0!
0%
#586835000000
1!
1%
#586840000000
0!
0%
#586845000000
1!
1%
#586850000000
0!
0%
#586855000000
1!
1%
#586860000000
0!
0%
#586865000000
1!
1%
#586870000000
0!
0%
#586875000000
1!
1%
#586880000000
0!
0%
#586885000000
1!
1%
#586890000000
0!
0%
#586895000000
1!
1%
#586900000000
0!
0%
#586905000000
1!
1%
#586910000000
0!
0%
#586915000000
1!
1%
#586920000000
0!
0%
#586925000000
1!
1%
#586930000000
0!
0%
#586935000000
1!
1%
#586940000000
0!
0%
#586945000000
1!
1%
#586950000000
0!
0%
#586955000000
1!
1%
#586960000000
0!
0%
#586965000000
1!
1%
#586970000000
0!
0%
#586975000000
1!
1%
#586980000000
0!
0%
#586985000000
1!
1%
#586990000000
0!
0%
#586995000000
1!
1%
#587000000000
0!
0%
#587005000000
1!
1%
#587010000000
0!
0%
#587015000000
1!
1%
#587020000000
0!
0%
#587025000000
1!
1%
#587030000000
0!
0%
#587035000000
1!
1%
#587040000000
0!
0%
#587045000000
1!
1%
#587050000000
0!
0%
#587055000000
1!
1%
#587060000000
0!
0%
#587065000000
1!
1%
#587070000000
0!
0%
#587075000000
1!
1%
#587080000000
0!
0%
#587085000000
1!
1%
#587090000000
0!
0%
#587095000000
1!
1%
#587100000000
0!
0%
#587105000000
1!
1%
#587110000000
0!
0%
#587115000000
1!
1%
#587120000000
0!
0%
#587125000000
1!
1%
#587130000000
0!
0%
#587135000000
1!
1%
#587140000000
0!
0%
#587145000000
1!
1%
#587150000000
0!
0%
#587155000000
1!
1%
#587160000000
0!
0%
#587165000000
1!
1%
#587170000000
0!
0%
#587175000000
1!
1%
#587180000000
0!
0%
#587185000000
1!
1%
#587190000000
0!
0%
#587195000000
1!
1%
#587200000000
0!
0%
#587205000000
1!
1%
#587210000000
0!
0%
#587215000000
1!
1%
#587220000000
0!
0%
#587225000000
1!
1%
#587230000000
0!
0%
#587235000000
1!
1%
#587240000000
0!
0%
#587245000000
1!
1%
#587250000000
0!
0%
#587255000000
1!
1%
#587260000000
0!
0%
#587265000000
1!
1%
#587270000000
0!
0%
#587275000000
1!
1%
#587280000000
0!
0%
#587285000000
1!
1%
#587290000000
0!
0%
#587295000000
1!
1%
#587300000000
0!
0%
#587305000000
1!
1%
#587310000000
0!
0%
#587315000000
1!
1%
#587320000000
0!
0%
#587325000000
1!
1%
#587330000000
0!
0%
#587335000000
1!
1%
#587340000000
0!
0%
#587345000000
1!
1%
#587350000000
0!
0%
#587355000000
1!
1%
#587360000000
0!
0%
#587365000000
1!
1%
#587370000000
0!
0%
#587375000000
1!
1%
#587380000000
0!
0%
#587385000000
1!
1%
#587390000000
0!
0%
#587395000000
1!
1%
#587400000000
0!
0%
#587405000000
1!
1%
#587410000000
0!
0%
#587415000000
1!
1%
#587420000000
0!
0%
#587425000000
1!
1%
#587430000000
0!
0%
#587435000000
1!
1%
#587440000000
0!
0%
#587445000000
1!
1%
#587450000000
0!
0%
#587455000000
1!
1%
#587460000000
0!
0%
#587465000000
1!
1%
#587470000000
0!
0%
#587475000000
1!
1%
#587480000000
0!
0%
#587485000000
1!
1%
#587490000000
0!
0%
#587495000000
1!
1%
#587500000000
0!
0%
#587505000000
1!
1%
#587510000000
0!
0%
#587515000000
1!
1%
#587520000000
0!
0%
#587525000000
1!
1%
#587530000000
0!
0%
#587535000000
1!
1%
#587540000000
0!
0%
#587545000000
1!
1%
#587550000000
0!
0%
#587555000000
1!
1%
#587560000000
0!
0%
#587565000000
1!
1%
#587570000000
0!
0%
#587575000000
1!
1%
#587580000000
0!
0%
#587585000000
1!
1%
#587590000000
0!
0%
#587595000000
1!
1%
#587600000000
0!
0%
#587605000000
1!
1%
#587610000000
0!
0%
#587615000000
1!
1%
#587620000000
0!
0%
#587625000000
1!
1%
#587630000000
0!
0%
#587635000000
1!
1%
#587640000000
0!
0%
#587645000000
1!
1%
#587650000000
0!
0%
#587655000000
1!
1%
#587660000000
0!
0%
#587665000000
1!
1%
#587670000000
0!
0%
#587675000000
1!
1%
#587680000000
0!
0%
#587685000000
1!
1%
#587690000000
0!
0%
#587695000000
1!
1%
#587700000000
0!
0%
#587705000000
1!
1%
#587710000000
0!
0%
#587715000000
1!
1%
#587720000000
0!
0%
#587725000000
1!
1%
#587730000000
0!
0%
#587735000000
1!
1%
#587740000000
0!
0%
#587745000000
1!
1%
#587750000000
0!
0%
#587755000000
1!
1%
#587760000000
0!
0%
#587765000000
1!
1%
#587770000000
0!
0%
#587775000000
1!
1%
#587780000000
0!
0%
#587785000000
1!
1%
#587790000000
0!
0%
#587795000000
1!
1%
#587800000000
0!
0%
#587805000000
1!
1%
#587810000000
0!
0%
#587815000000
1!
1%
#587820000000
0!
0%
#587825000000
1!
1%
#587830000000
0!
0%
#587835000000
1!
1%
#587840000000
0!
0%
#587845000000
1!
1%
#587850000000
0!
0%
#587855000000
1!
1%
#587860000000
0!
0%
#587865000000
1!
1%
#587870000000
0!
0%
#587875000000
1!
1%
#587880000000
0!
0%
#587885000000
1!
1%
#587890000000
0!
0%
#587895000000
1!
1%
#587900000000
0!
0%
#587905000000
1!
1%
#587910000000
0!
0%
#587915000000
1!
1%
#587920000000
0!
0%
#587925000000
1!
1%
#587930000000
0!
0%
#587935000000
1!
1%
#587940000000
0!
0%
#587945000000
1!
1%
#587950000000
0!
0%
#587955000000
1!
1%
#587960000000
0!
0%
#587965000000
1!
1%
#587970000000
0!
0%
#587975000000
1!
1%
#587980000000
0!
0%
#587985000000
1!
1%
#587990000000
0!
0%
#587995000000
1!
1%
#588000000000
0!
0%
#588005000000
1!
1%
#588010000000
0!
0%
#588015000000
1!
1%
#588020000000
0!
0%
#588025000000
1!
1%
#588030000000
0!
0%
#588035000000
1!
1%
#588040000000
0!
0%
#588045000000
1!
1%
#588050000000
0!
0%
#588055000000
1!
1%
#588060000000
0!
0%
#588065000000
1!
1%
#588070000000
0!
0%
#588075000000
1!
1%
#588080000000
0!
0%
#588085000000
1!
1%
#588090000000
0!
0%
#588095000000
1!
1%
#588100000000
0!
0%
#588105000000
1!
1%
#588110000000
0!
0%
#588115000000
1!
1%
#588120000000
0!
0%
#588125000000
1!
1%
#588130000000
0!
0%
#588135000000
1!
1%
#588140000000
0!
0%
#588145000000
1!
1%
#588150000000
0!
0%
#588155000000
1!
1%
#588160000000
0!
0%
#588165000000
1!
1%
#588170000000
0!
0%
#588175000000
1!
1%
#588180000000
0!
0%
#588185000000
1!
1%
#588190000000
0!
0%
#588195000000
1!
1%
#588200000000
0!
0%
#588205000000
1!
1%
#588210000000
0!
0%
#588215000000
1!
1%
#588220000000
0!
0%
#588225000000
1!
1%
#588230000000
0!
0%
#588235000000
1!
1%
#588240000000
0!
0%
#588245000000
1!
1%
#588250000000
0!
0%
#588255000000
1!
1%
#588260000000
0!
0%
#588265000000
1!
1%
#588270000000
0!
0%
#588275000000
1!
1%
#588280000000
0!
0%
#588285000000
1!
1%
#588290000000
0!
0%
#588295000000
1!
1%
#588300000000
0!
0%
#588305000000
1!
1%
#588310000000
0!
0%
#588315000000
1!
1%
#588320000000
0!
0%
#588325000000
1!
1%
#588330000000
0!
0%
#588335000000
1!
1%
#588340000000
0!
0%
#588345000000
1!
1%
#588350000000
0!
0%
#588355000000
1!
1%
#588360000000
0!
0%
#588365000000
1!
1%
#588370000000
0!
0%
#588375000000
1!
1%
#588380000000
0!
0%
#588385000000
1!
1%
#588390000000
0!
0%
#588395000000
1!
1%
#588400000000
0!
0%
#588405000000
1!
1%
#588410000000
0!
0%
#588415000000
1!
1%
#588420000000
0!
0%
#588425000000
1!
1%
#588430000000
0!
0%
#588435000000
1!
1%
#588440000000
0!
0%
#588445000000
1!
1%
#588450000000
0!
0%
#588455000000
1!
1%
#588460000000
0!
0%
#588465000000
1!
1%
#588470000000
0!
0%
#588475000000
1!
1%
#588480000000
0!
0%
#588485000000
1!
1%
#588490000000
0!
0%
#588495000000
1!
1%
#588500000000
0!
0%
#588505000000
1!
1%
#588510000000
0!
0%
#588515000000
1!
1%
#588520000000
0!
0%
#588525000000
1!
1%
#588530000000
0!
0%
#588535000000
1!
1%
#588540000000
0!
0%
#588545000000
1!
1%
#588550000000
0!
0%
#588555000000
1!
1%
#588560000000
0!
0%
#588565000000
1!
1%
#588570000000
0!
0%
#588575000000
1!
1%
#588580000000
0!
0%
#588585000000
1!
1%
#588590000000
0!
0%
#588595000000
1!
1%
#588600000000
0!
0%
#588605000000
1!
1%
#588610000000
0!
0%
#588615000000
1!
1%
#588620000000
0!
0%
#588625000000
1!
1%
#588630000000
0!
0%
#588635000000
1!
1%
#588640000000
0!
0%
#588645000000
1!
1%
#588650000000
0!
0%
#588655000000
1!
1%
#588660000000
0!
0%
#588665000000
1!
1%
#588670000000
0!
0%
#588675000000
1!
1%
#588680000000
0!
0%
#588685000000
1!
1%
#588690000000
0!
0%
#588695000000
1!
1%
#588700000000
0!
0%
#588705000000
1!
1%
#588710000000
0!
0%
#588715000000
1!
1%
#588720000000
0!
0%
#588725000000
1!
1%
#588730000000
0!
0%
#588735000000
1!
1%
#588740000000
0!
0%
#588745000000
1!
1%
#588750000000
0!
0%
#588755000000
1!
1%
#588760000000
0!
0%
#588765000000
1!
1%
#588770000000
0!
0%
#588775000000
1!
1%
#588780000000
0!
0%
#588785000000
1!
1%
#588790000000
0!
0%
#588795000000
1!
1%
#588800000000
0!
0%
#588805000000
1!
1%
#588810000000
0!
0%
#588815000000
1!
1%
#588820000000
0!
0%
#588825000000
1!
1%
#588830000000
0!
0%
#588835000000
1!
1%
#588840000000
0!
0%
#588845000000
1!
1%
#588850000000
0!
0%
#588855000000
1!
1%
#588860000000
0!
0%
#588865000000
1!
1%
#588870000000
0!
0%
#588875000000
1!
1%
#588880000000
0!
0%
#588885000000
1!
1%
#588890000000
0!
0%
#588895000000
1!
1%
#588900000000
0!
0%
#588905000000
1!
1%
#588910000000
0!
0%
#588915000000
1!
1%
#588920000000
0!
0%
#588925000000
1!
1%
#588930000000
0!
0%
#588935000000
1!
1%
#588940000000
0!
0%
#588945000000
1!
1%
#588950000000
0!
0%
#588955000000
1!
1%
#588960000000
0!
0%
#588965000000
1!
1%
#588970000000
0!
0%
#588975000000
1!
1%
#588980000000
0!
0%
#588985000000
1!
1%
#588990000000
0!
0%
#588995000000
1!
1%
#589000000000
0!
0%
#589005000000
1!
1%
#589010000000
0!
0%
#589015000000
1!
1%
#589020000000
0!
0%
#589025000000
1!
1%
#589030000000
0!
0%
#589035000000
1!
1%
#589040000000
0!
0%
#589045000000
1!
1%
#589050000000
0!
0%
#589055000000
1!
1%
#589060000000
0!
0%
#589065000000
1!
1%
#589070000000
0!
0%
#589075000000
1!
1%
#589080000000
0!
0%
#589085000000
1!
1%
#589090000000
0!
0%
#589095000000
1!
1%
#589100000000
0!
0%
#589105000000
1!
1%
#589110000000
0!
0%
#589115000000
1!
1%
#589120000000
0!
0%
#589125000000
1!
1%
#589130000000
0!
0%
#589135000000
1!
1%
#589140000000
0!
0%
#589145000000
1!
1%
#589150000000
0!
0%
#589155000000
1!
1%
#589160000000
0!
0%
#589165000000
1!
1%
#589170000000
0!
0%
#589175000000
1!
1%
#589180000000
0!
0%
#589185000000
1!
1%
#589190000000
0!
0%
#589195000000
1!
1%
#589200000000
0!
0%
#589205000000
1!
1%
#589210000000
0!
0%
#589215000000
1!
1%
#589220000000
0!
0%
#589225000000
1!
1%
#589230000000
0!
0%
#589235000000
1!
1%
#589240000000
0!
0%
#589245000000
1!
1%
#589250000000
0!
0%
#589255000000
1!
1%
#589260000000
0!
0%
#589265000000
1!
1%
#589270000000
0!
0%
#589275000000
1!
1%
#589280000000
0!
0%
#589285000000
1!
1%
#589290000000
0!
0%
#589295000000
1!
1%
#589300000000
0!
0%
#589305000000
1!
1%
#589310000000
0!
0%
#589315000000
1!
1%
#589320000000
0!
0%
#589325000000
1!
1%
#589330000000
0!
0%
#589335000000
1!
1%
#589340000000
0!
0%
#589345000000
1!
1%
#589350000000
0!
0%
#589355000000
1!
1%
#589360000000
0!
0%
#589365000000
1!
1%
#589370000000
0!
0%
#589375000000
1!
1%
#589380000000
0!
0%
#589385000000
1!
1%
#589390000000
0!
0%
#589395000000
1!
1%
#589400000000
0!
0%
#589405000000
1!
1%
#589410000000
0!
0%
#589415000000
1!
1%
#589420000000
0!
0%
#589425000000
1!
1%
#589430000000
0!
0%
#589435000000
1!
1%
#589440000000
0!
0%
#589445000000
1!
1%
#589450000000
0!
0%
#589455000000
1!
1%
#589460000000
0!
0%
#589465000000
1!
1%
#589470000000
0!
0%
#589475000000
1!
1%
#589480000000
0!
0%
#589485000000
1!
1%
#589490000000
0!
0%
#589495000000
1!
1%
#589500000000
0!
0%
#589505000000
1!
1%
#589510000000
0!
0%
#589515000000
1!
1%
#589520000000
0!
0%
#589525000000
1!
1%
#589530000000
0!
0%
#589535000000
1!
1%
#589540000000
0!
0%
#589545000000
1!
1%
#589550000000
0!
0%
#589555000000
1!
1%
#589560000000
0!
0%
#589565000000
1!
1%
#589570000000
0!
0%
#589575000000
1!
1%
#589580000000
0!
0%
#589585000000
1!
1%
#589590000000
0!
0%
#589595000000
1!
1%
#589600000000
0!
0%
#589605000000
1!
1%
#589610000000
0!
0%
#589615000000
1!
1%
#589620000000
0!
0%
#589625000000
1!
1%
#589630000000
0!
0%
#589635000000
1!
1%
#589640000000
0!
0%
#589645000000
1!
1%
#589650000000
0!
0%
#589655000000
1!
1%
#589660000000
0!
0%
#589665000000
1!
1%
#589670000000
0!
0%
#589675000000
1!
1%
#589680000000
0!
0%
#589685000000
1!
1%
#589690000000
0!
0%
#589695000000
1!
1%
#589700000000
0!
0%
#589705000000
1!
1%
#589710000000
0!
0%
#589715000000
1!
1%
#589720000000
0!
0%
#589725000000
1!
1%
#589730000000
0!
0%
#589735000000
1!
1%
#589740000000
0!
0%
#589745000000
1!
1%
#589750000000
0!
0%
#589755000000
1!
1%
#589760000000
0!
0%
#589765000000
1!
1%
#589770000000
0!
0%
#589775000000
1!
1%
#589780000000
0!
0%
#589785000000
1!
1%
#589790000000
0!
0%
#589795000000
1!
1%
#589800000000
0!
0%
#589805000000
1!
1%
#589810000000
0!
0%
#589815000000
1!
1%
#589820000000
0!
0%
#589825000000
1!
1%
#589830000000
0!
0%
#589835000000
1!
1%
#589840000000
0!
0%
#589845000000
1!
1%
#589850000000
0!
0%
#589855000000
1!
1%
#589860000000
0!
0%
#589865000000
1!
1%
#589870000000
0!
0%
#589875000000
1!
1%
#589880000000
0!
0%
#589885000000
1!
1%
#589890000000
0!
0%
#589895000000
1!
1%
#589900000000
0!
0%
#589905000000
1!
1%
#589910000000
0!
0%
#589915000000
1!
1%
#589920000000
0!
0%
#589925000000
1!
1%
#589930000000
0!
0%
#589935000000
1!
1%
#589940000000
0!
0%
#589945000000
1!
1%
#589950000000
0!
0%
#589955000000
1!
1%
#589960000000
0!
0%
#589965000000
1!
1%
#589970000000
0!
0%
#589975000000
1!
1%
#589980000000
0!
0%
#589985000000
1!
1%
#589990000000
0!
0%
#589995000000
1!
1%
#590000000000
0!
0%
#590005000000
1!
1%
#590010000000
0!
0%
#590015000000
1!
1%
#590020000000
0!
0%
#590025000000
1!
1%
#590030000000
0!
0%
#590035000000
1!
1%
#590040000000
0!
0%
#590045000000
1!
1%
#590050000000
0!
0%
#590055000000
1!
1%
#590060000000
0!
0%
#590065000000
1!
1%
#590070000000
0!
0%
#590075000000
1!
1%
#590080000000
0!
0%
#590085000000
1!
1%
#590090000000
0!
0%
#590095000000
1!
1%
#590100000000
0!
0%
#590105000000
1!
1%
#590110000000
0!
0%
#590115000000
1!
1%
#590120000000
0!
0%
#590125000000
1!
1%
#590130000000
0!
0%
#590135000000
1!
1%
#590140000000
0!
0%
#590145000000
1!
1%
#590150000000
0!
0%
#590155000000
1!
1%
#590160000000
0!
0%
#590165000000
1!
1%
#590170000000
0!
0%
#590175000000
1!
1%
#590180000000
0!
0%
#590185000000
1!
1%
#590190000000
0!
0%
#590195000000
1!
1%
#590200000000
0!
0%
#590205000000
1!
1%
#590210000000
0!
0%
#590215000000
1!
1%
#590220000000
0!
0%
#590225000000
1!
1%
#590230000000
0!
0%
#590235000000
1!
1%
#590240000000
0!
0%
#590245000000
1!
1%
#590250000000
0!
0%
#590255000000
1!
1%
#590260000000
0!
0%
#590265000000
1!
1%
#590270000000
0!
0%
#590275000000
1!
1%
#590280000000
0!
0%
#590285000000
1!
1%
#590290000000
0!
0%
#590295000000
1!
1%
#590300000000
0!
0%
#590305000000
1!
1%
#590310000000
0!
0%
#590315000000
1!
1%
#590320000000
0!
0%
#590325000000
1!
1%
#590330000000
0!
0%
#590335000000
1!
1%
#590340000000
0!
0%
#590345000000
1!
1%
#590350000000
0!
0%
#590355000000
1!
1%
#590360000000
0!
0%
#590365000000
1!
1%
#590370000000
0!
0%
#590375000000
1!
1%
#590380000000
0!
0%
#590385000000
1!
1%
#590390000000
0!
0%
#590395000000
1!
1%
#590400000000
0!
0%
#590405000000
1!
1%
#590410000000
0!
0%
#590415000000
1!
1%
#590420000000
0!
0%
#590425000000
1!
1%
#590430000000
0!
0%
#590435000000
1!
1%
#590440000000
0!
0%
#590445000000
1!
1%
#590450000000
0!
0%
#590455000000
1!
1%
#590460000000
0!
0%
#590465000000
1!
1%
#590470000000
0!
0%
#590475000000
1!
1%
#590480000000
0!
0%
#590485000000
1!
1%
#590490000000
0!
0%
#590495000000
1!
1%
#590500000000
0!
0%
#590505000000
1!
1%
#590510000000
0!
0%
#590515000000
1!
1%
#590520000000
0!
0%
#590525000000
1!
1%
#590530000000
0!
0%
#590535000000
1!
1%
#590540000000
0!
0%
#590545000000
1!
1%
#590550000000
0!
0%
#590555000000
1!
1%
#590560000000
0!
0%
#590565000000
1!
1%
#590570000000
0!
0%
#590575000000
1!
1%
#590580000000
0!
0%
#590585000000
1!
1%
#590590000000
0!
0%
#590595000000
1!
1%
#590600000000
0!
0%
#590605000000
1!
1%
#590610000000
0!
0%
#590615000000
1!
1%
#590620000000
0!
0%
#590625000000
1!
1%
#590630000000
0!
0%
#590635000000
1!
1%
#590640000000
0!
0%
#590645000000
1!
1%
#590650000000
0!
0%
#590655000000
1!
1%
#590660000000
0!
0%
#590665000000
1!
1%
#590670000000
0!
0%
#590675000000
1!
1%
#590680000000
0!
0%
#590685000000
1!
1%
#590690000000
0!
0%
#590695000000
1!
1%
#590700000000
0!
0%
#590705000000
1!
1%
#590710000000
0!
0%
#590715000000
1!
1%
#590720000000
0!
0%
#590725000000
1!
1%
#590730000000
0!
0%
#590735000000
1!
1%
#590740000000
0!
0%
#590745000000
1!
1%
#590750000000
0!
0%
#590755000000
1!
1%
#590760000000
0!
0%
#590765000000
1!
1%
#590770000000
0!
0%
#590775000000
1!
1%
#590780000000
0!
0%
#590785000000
1!
1%
#590790000000
0!
0%
#590795000000
1!
1%
#590800000000
0!
0%
#590805000000
1!
1%
#590810000000
0!
0%
#590815000000
1!
1%
#590820000000
0!
0%
#590825000000
1!
1%
#590830000000
0!
0%
#590835000000
1!
1%
#590840000000
0!
0%
#590845000000
1!
1%
#590850000000
0!
0%
#590855000000
1!
1%
#590860000000
0!
0%
#590865000000
1!
1%
#590870000000
0!
0%
#590875000000
1!
1%
#590880000000
0!
0%
#590885000000
1!
1%
#590890000000
0!
0%
#590895000000
1!
1%
#590900000000
0!
0%
#590905000000
1!
1%
#590910000000
0!
0%
#590915000000
1!
1%
#590920000000
0!
0%
#590925000000
1!
1%
#590930000000
0!
0%
#590935000000
1!
1%
#590940000000
0!
0%
#590945000000
1!
1%
#590950000000
0!
0%
#590955000000
1!
1%
#590960000000
0!
0%
#590965000000
1!
1%
#590970000000
0!
0%
#590975000000
1!
1%
#590980000000
0!
0%
#590985000000
1!
1%
#590990000000
0!
0%
#590995000000
1!
1%
#591000000000
0!
0%
#591005000000
1!
1%
#591010000000
0!
0%
#591015000000
1!
1%
#591020000000
0!
0%
#591025000000
1!
1%
#591030000000
0!
0%
#591035000000
1!
1%
#591040000000
0!
0%
#591045000000
1!
1%
#591050000000
0!
0%
#591055000000
1!
1%
#591060000000
0!
0%
#591065000000
1!
1%
#591070000000
0!
0%
#591075000000
1!
1%
#591080000000
0!
0%
#591085000000
1!
1%
#591090000000
0!
0%
#591095000000
1!
1%
#591100000000
0!
0%
#591105000000
1!
1%
#591110000000
0!
0%
#591115000000
1!
1%
#591120000000
0!
0%
#591125000000
1!
1%
#591130000000
0!
0%
#591135000000
1!
1%
#591140000000
0!
0%
#591145000000
1!
1%
#591150000000
0!
0%
#591155000000
1!
1%
#591160000000
0!
0%
#591165000000
1!
1%
#591170000000
0!
0%
#591175000000
1!
1%
#591180000000
0!
0%
#591185000000
1!
1%
#591190000000
0!
0%
#591195000000
1!
1%
#591200000000
0!
0%
#591205000000
1!
1%
#591210000000
0!
0%
#591215000000
1!
1%
#591220000000
0!
0%
#591225000000
1!
1%
#591230000000
0!
0%
#591235000000
1!
1%
#591240000000
0!
0%
#591245000000
1!
1%
#591250000000
0!
0%
#591255000000
1!
1%
#591260000000
0!
0%
#591265000000
1!
1%
#591270000000
0!
0%
#591275000000
1!
1%
#591280000000
0!
0%
#591285000000
1!
1%
#591290000000
0!
0%
#591295000000
1!
1%
#591300000000
0!
0%
#591305000000
1!
1%
#591310000000
0!
0%
#591315000000
1!
1%
#591320000000
0!
0%
#591325000000
1!
1%
#591330000000
0!
0%
#591335000000
1!
1%
#591340000000
0!
0%
#591345000000
1!
1%
#591350000000
0!
0%
#591355000000
1!
1%
#591360000000
0!
0%
#591365000000
1!
1%
#591370000000
0!
0%
#591375000000
1!
1%
#591380000000
0!
0%
#591385000000
1!
1%
#591390000000
0!
0%
#591395000000
1!
1%
#591400000000
0!
0%
#591405000000
1!
1%
#591410000000
0!
0%
#591415000000
1!
1%
#591420000000
0!
0%
#591425000000
1!
1%
#591430000000
0!
0%
#591435000000
1!
1%
#591440000000
0!
0%
#591445000000
1!
1%
#591450000000
0!
0%
#591455000000
1!
1%
#591460000000
0!
0%
#591465000000
1!
1%
#591470000000
0!
0%
#591475000000
1!
1%
#591480000000
0!
0%
#591485000000
1!
1%
#591490000000
0!
0%
#591495000000
1!
1%
#591500000000
0!
0%
#591505000000
1!
1%
#591510000000
0!
0%
#591515000000
1!
1%
#591520000000
0!
0%
#591525000000
1!
1%
#591530000000
0!
0%
#591535000000
1!
1%
#591540000000
0!
0%
#591545000000
1!
1%
#591550000000
0!
0%
#591555000000
1!
1%
#591560000000
0!
0%
#591565000000
1!
1%
#591570000000
0!
0%
#591575000000
1!
1%
#591580000000
0!
0%
#591585000000
1!
1%
#591590000000
0!
0%
#591595000000
1!
1%
#591600000000
0!
0%
#591605000000
1!
1%
#591610000000
0!
0%
#591615000000
1!
1%
#591620000000
0!
0%
#591625000000
1!
1%
#591630000000
0!
0%
#591635000000
1!
1%
#591640000000
0!
0%
#591645000000
1!
1%
#591650000000
0!
0%
#591655000000
1!
1%
#591660000000
0!
0%
#591665000000
1!
1%
#591670000000
0!
0%
#591675000000
1!
1%
#591680000000
0!
0%
#591685000000
1!
1%
#591690000000
0!
0%
#591695000000
1!
1%
#591700000000
0!
0%
#591705000000
1!
1%
#591710000000
0!
0%
#591715000000
1!
1%
#591720000000
0!
0%
#591725000000
1!
1%
#591730000000
0!
0%
#591735000000
1!
1%
#591740000000
0!
0%
#591745000000
1!
1%
#591750000000
0!
0%
#591755000000
1!
1%
#591760000000
0!
0%
#591765000000
1!
1%
#591770000000
0!
0%
#591775000000
1!
1%
#591780000000
0!
0%
#591785000000
1!
1%
#591790000000
0!
0%
#591795000000
1!
1%
#591800000000
0!
0%
#591805000000
1!
1%
#591810000000
0!
0%
#591815000000
1!
1%
#591820000000
0!
0%
#591825000000
1!
1%
#591830000000
0!
0%
#591835000000
1!
1%
#591840000000
0!
0%
#591845000000
1!
1%
#591850000000
0!
0%
#591855000000
1!
1%
#591860000000
0!
0%
#591865000000
1!
1%
#591870000000
0!
0%
#591875000000
1!
1%
#591880000000
0!
0%
#591885000000
1!
1%
#591890000000
0!
0%
#591895000000
1!
1%
#591900000000
0!
0%
#591905000000
1!
1%
#591910000000
0!
0%
#591915000000
1!
1%
#591920000000
0!
0%
#591925000000
1!
1%
#591930000000
0!
0%
#591935000000
1!
1%
#591940000000
0!
0%
#591945000000
1!
1%
#591950000000
0!
0%
#591955000000
1!
1%
#591960000000
0!
0%
#591965000000
1!
1%
#591970000000
0!
0%
#591975000000
1!
1%
#591980000000
0!
0%
#591985000000
1!
1%
#591990000000
0!
0%
#591995000000
1!
1%
#592000000000
0!
0%
#592005000000
1!
1%
#592010000000
0!
0%
#592015000000
1!
1%
#592020000000
0!
0%
#592025000000
1!
1%
#592030000000
0!
0%
#592035000000
1!
1%
#592040000000
0!
0%
#592045000000
1!
1%
#592050000000
0!
0%
#592055000000
1!
1%
#592060000000
0!
0%
#592065000000
1!
1%
#592070000000
0!
0%
#592075000000
1!
1%
#592080000000
0!
0%
#592085000000
1!
1%
#592090000000
0!
0%
#592095000000
1!
1%
#592100000000
0!
0%
#592105000000
1!
1%
#592110000000
0!
0%
#592115000000
1!
1%
#592120000000
0!
0%
#592125000000
1!
1%
#592130000000
0!
0%
#592135000000
1!
1%
#592140000000
0!
0%
#592145000000
1!
1%
#592150000000
0!
0%
#592155000000
1!
1%
#592160000000
0!
0%
#592165000000
1!
1%
#592170000000
0!
0%
#592175000000
1!
1%
#592180000000
0!
0%
#592185000000
1!
1%
#592190000000
0!
0%
#592195000000
1!
1%
#592200000000
0!
0%
#592205000000
1!
1%
#592210000000
0!
0%
#592215000000
1!
1%
#592220000000
0!
0%
#592225000000
1!
1%
#592230000000
0!
0%
#592235000000
1!
1%
#592240000000
0!
0%
#592245000000
1!
1%
#592250000000
0!
0%
#592255000000
1!
1%
#592260000000
0!
0%
#592265000000
1!
1%
#592270000000
0!
0%
#592275000000
1!
1%
#592280000000
0!
0%
#592285000000
1!
1%
#592290000000
0!
0%
#592295000000
1!
1%
#592300000000
0!
0%
#592305000000
1!
1%
#592310000000
0!
0%
#592315000000
1!
1%
#592320000000
0!
0%
#592325000000
1!
1%
#592330000000
0!
0%
#592335000000
1!
1%
#592340000000
0!
0%
#592345000000
1!
1%
#592350000000
0!
0%
#592355000000
1!
1%
#592360000000
0!
0%
#592365000000
1!
1%
#592370000000
0!
0%
#592375000000
1!
1%
#592380000000
0!
0%
#592385000000
1!
1%
#592390000000
0!
0%
#592395000000
1!
1%
#592400000000
0!
0%
#592405000000
1!
1%
#592410000000
0!
0%
#592415000000
1!
1%
#592420000000
0!
0%
#592425000000
1!
1%
#592430000000
0!
0%
#592435000000
1!
1%
#592440000000
0!
0%
#592445000000
1!
1%
#592450000000
0!
0%
#592455000000
1!
1%
#592460000000
0!
0%
#592465000000
1!
1%
#592470000000
0!
0%
#592475000000
1!
1%
#592480000000
0!
0%
#592485000000
1!
1%
#592490000000
0!
0%
#592495000000
1!
1%
#592500000000
0!
0%
#592505000000
1!
1%
#592510000000
0!
0%
#592515000000
1!
1%
#592520000000
0!
0%
#592525000000
1!
1%
#592530000000
0!
0%
#592535000000
1!
1%
#592540000000
0!
0%
#592545000000
1!
1%
#592550000000
0!
0%
#592555000000
1!
1%
#592560000000
0!
0%
#592565000000
1!
1%
#592570000000
0!
0%
#592575000000
1!
1%
#592580000000
0!
0%
#592585000000
1!
1%
#592590000000
0!
0%
#592595000000
1!
1%
#592600000000
0!
0%
#592605000000
1!
1%
#592610000000
0!
0%
#592615000000
1!
1%
#592620000000
0!
0%
#592625000000
1!
1%
#592630000000
0!
0%
#592635000000
1!
1%
#592640000000
0!
0%
#592645000000
1!
1%
#592650000000
0!
0%
#592655000000
1!
1%
#592660000000
0!
0%
#592665000000
1!
1%
#592670000000
0!
0%
#592675000000
1!
1%
#592680000000
0!
0%
#592685000000
1!
1%
#592690000000
0!
0%
#592695000000
1!
1%
#592700000000
0!
0%
#592705000000
1!
1%
#592710000000
0!
0%
#592715000000
1!
1%
#592720000000
0!
0%
#592725000000
1!
1%
#592730000000
0!
0%
#592735000000
1!
1%
#592740000000
0!
0%
#592745000000
1!
1%
#592750000000
0!
0%
#592755000000
1!
1%
#592760000000
0!
0%
#592765000000
1!
1%
#592770000000
0!
0%
#592775000000
1!
1%
#592780000000
0!
0%
#592785000000
1!
1%
#592790000000
0!
0%
#592795000000
1!
1%
#592800000000
0!
0%
#592805000000
1!
1%
#592810000000
0!
0%
#592815000000
1!
1%
#592820000000
0!
0%
#592825000000
1!
1%
#592830000000
0!
0%
#592835000000
1!
1%
#592840000000
0!
0%
#592845000000
1!
1%
#592850000000
0!
0%
#592855000000
1!
1%
#592860000000
0!
0%
#592865000000
1!
1%
#592870000000
0!
0%
#592875000000
1!
1%
#592880000000
0!
0%
#592885000000
1!
1%
#592890000000
0!
0%
#592895000000
1!
1%
#592900000000
0!
0%
#592905000000
1!
1%
#592910000000
0!
0%
#592915000000
1!
1%
#592920000000
0!
0%
#592925000000
1!
1%
#592930000000
0!
0%
#592935000000
1!
1%
#592940000000
0!
0%
#592945000000
1!
1%
#592950000000
0!
0%
#592955000000
1!
1%
#592960000000
0!
0%
#592965000000
1!
1%
#592970000000
0!
0%
#592975000000
1!
1%
#592980000000
0!
0%
#592985000000
1!
1%
#592990000000
0!
0%
#592995000000
1!
1%
#593000000000
0!
0%
#593005000000
1!
1%
#593010000000
0!
0%
#593015000000
1!
1%
#593020000000
0!
0%
#593025000000
1!
1%
#593030000000
0!
0%
#593035000000
1!
1%
#593040000000
0!
0%
#593045000000
1!
1%
#593050000000
0!
0%
#593055000000
1!
1%
#593060000000
0!
0%
#593065000000
1!
1%
#593070000000
0!
0%
#593075000000
1!
1%
#593080000000
0!
0%
#593085000000
1!
1%
#593090000000
0!
0%
#593095000000
1!
1%
#593100000000
0!
0%
#593105000000
1!
1%
#593110000000
0!
0%
#593115000000
1!
1%
#593120000000
0!
0%
#593125000000
1!
1%
#593130000000
0!
0%
#593135000000
1!
1%
#593140000000
0!
0%
#593145000000
1!
1%
#593150000000
0!
0%
#593155000000
1!
1%
#593160000000
0!
0%
#593165000000
1!
1%
#593170000000
0!
0%
#593175000000
1!
1%
#593180000000
0!
0%
#593185000000
1!
1%
#593190000000
0!
0%
#593195000000
1!
1%
#593200000000
0!
0%
#593205000000
1!
1%
#593210000000
0!
0%
#593215000000
1!
1%
#593220000000
0!
0%
#593225000000
1!
1%
#593230000000
0!
0%
#593235000000
1!
1%
#593240000000
0!
0%
#593245000000
1!
1%
#593250000000
0!
0%
#593255000000
1!
1%
#593260000000
0!
0%
#593265000000
1!
1%
#593270000000
0!
0%
#593275000000
1!
1%
#593280000000
0!
0%
#593285000000
1!
1%
#593290000000
0!
0%
#593295000000
1!
1%
#593300000000
0!
0%
#593305000000
1!
1%
#593310000000
0!
0%
#593315000000
1!
1%
#593320000000
0!
0%
#593325000000
1!
1%
#593330000000
0!
0%
#593335000000
1!
1%
#593340000000
0!
0%
#593345000000
1!
1%
#593350000000
0!
0%
#593355000000
1!
1%
#593360000000
0!
0%
#593365000000
1!
1%
#593370000000
0!
0%
#593375000000
1!
1%
#593380000000
0!
0%
#593385000000
1!
1%
#593390000000
0!
0%
#593395000000
1!
1%
#593400000000
0!
0%
#593405000000
1!
1%
#593410000000
0!
0%
#593415000000
1!
1%
#593420000000
0!
0%
#593425000000
1!
1%
#593430000000
0!
0%
#593435000000
1!
1%
#593440000000
0!
0%
#593445000000
1!
1%
#593450000000
0!
0%
#593455000000
1!
1%
#593460000000
0!
0%
#593465000000
1!
1%
#593470000000
0!
0%
#593475000000
1!
1%
#593480000000
0!
0%
#593485000000
1!
1%
#593490000000
0!
0%
#593495000000
1!
1%
#593500000000
0!
0%
#593505000000
1!
1%
#593510000000
0!
0%
#593515000000
1!
1%
#593520000000
0!
0%
#593525000000
1!
1%
#593530000000
0!
0%
#593535000000
1!
1%
#593540000000
0!
0%
#593545000000
1!
1%
#593550000000
0!
0%
#593555000000
1!
1%
#593560000000
0!
0%
#593565000000
1!
1%
#593570000000
0!
0%
#593575000000
1!
1%
#593580000000
0!
0%
#593585000000
1!
1%
#593590000000
0!
0%
#593595000000
1!
1%
#593600000000
0!
0%
#593605000000
1!
1%
#593610000000
0!
0%
#593615000000
1!
1%
#593620000000
0!
0%
#593625000000
1!
1%
#593630000000
0!
0%
#593635000000
1!
1%
#593640000000
0!
0%
#593645000000
1!
1%
#593650000000
0!
0%
#593655000000
1!
1%
#593660000000
0!
0%
#593665000000
1!
1%
#593670000000
0!
0%
#593675000000
1!
1%
#593680000000
0!
0%
#593685000000
1!
1%
#593690000000
0!
0%
#593695000000
1!
1%
#593700000000
0!
0%
#593705000000
1!
1%
#593710000000
0!
0%
#593715000000
1!
1%
#593720000000
0!
0%
#593725000000
1!
1%
#593730000000
0!
0%
#593735000000
1!
1%
#593740000000
0!
0%
#593745000000
1!
1%
#593750000000
0!
0%
#593755000000
1!
1%
#593760000000
0!
0%
#593765000000
1!
1%
#593770000000
0!
0%
#593775000000
1!
1%
#593780000000
0!
0%
#593785000000
1!
1%
#593790000000
0!
0%
#593795000000
1!
1%
#593800000000
0!
0%
#593805000000
1!
1%
#593810000000
0!
0%
#593815000000
1!
1%
#593820000000
0!
0%
#593825000000
1!
1%
#593830000000
0!
0%
#593835000000
1!
1%
#593840000000
0!
0%
#593845000000
1!
1%
#593850000000
0!
0%
#593855000000
1!
1%
#593860000000
0!
0%
#593865000000
1!
1%
#593870000000
0!
0%
#593875000000
1!
1%
#593880000000
0!
0%
#593885000000
1!
1%
#593890000000
0!
0%
#593895000000
1!
1%
#593900000000
0!
0%
#593905000000
1!
1%
#593910000000
0!
0%
#593915000000
1!
1%
#593920000000
0!
0%
#593925000000
1!
1%
#593930000000
0!
0%
#593935000000
1!
1%
#593940000000
0!
0%
#593945000000
1!
1%
#593950000000
0!
0%
#593955000000
1!
1%
#593960000000
0!
0%
#593965000000
1!
1%
#593970000000
0!
0%
#593975000000
1!
1%
#593980000000
0!
0%
#593985000000
1!
1%
#593990000000
0!
0%
#593995000000
1!
1%
#594000000000
0!
0%
#594005000000
1!
1%
#594010000000
0!
0%
#594015000000
1!
1%
#594020000000
0!
0%
#594025000000
1!
1%
#594030000000
0!
0%
#594035000000
1!
1%
#594040000000
0!
0%
#594045000000
1!
1%
#594050000000
0!
0%
#594055000000
1!
1%
#594060000000
0!
0%
#594065000000
1!
1%
#594070000000
0!
0%
#594075000000
1!
1%
#594080000000
0!
0%
#594085000000
1!
1%
#594090000000
0!
0%
#594095000000
1!
1%
#594100000000
0!
0%
#594105000000
1!
1%
#594110000000
0!
0%
#594115000000
1!
1%
#594120000000
0!
0%
#594125000000
1!
1%
#594130000000
0!
0%
#594135000000
1!
1%
#594140000000
0!
0%
#594145000000
1!
1%
#594150000000
0!
0%
#594155000000
1!
1%
#594160000000
0!
0%
#594165000000
1!
1%
#594170000000
0!
0%
#594175000000
1!
1%
#594180000000
0!
0%
#594185000000
1!
1%
#594190000000
0!
0%
#594195000000
1!
1%
#594200000000
0!
0%
#594205000000
1!
1%
#594210000000
0!
0%
#594215000000
1!
1%
#594220000000
0!
0%
#594225000000
1!
1%
#594230000000
0!
0%
#594235000000
1!
1%
#594240000000
0!
0%
#594245000000
1!
1%
#594250000000
0!
0%
#594255000000
1!
1%
#594260000000
0!
0%
#594265000000
1!
1%
#594270000000
0!
0%
#594275000000
1!
1%
#594280000000
0!
0%
#594285000000
1!
1%
#594290000000
0!
0%
#594295000000
1!
1%
#594300000000
0!
0%
#594305000000
1!
1%
#594310000000
0!
0%
#594315000000
1!
1%
#594320000000
0!
0%
#594325000000
1!
1%
#594330000000
0!
0%
#594335000000
1!
1%
#594340000000
0!
0%
#594345000000
1!
1%
#594350000000
0!
0%
#594355000000
1!
1%
#594360000000
0!
0%
#594365000000
1!
1%
#594370000000
0!
0%
#594375000000
1!
1%
#594380000000
0!
0%
#594385000000
1!
1%
#594390000000
0!
0%
#594395000000
1!
1%
#594400000000
0!
0%
#594405000000
1!
1%
#594410000000
0!
0%
#594415000000
1!
1%
#594420000000
0!
0%
#594425000000
1!
1%
#594430000000
0!
0%
#594435000000
1!
1%
#594440000000
0!
0%
#594445000000
1!
1%
#594450000000
0!
0%
#594455000000
1!
1%
#594460000000
0!
0%
#594465000000
1!
1%
#594470000000
0!
0%
#594475000000
1!
1%
#594480000000
0!
0%
#594485000000
1!
1%
#594490000000
0!
0%
#594495000000
1!
1%
#594500000000
0!
0%
#594505000000
1!
1%
#594510000000
0!
0%
#594515000000
1!
1%
#594520000000
0!
0%
#594525000000
1!
1%
#594530000000
0!
0%
#594535000000
1!
1%
#594540000000
0!
0%
#594545000000
1!
1%
#594550000000
0!
0%
#594555000000
1!
1%
#594560000000
0!
0%
#594565000000
1!
1%
#594570000000
0!
0%
#594575000000
1!
1%
#594580000000
0!
0%
#594585000000
1!
1%
#594590000000
0!
0%
#594595000000
1!
1%
#594600000000
0!
0%
#594605000000
1!
1%
#594610000000
0!
0%
#594615000000
1!
1%
#594620000000
0!
0%
#594625000000
1!
1%
#594630000000
0!
0%
#594635000000
1!
1%
#594640000000
0!
0%
#594645000000
1!
1%
#594650000000
0!
0%
#594655000000
1!
1%
#594660000000
0!
0%
#594665000000
1!
1%
#594670000000
0!
0%
#594675000000
1!
1%
#594680000000
0!
0%
#594685000000
1!
1%
#594690000000
0!
0%
#594695000000
1!
1%
#594700000000
0!
0%
#594705000000
1!
1%
#594710000000
0!
0%
#594715000000
1!
1%
#594720000000
0!
0%
#594725000000
1!
1%
#594730000000
0!
0%
#594735000000
1!
1%
#594740000000
0!
0%
#594745000000
1!
1%
#594750000000
0!
0%
#594755000000
1!
1%
#594760000000
0!
0%
#594765000000
1!
1%
#594770000000
0!
0%
#594775000000
1!
1%
#594780000000
0!
0%
#594785000000
1!
1%
#594790000000
0!
0%
#594795000000
1!
1%
#594800000000
0!
0%
#594805000000
1!
1%
#594810000000
0!
0%
#594815000000
1!
1%
#594820000000
0!
0%
#594825000000
1!
1%
#594830000000
0!
0%
#594835000000
1!
1%
#594840000000
0!
0%
#594845000000
1!
1%
#594850000000
0!
0%
#594855000000
1!
1%
#594860000000
0!
0%
#594865000000
1!
1%
#594870000000
0!
0%
#594875000000
1!
1%
#594880000000
0!
0%
#594885000000
1!
1%
#594890000000
0!
0%
#594895000000
1!
1%
#594900000000
0!
0%
#594905000000
1!
1%
#594910000000
0!
0%
#594915000000
1!
1%
#594920000000
0!
0%
#594925000000
1!
1%
#594930000000
0!
0%
#594935000000
1!
1%
#594940000000
0!
0%
#594945000000
1!
1%
#594950000000
0!
0%
#594955000000
1!
1%
#594960000000
0!
0%
#594965000000
1!
1%
#594970000000
0!
0%
#594975000000
1!
1%
#594980000000
0!
0%
#594985000000
1!
1%
#594990000000
0!
0%
#594995000000
1!
1%
#595000000000
0!
0%
#595005000000
1!
1%
#595010000000
0!
0%
#595015000000
1!
1%
#595020000000
0!
0%
#595025000000
1!
1%
#595030000000
0!
0%
#595035000000
1!
1%
#595040000000
0!
0%
#595045000000
1!
1%
#595050000000
0!
0%
#595055000000
1!
1%
#595060000000
0!
0%
#595065000000
1!
1%
#595070000000
0!
0%
#595075000000
1!
1%
#595080000000
0!
0%
#595085000000
1!
1%
#595090000000
0!
0%
#595095000000
1!
1%
#595100000000
0!
0%
#595105000000
1!
1%
#595110000000
0!
0%
#595115000000
1!
1%
#595120000000
0!
0%
#595125000000
1!
1%
#595130000000
0!
0%
#595135000000
1!
1%
#595140000000
0!
0%
#595145000000
1!
1%
#595150000000
0!
0%
#595155000000
1!
1%
#595160000000
0!
0%
#595165000000
1!
1%
#595170000000
0!
0%
#595175000000
1!
1%
#595180000000
0!
0%
#595185000000
1!
1%
#595190000000
0!
0%
#595195000000
1!
1%
#595200000000
0!
0%
#595205000000
1!
1%
#595210000000
0!
0%
#595215000000
1!
1%
#595220000000
0!
0%
#595225000000
1!
1%
#595230000000
0!
0%
#595235000000
1!
1%
#595240000000
0!
0%
#595245000000
1!
1%
#595250000000
0!
0%
#595255000000
1!
1%
#595260000000
0!
0%
#595265000000
1!
1%
#595270000000
0!
0%
#595275000000
1!
1%
#595280000000
0!
0%
#595285000000
1!
1%
#595290000000
0!
0%
#595295000000
1!
1%
#595300000000
0!
0%
#595305000000
1!
1%
#595310000000
0!
0%
#595315000000
1!
1%
#595320000000
0!
0%
#595325000000
1!
1%
#595330000000
0!
0%
#595335000000
1!
1%
#595340000000
0!
0%
#595345000000
1!
1%
#595350000000
0!
0%
#595355000000
1!
1%
#595360000000
0!
0%
#595365000000
1!
1%
#595370000000
0!
0%
#595375000000
1!
1%
#595380000000
0!
0%
#595385000000
1!
1%
#595390000000
0!
0%
#595395000000
1!
1%
#595400000000
0!
0%
#595405000000
1!
1%
#595410000000
0!
0%
#595415000000
1!
1%
#595420000000
0!
0%
#595425000000
1!
1%
#595430000000
0!
0%
#595435000000
1!
1%
#595440000000
0!
0%
#595445000000
1!
1%
#595450000000
0!
0%
#595455000000
1!
1%
#595460000000
0!
0%
#595465000000
1!
1%
#595470000000
0!
0%
#595475000000
1!
1%
#595480000000
0!
0%
#595485000000
1!
1%
#595490000000
0!
0%
#595495000000
1!
1%
#595500000000
0!
0%
#595505000000
1!
1%
#595510000000
0!
0%
#595515000000
1!
1%
#595520000000
0!
0%
#595525000000
1!
1%
#595530000000
0!
0%
#595535000000
1!
1%
#595540000000
0!
0%
#595545000000
1!
1%
#595550000000
0!
0%
#595555000000
1!
1%
#595560000000
0!
0%
#595565000000
1!
1%
#595570000000
0!
0%
#595575000000
1!
1%
#595580000000
0!
0%
#595585000000
1!
1%
#595590000000
0!
0%
#595595000000
1!
1%
#595600000000
0!
0%
#595605000000
1!
1%
#595610000000
0!
0%
#595615000000
1!
1%
#595620000000
0!
0%
#595625000000
1!
1%
#595630000000
0!
0%
#595635000000
1!
1%
#595640000000
0!
0%
#595645000000
1!
1%
#595650000000
0!
0%
#595655000000
1!
1%
#595660000000
0!
0%
#595665000000
1!
1%
#595670000000
0!
0%
#595675000000
1!
1%
#595680000000
0!
0%
#595685000000
1!
1%
#595690000000
0!
0%
#595695000000
1!
1%
#595700000000
0!
0%
#595705000000
1!
1%
#595710000000
0!
0%
#595715000000
1!
1%
#595720000000
0!
0%
#595725000000
1!
1%
#595730000000
0!
0%
#595735000000
1!
1%
#595740000000
0!
0%
#595745000000
1!
1%
#595750000000
0!
0%
#595755000000
1!
1%
#595760000000
0!
0%
#595765000000
1!
1%
#595770000000
0!
0%
#595775000000
1!
1%
#595780000000
0!
0%
#595785000000
1!
1%
#595790000000
0!
0%
#595795000000
1!
1%
#595800000000
0!
0%
#595805000000
1!
1%
#595810000000
0!
0%
#595815000000
1!
1%
#595820000000
0!
0%
#595825000000
1!
1%
#595830000000
0!
0%
#595835000000
1!
1%
#595840000000
0!
0%
#595845000000
1!
1%
#595850000000
0!
0%
#595855000000
1!
1%
#595860000000
0!
0%
#595865000000
1!
1%
#595870000000
0!
0%
#595875000000
1!
1%
#595880000000
0!
0%
#595885000000
1!
1%
#595890000000
0!
0%
#595895000000
1!
1%
#595900000000
0!
0%
#595905000000
1!
1%
#595910000000
0!
0%
#595915000000
1!
1%
#595920000000
0!
0%
#595925000000
1!
1%
#595930000000
0!
0%
#595935000000
1!
1%
#595940000000
0!
0%
#595945000000
1!
1%
#595950000000
0!
0%
#595955000000
1!
1%
#595960000000
0!
0%
#595965000000
1!
1%
#595970000000
0!
0%
#595975000000
1!
1%
#595980000000
0!
0%
#595985000000
1!
1%
#595990000000
0!
0%
#595995000000
1!
1%
#596000000000
0!
0%
#596005000000
1!
1%
#596010000000
0!
0%
#596015000000
1!
1%
#596020000000
0!
0%
#596025000000
1!
1%
#596030000000
0!
0%
#596035000000
1!
1%
#596040000000
0!
0%
#596045000000
1!
1%
#596050000000
0!
0%
#596055000000
1!
1%
#596060000000
0!
0%
#596065000000
1!
1%
#596070000000
0!
0%
#596075000000
1!
1%
#596080000000
0!
0%
#596085000000
1!
1%
#596090000000
0!
0%
#596095000000
1!
1%
#596100000000
0!
0%
#596105000000
1!
1%
#596110000000
0!
0%
#596115000000
1!
1%
#596120000000
0!
0%
#596125000000
1!
1%
#596130000000
0!
0%
#596135000000
1!
1%
#596140000000
0!
0%
#596145000000
1!
1%
#596150000000
0!
0%
#596155000000
1!
1%
#596160000000
0!
0%
#596165000000
1!
1%
#596170000000
0!
0%
#596175000000
1!
1%
#596180000000
0!
0%
#596185000000
1!
1%
#596190000000
0!
0%
#596195000000
1!
1%
#596200000000
0!
0%
#596205000000
1!
1%
#596210000000
0!
0%
#596215000000
1!
1%
#596220000000
0!
0%
#596225000000
1!
1%
#596230000000
0!
0%
#596235000000
1!
1%
#596240000000
0!
0%
#596245000000
1!
1%
#596250000000
0!
0%
#596255000000
1!
1%
#596260000000
0!
0%
#596265000000
1!
1%
#596270000000
0!
0%
#596275000000
1!
1%
#596280000000
0!
0%
#596285000000
1!
1%
#596290000000
0!
0%
#596295000000
1!
1%
#596300000000
0!
0%
#596305000000
1!
1%
#596310000000
0!
0%
#596315000000
1!
1%
#596320000000
0!
0%
#596325000000
1!
1%
#596330000000
0!
0%
#596335000000
1!
1%
#596340000000
0!
0%
#596345000000
1!
1%
#596350000000
0!
0%
#596355000000
1!
1%
#596360000000
0!
0%
#596365000000
1!
1%
#596370000000
0!
0%
#596375000000
1!
1%
#596380000000
0!
0%
#596385000000
1!
1%
#596390000000
0!
0%
#596395000000
1!
1%
#596400000000
0!
0%
#596405000000
1!
1%
#596410000000
0!
0%
#596415000000
1!
1%
#596420000000
0!
0%
#596425000000
1!
1%
#596430000000
0!
0%
#596435000000
1!
1%
#596440000000
0!
0%
#596445000000
1!
1%
#596450000000
0!
0%
#596455000000
1!
1%
#596460000000
0!
0%
#596465000000
1!
1%
#596470000000
0!
0%
#596475000000
1!
1%
#596480000000
0!
0%
#596485000000
1!
1%
#596490000000
0!
0%
#596495000000
1!
1%
#596500000000
0!
0%
#596505000000
1!
1%
#596510000000
0!
0%
#596515000000
1!
1%
#596520000000
0!
0%
#596525000000
1!
1%
#596530000000
0!
0%
#596535000000
1!
1%
#596540000000
0!
0%
#596545000000
1!
1%
#596550000000
0!
0%
#596555000000
1!
1%
#596560000000
0!
0%
#596565000000
1!
1%
#596570000000
0!
0%
#596575000000
1!
1%
#596580000000
0!
0%
#596585000000
1!
1%
#596590000000
0!
0%
#596595000000
1!
1%
#596600000000
0!
0%
#596605000000
1!
1%
#596610000000
0!
0%
#596615000000
1!
1%
#596620000000
0!
0%
#596625000000
1!
1%
#596630000000
0!
0%
#596635000000
1!
1%
#596640000000
0!
0%
#596645000000
1!
1%
#596650000000
0!
0%
#596655000000
1!
1%
#596660000000
0!
0%
#596665000000
1!
1%
#596670000000
0!
0%
#596675000000
1!
1%
#596680000000
0!
0%
#596685000000
1!
1%
#596690000000
0!
0%
#596695000000
1!
1%
#596700000000
0!
0%
#596705000000
1!
1%
#596710000000
0!
0%
#596715000000
1!
1%
#596720000000
0!
0%
#596725000000
1!
1%
#596730000000
0!
0%
#596735000000
1!
1%
#596740000000
0!
0%
#596745000000
1!
1%
#596750000000
0!
0%
#596755000000
1!
1%
#596760000000
0!
0%
#596765000000
1!
1%
#596770000000
0!
0%
#596775000000
1!
1%
#596780000000
0!
0%
#596785000000
1!
1%
#596790000000
0!
0%
#596795000000
1!
1%
#596800000000
0!
0%
#596805000000
1!
1%
#596810000000
0!
0%
#596815000000
1!
1%
#596820000000
0!
0%
#596825000000
1!
1%
#596830000000
0!
0%
#596835000000
1!
1%
#596840000000
0!
0%
#596845000000
1!
1%
#596850000000
0!
0%
#596855000000
1!
1%
#596860000000
0!
0%
#596865000000
1!
1%
#596870000000
0!
0%
#596875000000
1!
1%
#596880000000
0!
0%
#596885000000
1!
1%
#596890000000
0!
0%
#596895000000
1!
1%
#596900000000
0!
0%
#596905000000
1!
1%
#596910000000
0!
0%
#596915000000
1!
1%
#596920000000
0!
0%
#596925000000
1!
1%
#596930000000
0!
0%
#596935000000
1!
1%
#596940000000
0!
0%
#596945000000
1!
1%
#596950000000
0!
0%
#596955000000
1!
1%
#596960000000
0!
0%
#596965000000
1!
1%
#596970000000
0!
0%
#596975000000
1!
1%
#596980000000
0!
0%
#596985000000
1!
1%
#596990000000
0!
0%
#596995000000
1!
1%
#597000000000
0!
0%
#597005000000
1!
1%
#597010000000
0!
0%
#597015000000
1!
1%
#597020000000
0!
0%
#597025000000
1!
1%
#597030000000
0!
0%
#597035000000
1!
1%
#597040000000
0!
0%
#597045000000
1!
1%
#597050000000
0!
0%
#597055000000
1!
1%
#597060000000
0!
0%
#597065000000
1!
1%
#597070000000
0!
0%
#597075000000
1!
1%
#597080000000
0!
0%
#597085000000
1!
1%
#597090000000
0!
0%
#597095000000
1!
1%
#597100000000
0!
0%
#597105000000
1!
1%
#597110000000
0!
0%
#597115000000
1!
1%
#597120000000
0!
0%
#597125000000
1!
1%
#597130000000
0!
0%
#597135000000
1!
1%
#597140000000
0!
0%
#597145000000
1!
1%
#597150000000
0!
0%
#597155000000
1!
1%
#597160000000
0!
0%
#597165000000
1!
1%
#597170000000
0!
0%
#597175000000
1!
1%
#597180000000
0!
0%
#597185000000
1!
1%
#597190000000
0!
0%
#597195000000
1!
1%
#597200000000
0!
0%
#597205000000
1!
1%
#597210000000
0!
0%
#597215000000
1!
1%
#597220000000
0!
0%
#597225000000
1!
1%
#597230000000
0!
0%
#597235000000
1!
1%
#597240000000
0!
0%
#597245000000
1!
1%
#597250000000
0!
0%
#597255000000
1!
1%
#597260000000
0!
0%
#597265000000
1!
1%
#597270000000
0!
0%
#597275000000
1!
1%
#597280000000
0!
0%
#597285000000
1!
1%
#597290000000
0!
0%
#597295000000
1!
1%
#597300000000
0!
0%
#597305000000
1!
1%
#597310000000
0!
0%
#597315000000
1!
1%
#597320000000
0!
0%
#597325000000
1!
1%
#597330000000
0!
0%
#597335000000
1!
1%
#597340000000
0!
0%
#597345000000
1!
1%
#597350000000
0!
0%
#597355000000
1!
1%
#597360000000
0!
0%
#597365000000
1!
1%
#597370000000
0!
0%
#597375000000
1!
1%
#597380000000
0!
0%
#597385000000
1!
1%
#597390000000
0!
0%
#597395000000
1!
1%
#597400000000
0!
0%
#597405000000
1!
1%
#597410000000
0!
0%
#597415000000
1!
1%
#597420000000
0!
0%
#597425000000
1!
1%
#597430000000
0!
0%
#597435000000
1!
1%
#597440000000
0!
0%
#597445000000
1!
1%
#597450000000
0!
0%
#597455000000
1!
1%
#597460000000
0!
0%
#597465000000
1!
1%
#597470000000
0!
0%
#597475000000
1!
1%
#597480000000
0!
0%
#597485000000
1!
1%
#597490000000
0!
0%
#597495000000
1!
1%
#597500000000
0!
0%
#597505000000
1!
1%
#597510000000
0!
0%
#597515000000
1!
1%
#597520000000
0!
0%
#597525000000
1!
1%
#597530000000
0!
0%
#597535000000
1!
1%
#597540000000
0!
0%
#597545000000
1!
1%
#597550000000
0!
0%
#597555000000
1!
1%
#597560000000
0!
0%
#597565000000
1!
1%
#597570000000
0!
0%
#597575000000
1!
1%
#597580000000
0!
0%
#597585000000
1!
1%
#597590000000
0!
0%
#597595000000
1!
1%
#597600000000
0!
0%
#597605000000
1!
1%
#597610000000
0!
0%
#597615000000
1!
1%
#597620000000
0!
0%
#597625000000
1!
1%
#597630000000
0!
0%
#597635000000
1!
1%
#597640000000
0!
0%
#597645000000
1!
1%
#597650000000
0!
0%
#597655000000
1!
1%
#597660000000
0!
0%
#597665000000
1!
1%
#597670000000
0!
0%
#597675000000
1!
1%
#597680000000
0!
0%
#597685000000
1!
1%
#597690000000
0!
0%
#597695000000
1!
1%
#597700000000
0!
0%
#597705000000
1!
1%
#597710000000
0!
0%
#597715000000
1!
1%
#597720000000
0!
0%
#597725000000
1!
1%
#597730000000
0!
0%
#597735000000
1!
1%
#597740000000
0!
0%
#597745000000
1!
1%
#597750000000
0!
0%
#597755000000
1!
1%
#597760000000
0!
0%
#597765000000
1!
1%
#597770000000
0!
0%
#597775000000
1!
1%
#597780000000
0!
0%
#597785000000
1!
1%
#597790000000
0!
0%
#597795000000
1!
1%
#597800000000
0!
0%
#597805000000
1!
1%
#597810000000
0!
0%
#597815000000
1!
1%
#597820000000
0!
0%
#597825000000
1!
1%
#597830000000
0!
0%
#597835000000
1!
1%
#597840000000
0!
0%
#597845000000
1!
1%
#597850000000
0!
0%
#597855000000
1!
1%
#597860000000
0!
0%
#597865000000
1!
1%
#597870000000
0!
0%
#597875000000
1!
1%
#597880000000
0!
0%
#597885000000
1!
1%
#597890000000
0!
0%
#597895000000
1!
1%
#597900000000
0!
0%
#597905000000
1!
1%
#597910000000
0!
0%
#597915000000
1!
1%
#597920000000
0!
0%
#597925000000
1!
1%
#597930000000
0!
0%
#597935000000
1!
1%
#597940000000
0!
0%
#597945000000
1!
1%
#597950000000
0!
0%
#597955000000
1!
1%
#597960000000
0!
0%
#597965000000
1!
1%
#597970000000
0!
0%
#597975000000
1!
1%
#597980000000
0!
0%
#597985000000
1!
1%
#597990000000
0!
0%
#597995000000
1!
1%
#598000000000
0!
0%
#598005000000
1!
1%
#598010000000
0!
0%
#598015000000
1!
1%
#598020000000
0!
0%
#598025000000
1!
1%
#598030000000
0!
0%
#598035000000
1!
1%
#598040000000
0!
0%
#598045000000
1!
1%
#598050000000
0!
0%
#598055000000
1!
1%
#598060000000
0!
0%
#598065000000
1!
1%
#598070000000
0!
0%
#598075000000
1!
1%
#598080000000
0!
0%
#598085000000
1!
1%
#598090000000
0!
0%
#598095000000
1!
1%
#598100000000
0!
0%
#598105000000
1!
1%
#598110000000
0!
0%
#598115000000
1!
1%
#598120000000
0!
0%
#598125000000
1!
1%
#598130000000
0!
0%
#598135000000
1!
1%
#598140000000
0!
0%
#598145000000
1!
1%
#598150000000
0!
0%
#598155000000
1!
1%
#598160000000
0!
0%
#598165000000
1!
1%
#598170000000
0!
0%
#598175000000
1!
1%
#598180000000
0!
0%
#598185000000
1!
1%
#598190000000
0!
0%
#598195000000
1!
1%
#598200000000
0!
0%
#598205000000
1!
1%
#598210000000
0!
0%
#598215000000
1!
1%
#598220000000
0!
0%
#598225000000
1!
1%
#598230000000
0!
0%
#598235000000
1!
1%
#598240000000
0!
0%
#598245000000
1!
1%
#598250000000
0!
0%
#598255000000
1!
1%
#598260000000
0!
0%
#598265000000
1!
1%
#598270000000
0!
0%
#598275000000
1!
1%
#598280000000
0!
0%
#598285000000
1!
1%
#598290000000
0!
0%
#598295000000
1!
1%
#598300000000
0!
0%
#598305000000
1!
1%
#598310000000
0!
0%
#598315000000
1!
1%
#598320000000
0!
0%
#598325000000
1!
1%
#598330000000
0!
0%
#598335000000
1!
1%
#598340000000
0!
0%
#598345000000
1!
1%
#598350000000
0!
0%
#598355000000
1!
1%
#598360000000
0!
0%
#598365000000
1!
1%
#598370000000
0!
0%
#598375000000
1!
1%
#598380000000
0!
0%
#598385000000
1!
1%
#598390000000
0!
0%
#598395000000
1!
1%
#598400000000
0!
0%
#598405000000
1!
1%
#598410000000
0!
0%
#598415000000
1!
1%
#598420000000
0!
0%
#598425000000
1!
1%
#598430000000
0!
0%
#598435000000
1!
1%
#598440000000
0!
0%
#598445000000
1!
1%
#598450000000
0!
0%
#598455000000
1!
1%
#598460000000
0!
0%
#598465000000
1!
1%
#598470000000
0!
0%
#598475000000
1!
1%
#598480000000
0!
0%
#598485000000
1!
1%
#598490000000
0!
0%
#598495000000
1!
1%
#598500000000
0!
0%
#598505000000
1!
1%
#598510000000
0!
0%
#598515000000
1!
1%
#598520000000
0!
0%
#598525000000
1!
1%
#598530000000
0!
0%
#598535000000
1!
1%
#598540000000
0!
0%
#598545000000
1!
1%
#598550000000
0!
0%
#598555000000
1!
1%
#598560000000
0!
0%
#598565000000
1!
1%
#598570000000
0!
0%
#598575000000
1!
1%
#598580000000
0!
0%
#598585000000
1!
1%
#598590000000
0!
0%
#598595000000
1!
1%
#598600000000
0!
0%
#598605000000
1!
1%
#598610000000
0!
0%
#598615000000
1!
1%
#598620000000
0!
0%
#598625000000
1!
1%
#598630000000
0!
0%
#598635000000
1!
1%
#598640000000
0!
0%
#598645000000
1!
1%
#598650000000
0!
0%
#598655000000
1!
1%
#598660000000
0!
0%
#598665000000
1!
1%
#598670000000
0!
0%
#598675000000
1!
1%
#598680000000
0!
0%
#598685000000
1!
1%
#598690000000
0!
0%
#598695000000
1!
1%
#598700000000
0!
0%
#598705000000
1!
1%
#598710000000
0!
0%
#598715000000
1!
1%
#598720000000
0!
0%
#598725000000
1!
1%
#598730000000
0!
0%
#598735000000
1!
1%
#598740000000
0!
0%
#598745000000
1!
1%
#598750000000
0!
0%
#598755000000
1!
1%
#598760000000
0!
0%
#598765000000
1!
1%
#598770000000
0!
0%
#598775000000
1!
1%
#598780000000
0!
0%
#598785000000
1!
1%
#598790000000
0!
0%
#598795000000
1!
1%
#598800000000
0!
0%
#598805000000
1!
1%
#598810000000
0!
0%
#598815000000
1!
1%
#598820000000
0!
0%
#598825000000
1!
1%
#598830000000
0!
0%
#598835000000
1!
1%
#598840000000
0!
0%
#598845000000
1!
1%
#598850000000
0!
0%
#598855000000
1!
1%
#598860000000
0!
0%
#598865000000
1!
1%
#598870000000
0!
0%
#598875000000
1!
1%
#598880000000
0!
0%
#598885000000
1!
1%
#598890000000
0!
0%
#598895000000
1!
1%
#598900000000
0!
0%
#598905000000
1!
1%
#598910000000
0!
0%
#598915000000
1!
1%
#598920000000
0!
0%
#598925000000
1!
1%
#598930000000
0!
0%
#598935000000
1!
1%
#598940000000
0!
0%
#598945000000
1!
1%
#598950000000
0!
0%
#598955000000
1!
1%
#598960000000
0!
0%
#598965000000
1!
1%
#598970000000
0!
0%
#598975000000
1!
1%
#598980000000
0!
0%
#598985000000
1!
1%
#598990000000
0!
0%
#598995000000
1!
1%
#599000000000
0!
0%
#599005000000
1!
1%
#599010000000
0!
0%
#599015000000
1!
1%
#599020000000
0!
0%
#599025000000
1!
1%
#599030000000
0!
0%
#599035000000
1!
1%
#599040000000
0!
0%
#599045000000
1!
1%
#599050000000
0!
0%
#599055000000
1!
1%
#599060000000
0!
0%
#599065000000
1!
1%
#599070000000
0!
0%
#599075000000
1!
1%
#599080000000
0!
0%
#599085000000
1!
1%
#599090000000
0!
0%
#599095000000
1!
1%
#599100000000
0!
0%
#599105000000
1!
1%
#599110000000
0!
0%
#599115000000
1!
1%
#599120000000
0!
0%
#599125000000
1!
1%
#599130000000
0!
0%
#599135000000
1!
1%
#599140000000
0!
0%
#599145000000
1!
1%
#599150000000
0!
0%
#599155000000
1!
1%
#599160000000
0!
0%
#599165000000
1!
1%
#599170000000
0!
0%
#599175000000
1!
1%
#599180000000
0!
0%
#599185000000
1!
1%
#599190000000
0!
0%
#599195000000
1!
1%
#599200000000
0!
0%
#599205000000
1!
1%
#599210000000
0!
0%
#599215000000
1!
1%
#599220000000
0!
0%
#599225000000
1!
1%
#599230000000
0!
0%
#599235000000
1!
1%
#599240000000
0!
0%
#599245000000
1!
1%
#599250000000
0!
0%
#599255000000
1!
1%
#599260000000
0!
0%
#599265000000
1!
1%
#599270000000
0!
0%
#599275000000
1!
1%
#599280000000
0!
0%
#599285000000
1!
1%
#599290000000
0!
0%
#599295000000
1!
1%
#599300000000
0!
0%
#599305000000
1!
1%
#599310000000
0!
0%
#599315000000
1!
1%
#599320000000
0!
0%
#599325000000
1!
1%
#599330000000
0!
0%
#599335000000
1!
1%
#599340000000
0!
0%
#599345000000
1!
1%
#599350000000
0!
0%
#599355000000
1!
1%
#599360000000
0!
0%
#599365000000
1!
1%
#599370000000
0!
0%
#599375000000
1!
1%
#599380000000
0!
0%
#599385000000
1!
1%
#599390000000
0!
0%
#599395000000
1!
1%
#599400000000
0!
0%
#599405000000
1!
1%
#599410000000
0!
0%
#599415000000
1!
1%
#599420000000
0!
0%
#599425000000
1!
1%
#599430000000
0!
0%
#599435000000
1!
1%
#599440000000
0!
0%
#599445000000
1!
1%
#599450000000
0!
0%
#599455000000
1!
1%
#599460000000
0!
0%
#599465000000
1!
1%
#599470000000
0!
0%
#599475000000
1!
1%
#599480000000
0!
0%
#599485000000
1!
1%
#599490000000
0!
0%
#599495000000
1!
1%
#599500000000
0!
0%
#599505000000
1!
1%
#599510000000
0!
0%
#599515000000
1!
1%
#599520000000
0!
0%
#599525000000
1!
1%
#599530000000
0!
0%
#599535000000
1!
1%
#599540000000
0!
0%
#599545000000
1!
1%
#599550000000
0!
0%
#599555000000
1!
1%
#599560000000
0!
0%
#599565000000
1!
1%
#599570000000
0!
0%
#599575000000
1!
1%
#599580000000
0!
0%
#599585000000
1!
1%
#599590000000
0!
0%
#599595000000
1!
1%
#599600000000
0!
0%
#599605000000
1!
1%
#599610000000
0!
0%
#599615000000
1!
1%
#599620000000
0!
0%
#599625000000
1!
1%
#599630000000
0!
0%
#599635000000
1!
1%
#599640000000
0!
0%
#599645000000
1!
1%
#599650000000
0!
0%
#599655000000
1!
1%
#599660000000
0!
0%
#599665000000
1!
1%
#599670000000
0!
0%
#599675000000
1!
1%
#599680000000
0!
0%
#599685000000
1!
1%
#599690000000
0!
0%
#599695000000
1!
1%
#599700000000
0!
0%
#599705000000
1!
1%
#599710000000
0!
0%
#599715000000
1!
1%
#599720000000
0!
0%
#599725000000
1!
1%
#599730000000
0!
0%
#599735000000
1!
1%
#599740000000
0!
0%
#599745000000
1!
1%
#599750000000
0!
0%
#599755000000
1!
1%
#599760000000
0!
0%
#599765000000
1!
1%
#599770000000
0!
0%
#599775000000
1!
1%
#599780000000
0!
0%
#599785000000
1!
1%
#599790000000
0!
0%
#599795000000
1!
1%
#599800000000
0!
0%
#599805000000
1!
1%
#599810000000
0!
0%
#599815000000
1!
1%
#599820000000
0!
0%
#599825000000
1!
1%
#599830000000
0!
0%
#599835000000
1!
1%
#599840000000
0!
0%
#599845000000
1!
1%
#599850000000
0!
0%
#599855000000
1!
1%
#599860000000
0!
0%
#599865000000
1!
1%
#599870000000
0!
0%
#599875000000
1!
1%
#599880000000
0!
0%
#599885000000
1!
1%
#599890000000
0!
0%
#599895000000
1!
1%
#599900000000
0!
0%
#599905000000
1!
1%
#599910000000
0!
0%
#599915000000
1!
1%
#599920000000
0!
0%
#599925000000
1!
1%
#599930000000
0!
0%
#599935000000
1!
1%
#599940000000
0!
0%
#599945000000
1!
1%
#599950000000
0!
0%
#599955000000
1!
1%
#599960000000
0!
0%
#599965000000
1!
1%
#599970000000
0!
0%
#599975000000
1!
1%
#599980000000
0!
0%
#599985000000
1!
1%
#599990000000
0!
0%
#599995000000
1!
1%
#600000000000
0!
0%
#600005000000
1!
1%
#600010000000
0!
0%
#600015000000
1!
1%
#600020000000
0!
0%
#600025000000
1!
1%
#600030000000
0!
0%
#600035000000
1!
1%
#600040000000
0!
0%
#600045000000
1!
1%
#600050000000
0!
0%
#600055000000
1!
1%
#600060000000
0!
0%
#600065000000
1!
1%
#600070000000
0!
0%
#600075000000
1!
1%
#600080000000
0!
0%
#600085000000
1!
1%
#600090000000
0!
0%
#600095000000
1!
1%
#600100000000
0!
0%
#600105000000
1!
1%
#600110000000
0!
0%
#600115000000
1!
1%
#600120000000
0!
0%
#600125000000
1!
1%
#600130000000
0!
0%
#600135000000
1!
1%
#600140000000
0!
0%
#600145000000
1!
1%
#600150000000
0!
0%
#600155000000
1!
1%
#600160000000
0!
0%
#600165000000
1!
1%
#600170000000
0!
0%
#600175000000
1!
1%
#600180000000
0!
0%
#600185000000
1!
1%
#600190000000
0!
0%
#600195000000
1!
1%
#600200000000
0!
0%
#600205000000
1!
1%
#600210000000
0!
0%
#600215000000
1!
1%
#600220000000
0!
0%
#600225000000
1!
1%
#600230000000
0!
0%
#600235000000
1!
1%
#600240000000
0!
0%
#600245000000
1!
1%
#600250000000
0!
0%
#600255000000
1!
1%
#600260000000
0!
0%
#600265000000
1!
1%
#600270000000
0!
0%
#600275000000
1!
1%
#600280000000
0!
0%
#600285000000
1!
1%
#600290000000
0!
0%
#600295000000
1!
1%
#600300000000
0!
0%
#600305000000
1!
1%
#600310000000
0!
0%
#600315000000
1!
1%
#600320000000
0!
0%
#600325000000
1!
1%
#600330000000
0!
0%
#600335000000
1!
1%
#600340000000
0!
0%
#600345000000
1!
1%
#600350000000
0!
0%
#600355000000
1!
1%
#600360000000
0!
0%
#600365000000
1!
1%
#600370000000
0!
0%
#600375000000
1!
1%
#600380000000
0!
0%
#600385000000
1!
1%
#600390000000
0!
0%
#600395000000
1!
1%
#600400000000
0!
0%
#600405000000
1!
1%
#600410000000
0!
0%
#600415000000
1!
1%
#600420000000
0!
0%
#600425000000
1!
1%
#600430000000
0!
0%
#600435000000
1!
1%
#600440000000
0!
0%
#600445000000
1!
1%
#600450000000
0!
0%
#600455000000
1!
1%
#600460000000
0!
0%
#600465000000
1!
1%
#600470000000
0!
0%
#600475000000
1!
1%
#600480000000
0!
0%
#600485000000
1!
1%
#600490000000
0!
0%
#600495000000
1!
1%
#600500000000
0!
0%
#600505000000
1!
1%
#600510000000
0!
0%
#600515000000
1!
1%
#600520000000
0!
0%
#600525000000
1!
1%
#600530000000
0!
0%
#600535000000
1!
1%
#600540000000
0!
0%
#600545000000
1!
1%
#600550000000
0!
0%
#600555000000
1!
1%
#600560000000
0!
0%
#600565000000
1!
1%
#600570000000
0!
0%
#600575000000
1!
1%
#600580000000
0!
0%
#600585000000
1!
1%
#600590000000
0!
0%
#600595000000
1!
1%
#600600000000
0!
0%
#600605000000
1!
1%
#600610000000
0!
0%
#600615000000
1!
1%
#600620000000
0!
0%
#600625000000
1!
1%
#600630000000
0!
0%
#600635000000
1!
1%
#600640000000
0!
0%
#600645000000
1!
1%
#600650000000
0!
0%
#600655000000
1!
1%
#600660000000
0!
0%
#600665000000
1!
1%
#600670000000
0!
0%
#600675000000
1!
1%
#600680000000
0!
0%
#600685000000
1!
1%
#600690000000
0!
0%
#600695000000
1!
1%
#600700000000
0!
0%
#600705000000
1!
1%
#600710000000
0!
0%
#600715000000
1!
1%
#600720000000
0!
0%
#600725000000
1!
1%
#600730000000
0!
0%
#600735000000
1!
1%
#600740000000
0!
0%
#600745000000
1!
1%
#600750000000
0!
0%
#600755000000
1!
1%
#600760000000
0!
0%
#600765000000
1!
1%
#600770000000
0!
0%
#600775000000
1!
1%
#600780000000
0!
0%
#600785000000
1!
1%
#600790000000
0!
0%
#600795000000
1!
1%
#600800000000
0!
0%
#600805000000
1!
1%
#600810000000
0!
0%
#600815000000
1!
1%
#600820000000
0!
0%
#600825000000
1!
1%
#600830000000
0!
0%
#600835000000
1!
1%
#600840000000
0!
0%
#600845000000
1!
1%
#600850000000
0!
0%
#600855000000
1!
1%
#600860000000
0!
0%
#600865000000
1!
1%
#600870000000
0!
0%
#600875000000
1!
1%
#600880000000
0!
0%
#600885000000
1!
1%
#600890000000
0!
0%
#600895000000
1!
1%
#600900000000
0!
0%
#600905000000
1!
1%
#600910000000
0!
0%
#600915000000
1!
1%
#600920000000
0!
0%
#600925000000
1!
1%
#600930000000
0!
0%
#600935000000
1!
1%
#600940000000
0!
0%
#600945000000
1!
1%
#600950000000
0!
0%
#600955000000
1!
1%
#600960000000
0!
0%
#600965000000
1!
1%
#600970000000
0!
0%
#600975000000
1!
1%
#600980000000
0!
0%
#600985000000
1!
1%
#600990000000
0!
0%
#600995000000
1!
1%
#601000000000
0!
0%
#601005000000
1!
1%
#601010000000
0!
0%
#601015000000
1!
1%
#601020000000
0!
0%
#601025000000
1!
1%
#601030000000
0!
0%
#601035000000
1!
1%
#601040000000
0!
0%
#601045000000
1!
1%
#601050000000
0!
0%
#601055000000
1!
1%
#601060000000
0!
0%
#601065000000
1!
1%
#601070000000
0!
0%
#601075000000
1!
1%
#601080000000
0!
0%
#601085000000
1!
1%
#601090000000
0!
0%
#601095000000
1!
1%
#601100000000
0!
0%
#601105000000
1!
1%
#601110000000
0!
0%
#601115000000
1!
1%
#601120000000
0!
0%
#601125000000
1!
1%
#601130000000
0!
0%
#601135000000
1!
1%
#601140000000
0!
0%
#601145000000
1!
1%
#601150000000
0!
0%
#601155000000
1!
1%
#601160000000
0!
0%
#601165000000
1!
1%
#601170000000
0!
0%
#601175000000
1!
1%
#601180000000
0!
0%
#601185000000
1!
1%
#601190000000
0!
0%
#601195000000
1!
1%
#601200000000
0!
0%
#601205000000
1!
1%
#601210000000
0!
0%
#601215000000
1!
1%
#601220000000
0!
0%
#601225000000
1!
1%
#601230000000
0!
0%
#601235000000
1!
1%
#601240000000
0!
0%
#601245000000
1!
1%
#601250000000
0!
0%
#601255000000
1!
1%
#601260000000
0!
0%
#601265000000
1!
1%
#601270000000
0!
0%
#601275000000
1!
1%
#601280000000
0!
0%
#601285000000
1!
1%
#601290000000
0!
0%
#601295000000
1!
1%
#601300000000
0!
0%
#601305000000
1!
1%
#601310000000
0!
0%
#601315000000
1!
1%
#601320000000
0!
0%
#601325000000
1!
1%
#601330000000
0!
0%
#601335000000
1!
1%
#601340000000
0!
0%
#601345000000
1!
1%
#601350000000
0!
0%
#601355000000
1!
1%
#601360000000
0!
0%
#601365000000
1!
1%
#601370000000
0!
0%
#601375000000
1!
1%
#601380000000
0!
0%
#601385000000
1!
1%
#601390000000
0!
0%
#601395000000
1!
1%
#601400000000
0!
0%
#601405000000
1!
1%
#601410000000
0!
0%
#601415000000
1!
1%
#601420000000
0!
0%
#601425000000
1!
1%
#601430000000
0!
0%
#601435000000
1!
1%
#601440000000
0!
0%
#601445000000
1!
1%
#601450000000
0!
0%
#601455000000
1!
1%
#601460000000
0!
0%
#601465000000
1!
1%
#601470000000
0!
0%
#601475000000
1!
1%
#601480000000
0!
0%
#601485000000
1!
1%
#601490000000
0!
0%
#601495000000
1!
1%
#601500000000
0!
0%
#601505000000
1!
1%
#601510000000
0!
0%
#601515000000
1!
1%
#601520000000
0!
0%
#601525000000
1!
1%
#601530000000
0!
0%
#601535000000
1!
1%
#601540000000
0!
0%
#601545000000
1!
1%
#601550000000
0!
0%
#601555000000
1!
1%
#601560000000
0!
0%
#601565000000
1!
1%
#601570000000
0!
0%
#601575000000
1!
1%
#601580000000
0!
0%
#601585000000
1!
1%
#601590000000
0!
0%
#601595000000
1!
1%
#601600000000
0!
0%
#601605000000
1!
1%
#601610000000
0!
0%
#601615000000
1!
1%
#601620000000
0!
0%
#601625000000
1!
1%
#601630000000
0!
0%
#601635000000
1!
1%
#601640000000
0!
0%
#601645000000
1!
1%
#601650000000
0!
0%
#601655000000
1!
1%
#601660000000
0!
0%
#601665000000
1!
1%
#601670000000
0!
0%
#601675000000
1!
1%
#601680000000
0!
0%
#601685000000
1!
1%
#601690000000
0!
0%
#601695000000
1!
1%
#601700000000
0!
0%
#601705000000
1!
1%
#601710000000
0!
0%
#601715000000
1!
1%
#601720000000
0!
0%
#601725000000
1!
1%
#601730000000
0!
0%
#601735000000
1!
1%
#601740000000
0!
0%
#601745000000
1!
1%
#601750000000
0!
0%
#601755000000
1!
1%
#601760000000
0!
0%
#601765000000
1!
1%
#601770000000
0!
0%
#601775000000
1!
1%
#601780000000
0!
0%
#601785000000
1!
1%
#601790000000
0!
0%
#601795000000
1!
1%
#601800000000
0!
0%
#601805000000
1!
1%
#601810000000
0!
0%
#601815000000
1!
1%
#601820000000
0!
0%
#601825000000
1!
1%
#601830000000
0!
0%
#601835000000
1!
1%
#601840000000
0!
0%
#601845000000
1!
1%
#601850000000
0!
0%
#601855000000
1!
1%
#601860000000
0!
0%
#601865000000
1!
1%
#601870000000
0!
0%
#601875000000
1!
1%
#601880000000
0!
0%
#601885000000
1!
1%
#601890000000
0!
0%
#601895000000
1!
1%
#601900000000
0!
0%
#601905000000
1!
1%
#601910000000
0!
0%
#601915000000
1!
1%
#601920000000
0!
0%
#601925000000
1!
1%
#601930000000
0!
0%
#601935000000
1!
1%
#601940000000
0!
0%
#601945000000
1!
1%
#601950000000
0!
0%
#601955000000
1!
1%
#601960000000
0!
0%
#601965000000
1!
1%
#601970000000
0!
0%
#601975000000
1!
1%
#601980000000
0!
0%
#601985000000
1!
1%
#601990000000
0!
0%
#601995000000
1!
1%
#602000000000
0!
0%
#602005000000
1!
1%
#602010000000
0!
0%
#602015000000
1!
1%
#602020000000
0!
0%
#602025000000
1!
1%
#602030000000
0!
0%
#602035000000
1!
1%
#602040000000
0!
0%
#602045000000
1!
1%
#602050000000
0!
0%
#602055000000
1!
1%
#602060000000
0!
0%
#602065000000
1!
1%
#602070000000
0!
0%
#602075000000
1!
1%
#602080000000
0!
0%
#602085000000
1!
1%
#602090000000
0!
0%
#602095000000
1!
1%
#602100000000
0!
0%
#602105000000
1!
1%
#602110000000
0!
0%
#602115000000
1!
1%
#602120000000
0!
0%
#602125000000
1!
1%
#602130000000
0!
0%
#602135000000
1!
1%
#602140000000
0!
0%
#602145000000
1!
1%
#602150000000
0!
0%
#602155000000
1!
1%
#602160000000
0!
0%
#602165000000
1!
1%
#602170000000
0!
0%
#602175000000
1!
1%
#602180000000
0!
0%
#602185000000
1!
1%
#602190000000
0!
0%
#602195000000
1!
1%
#602200000000
0!
0%
#602205000000
1!
1%
#602210000000
0!
0%
#602215000000
1!
1%
#602220000000
0!
0%
#602225000000
1!
1%
#602230000000
0!
0%
#602235000000
1!
1%
#602240000000
0!
0%
#602245000000
1!
1%
#602250000000
0!
0%
#602255000000
1!
1%
#602260000000
0!
0%
#602265000000
1!
1%
#602270000000
0!
0%
#602275000000
1!
1%
#602280000000
0!
0%
#602285000000
1!
1%
#602290000000
0!
0%
#602295000000
1!
1%
#602300000000
0!
0%
#602305000000
1!
1%
#602310000000
0!
0%
#602315000000
1!
1%
#602320000000
0!
0%
#602325000000
1!
1%
#602330000000
0!
0%
#602335000000
1!
1%
#602340000000
0!
0%
#602345000000
1!
1%
#602350000000
0!
0%
#602355000000
1!
1%
#602360000000
0!
0%
#602365000000
1!
1%
#602370000000
0!
0%
#602375000000
1!
1%
#602380000000
0!
0%
#602385000000
1!
1%
#602390000000
0!
0%
#602395000000
1!
1%
#602400000000
0!
0%
#602405000000
1!
1%
#602410000000
0!
0%
#602415000000
1!
1%
#602420000000
0!
0%
#602425000000
1!
1%
#602430000000
0!
0%
#602435000000
1!
1%
#602440000000
0!
0%
#602445000000
1!
1%
#602450000000
0!
0%
#602455000000
1!
1%
#602460000000
0!
0%
#602465000000
1!
1%
#602470000000
0!
0%
#602475000000
1!
1%
#602480000000
0!
0%
#602485000000
1!
1%
#602490000000
0!
0%
#602495000000
1!
1%
#602500000000
0!
0%
#602505000000
1!
1%
#602510000000
0!
0%
#602515000000
1!
1%
#602520000000
0!
0%
#602525000000
1!
1%
#602530000000
0!
0%
#602535000000
1!
1%
#602540000000
0!
0%
#602545000000
1!
1%
#602550000000
0!
0%
#602555000000
1!
1%
#602560000000
0!
0%
#602565000000
1!
1%
#602570000000
0!
0%
#602575000000
1!
1%
#602580000000
0!
0%
#602585000000
1!
1%
#602590000000
0!
0%
#602595000000
1!
1%
#602600000000
0!
0%
#602605000000
1!
1%
#602610000000
0!
0%
#602615000000
1!
1%
#602620000000
0!
0%
#602625000000
1!
1%
#602630000000
0!
0%
#602635000000
1!
1%
#602640000000
0!
0%
#602645000000
1!
1%
#602650000000
0!
0%
#602655000000
1!
1%
#602660000000
0!
0%
#602665000000
1!
1%
#602670000000
0!
0%
#602675000000
1!
1%
#602680000000
0!
0%
#602685000000
1!
1%
#602690000000
0!
0%
#602695000000
1!
1%
#602700000000
0!
0%
#602705000000
1!
1%
#602710000000
0!
0%
#602715000000
1!
1%
#602720000000
0!
0%
#602725000000
1!
1%
#602730000000
0!
0%
#602735000000
1!
1%
#602740000000
0!
0%
#602745000000
1!
1%
#602750000000
0!
0%
#602755000000
1!
1%
#602760000000
0!
0%
#602765000000
1!
1%
#602770000000
0!
0%
#602775000000
1!
1%
#602780000000
0!
0%
#602785000000
1!
1%
#602790000000
0!
0%
#602795000000
1!
1%
#602800000000
0!
0%
#602805000000
1!
1%
#602810000000
0!
0%
#602815000000
1!
1%
#602820000000
0!
0%
#602825000000
1!
1%
#602830000000
0!
0%
#602835000000
1!
1%
#602840000000
0!
0%
#602845000000
1!
1%
#602850000000
0!
0%
#602855000000
1!
1%
#602860000000
0!
0%
#602865000000
1!
1%
#602870000000
0!
0%
#602875000000
1!
1%
#602880000000
0!
0%
#602885000000
1!
1%
#602890000000
0!
0%
#602895000000
1!
1%
#602900000000
0!
0%
#602905000000
1!
1%
#602910000000
0!
0%
#602915000000
1!
1%
#602920000000
0!
0%
#602925000000
1!
1%
#602930000000
0!
0%
#602935000000
1!
1%
#602940000000
0!
0%
#602945000000
1!
1%
#602950000000
0!
0%
#602955000000
1!
1%
#602960000000
0!
0%
#602965000000
1!
1%
#602970000000
0!
0%
#602975000000
1!
1%
#602980000000
0!
0%
#602985000000
1!
1%
#602990000000
0!
0%
#602995000000
1!
1%
#603000000000
0!
0%
#603005000000
1!
1%
#603010000000
0!
0%
#603015000000
1!
1%
#603020000000
0!
0%
#603025000000
1!
1%
#603030000000
0!
0%
#603035000000
1!
1%
#603040000000
0!
0%
#603045000000
1!
1%
#603050000000
0!
0%
#603055000000
1!
1%
#603060000000
0!
0%
#603065000000
1!
1%
#603070000000
0!
0%
#603075000000
1!
1%
#603080000000
0!
0%
#603085000000
1!
1%
#603090000000
0!
0%
#603095000000
1!
1%
#603100000000
0!
0%
#603105000000
1!
1%
#603110000000
0!
0%
#603115000000
1!
1%
#603120000000
0!
0%
#603125000000
1!
1%
#603130000000
0!
0%
#603135000000
1!
1%
#603140000000
0!
0%
#603145000000
1!
1%
#603150000000
0!
0%
#603155000000
1!
1%
#603160000000
0!
0%
#603165000000
1!
1%
#603170000000
0!
0%
#603175000000
1!
1%
#603180000000
0!
0%
#603185000000
1!
1%
#603190000000
0!
0%
#603195000000
1!
1%
#603200000000
0!
0%
#603205000000
1!
1%
#603210000000
0!
0%
#603215000000
1!
1%
#603220000000
0!
0%
#603225000000
1!
1%
#603230000000
0!
0%
#603235000000
1!
1%
#603240000000
0!
0%
#603245000000
1!
1%
#603250000000
0!
0%
#603255000000
1!
1%
#603260000000
0!
0%
#603265000000
1!
1%
#603270000000
0!
0%
#603275000000
1!
1%
#603280000000
0!
0%
#603285000000
1!
1%
#603290000000
0!
0%
#603295000000
1!
1%
#603300000000
0!
0%
#603305000000
1!
1%
#603310000000
0!
0%
#603315000000
1!
1%
#603320000000
0!
0%
#603325000000
1!
1%
#603330000000
0!
0%
#603335000000
1!
1%
#603340000000
0!
0%
#603345000000
1!
1%
#603350000000
0!
0%
#603355000000
1!
1%
#603360000000
0!
0%
#603365000000
1!
1%
#603370000000
0!
0%
#603375000000
1!
1%
#603380000000
0!
0%
#603385000000
1!
1%
#603390000000
0!
0%
#603395000000
1!
1%
#603400000000
0!
0%
#603405000000
1!
1%
#603410000000
0!
0%
#603415000000
1!
1%
#603420000000
0!
0%
#603425000000
1!
1%
#603430000000
0!
0%
#603435000000
1!
1%
#603440000000
0!
0%
#603445000000
1!
1%
#603450000000
0!
0%
#603455000000
1!
1%
#603460000000
0!
0%
#603465000000
1!
1%
#603470000000
0!
0%
#603475000000
1!
1%
#603480000000
0!
0%
#603485000000
1!
1%
#603490000000
0!
0%
#603495000000
1!
1%
#603500000000
0!
0%
#603505000000
1!
1%
#603510000000
0!
0%
#603515000000
1!
1%
#603520000000
0!
0%
#603525000000
1!
1%
#603530000000
0!
0%
#603535000000
1!
1%
#603540000000
0!
0%
#603545000000
1!
1%
#603550000000
0!
0%
#603555000000
1!
1%
#603560000000
0!
0%
#603565000000
1!
1%
#603570000000
0!
0%
#603575000000
1!
1%
#603580000000
0!
0%
#603585000000
1!
1%
#603590000000
0!
0%
#603595000000
1!
1%
#603600000000
0!
0%
#603605000000
1!
1%
#603610000000
0!
0%
#603615000000
1!
1%
#603620000000
0!
0%
#603625000000
1!
1%
#603630000000
0!
0%
#603635000000
1!
1%
#603640000000
0!
0%
#603645000000
1!
1%
#603650000000
0!
0%
#603655000000
1!
1%
#603660000000
0!
0%
#603665000000
1!
1%
#603670000000
0!
0%
#603675000000
1!
1%
#603680000000
0!
0%
#603685000000
1!
1%
#603690000000
0!
0%
#603695000000
1!
1%
#603700000000
0!
0%
#603705000000
1!
1%
#603710000000
0!
0%
#603715000000
1!
1%
#603720000000
0!
0%
#603725000000
1!
1%
#603730000000
0!
0%
#603735000000
1!
1%
#603740000000
0!
0%
#603745000000
1!
1%
#603750000000
0!
0%
#603755000000
1!
1%
#603760000000
0!
0%
#603765000000
1!
1%
#603770000000
0!
0%
#603775000000
1!
1%
#603780000000
0!
0%
#603785000000
1!
1%
#603790000000
0!
0%
#603795000000
1!
1%
#603800000000
0!
0%
#603805000000
1!
1%
#603810000000
0!
0%
#603815000000
1!
1%
#603820000000
0!
0%
#603825000000
1!
1%
#603830000000
0!
0%
#603835000000
1!
1%
#603840000000
0!
0%
#603845000000
1!
1%
#603850000000
0!
0%
#603855000000
1!
1%
#603860000000
0!
0%
#603865000000
1!
1%
#603870000000
0!
0%
#603875000000
1!
1%
#603880000000
0!
0%
#603885000000
1!
1%
#603890000000
0!
0%
#603895000000
1!
1%
#603900000000
0!
0%
#603905000000
1!
1%
#603910000000
0!
0%
#603915000000
1!
1%
#603920000000
0!
0%
#603925000000
1!
1%
#603930000000
0!
0%
#603935000000
1!
1%
#603940000000
0!
0%
#603945000000
1!
1%
#603950000000
0!
0%
#603955000000
1!
1%
#603960000000
0!
0%
#603965000000
1!
1%
#603970000000
0!
0%
#603975000000
1!
1%
#603980000000
0!
0%
#603985000000
1!
1%
#603990000000
0!
0%
#603995000000
1!
1%
#604000000000
0!
0%
#604005000000
1!
1%
#604010000000
0!
0%
#604015000000
1!
1%
#604020000000
0!
0%
#604025000000
1!
1%
#604030000000
0!
0%
#604035000000
1!
1%
#604040000000
0!
0%
#604045000000
1!
1%
#604050000000
0!
0%
#604055000000
1!
1%
#604060000000
0!
0%
#604065000000
1!
1%
#604070000000
0!
0%
#604075000000
1!
1%
#604080000000
0!
0%
#604085000000
1!
1%
#604090000000
0!
0%
#604095000000
1!
1%
#604100000000
0!
0%
#604105000000
1!
1%
#604110000000
0!
0%
#604115000000
1!
1%
#604120000000
0!
0%
#604125000000
1!
1%
#604130000000
0!
0%
#604135000000
1!
1%
#604140000000
0!
0%
#604145000000
1!
1%
#604150000000
0!
0%
#604155000000
1!
1%
#604160000000
0!
0%
#604165000000
1!
1%
#604170000000
0!
0%
#604175000000
1!
1%
#604180000000
0!
0%
#604185000000
1!
1%
#604190000000
0!
0%
#604195000000
1!
1%
#604200000000
0!
0%
#604205000000
1!
1%
#604210000000
0!
0%
#604215000000
1!
1%
#604220000000
0!
0%
#604225000000
1!
1%
#604230000000
0!
0%
#604235000000
1!
1%
#604240000000
0!
0%
#604245000000
1!
1%
#604250000000
0!
0%
#604255000000
1!
1%
#604260000000
0!
0%
#604265000000
1!
1%
#604270000000
0!
0%
#604275000000
1!
1%
#604280000000
0!
0%
#604285000000
1!
1%
#604290000000
0!
0%
#604295000000
1!
1%
#604300000000
0!
0%
#604305000000
1!
1%
#604310000000
0!
0%
#604315000000
1!
1%
#604320000000
0!
0%
#604325000000
1!
1%
#604330000000
0!
0%
#604335000000
1!
1%
#604340000000
0!
0%
#604345000000
1!
1%
#604350000000
0!
0%
#604355000000
1!
1%
#604360000000
0!
0%
#604365000000
1!
1%
#604370000000
0!
0%
#604375000000
1!
1%
#604380000000
0!
0%
#604385000000
1!
1%
#604390000000
0!
0%
#604395000000
1!
1%
#604400000000
0!
0%
#604405000000
1!
1%
#604410000000
0!
0%
#604415000000
1!
1%
#604420000000
0!
0%
#604425000000
1!
1%
#604430000000
0!
0%
#604435000000
1!
1%
#604440000000
0!
0%
#604445000000
1!
1%
#604450000000
0!
0%
#604455000000
1!
1%
#604460000000
0!
0%
#604465000000
1!
1%
#604470000000
0!
0%
#604475000000
1!
1%
#604480000000
0!
0%
#604485000000
1!
1%
#604490000000
0!
0%
#604495000000
1!
1%
#604500000000
0!
0%
#604505000000
1!
1%
#604510000000
0!
0%
#604515000000
1!
1%
#604520000000
0!
0%
#604525000000
1!
1%
#604530000000
0!
0%
#604535000000
1!
1%
#604540000000
0!
0%
#604545000000
1!
1%
#604550000000
0!
0%
#604555000000
1!
1%
#604560000000
0!
0%
#604565000000
1!
1%
#604570000000
0!
0%
#604575000000
1!
1%
#604580000000
0!
0%
#604585000000
1!
1%
#604590000000
0!
0%
#604595000000
1!
1%
#604600000000
0!
0%
#604605000000
1!
1%
#604610000000
0!
0%
#604615000000
1!
1%
#604620000000
0!
0%
#604625000000
1!
1%
#604630000000
0!
0%
#604635000000
1!
1%
#604640000000
0!
0%
#604645000000
1!
1%
#604650000000
0!
0%
#604655000000
1!
1%
#604660000000
0!
0%
#604665000000
1!
1%
#604670000000
0!
0%
#604675000000
1!
1%
#604680000000
0!
0%
#604685000000
1!
1%
#604690000000
0!
0%
#604695000000
1!
1%
#604700000000
0!
0%
#604705000000
1!
1%
#604710000000
0!
0%
#604715000000
1!
1%
#604720000000
0!
0%
#604725000000
1!
1%
#604730000000
0!
0%
#604735000000
1!
1%
#604740000000
0!
0%
#604745000000
1!
1%
#604750000000
0!
0%
#604755000000
1!
1%
#604760000000
0!
0%
#604765000000
1!
1%
#604770000000
0!
0%
#604775000000
1!
1%
#604780000000
0!
0%
#604785000000
1!
1%
#604790000000
0!
0%
#604795000000
1!
1%
#604800000000
0!
0%
#604805000000
1!
1%
#604810000000
0!
0%
#604815000000
1!
1%
#604820000000
0!
0%
#604825000000
1!
1%
#604830000000
0!
0%
#604835000000
1!
1%
#604840000000
0!
0%
#604845000000
1!
1%
#604850000000
0!
0%
#604855000000
1!
1%
#604860000000
0!
0%
#604865000000
1!
1%
#604870000000
0!
0%
#604875000000
1!
1%
#604880000000
0!
0%
#604885000000
1!
1%
#604890000000
0!
0%
#604895000000
1!
1%
#604900000000
0!
0%
#604905000000
1!
1%
#604910000000
0!
0%
#604915000000
1!
1%
#604920000000
0!
0%
#604925000000
1!
1%
#604930000000
0!
0%
#604935000000
1!
1%
#604940000000
0!
0%
#604945000000
1!
1%
#604950000000
0!
0%
#604955000000
1!
1%
#604960000000
0!
0%
#604965000000
1!
1%
#604970000000
0!
0%
#604975000000
1!
1%
#604980000000
0!
0%
#604985000000
1!
1%
#604990000000
0!
0%
#604995000000
1!
1%
#605000000000
0!
0%
#605005000000
1!
1%
#605010000000
0!
0%
#605015000000
1!
1%
#605020000000
0!
0%
#605025000000
1!
1%
#605030000000
0!
0%
#605035000000
1!
1%
#605040000000
0!
0%
#605045000000
1!
1%
#605050000000
0!
0%
#605055000000
1!
1%
#605060000000
0!
0%
#605065000000
1!
1%
#605070000000
0!
0%
#605075000000
1!
1%
#605080000000
0!
0%
#605085000000
1!
1%
#605090000000
0!
0%
#605095000000
1!
1%
#605100000000
0!
0%
#605105000000
1!
1%
#605110000000
0!
0%
#605115000000
1!
1%
#605120000000
0!
0%
#605125000000
1!
1%
#605130000000
0!
0%
#605135000000
1!
1%
#605140000000
0!
0%
#605145000000
1!
1%
#605150000000
0!
0%
#605155000000
1!
1%
#605160000000
0!
0%
#605165000000
1!
1%
#605170000000
0!
0%
#605175000000
1!
1%
#605180000000
0!
0%
#605185000000
1!
1%
#605190000000
0!
0%
#605195000000
1!
1%
#605200000000
0!
0%
#605205000000
1!
1%
#605210000000
0!
0%
#605215000000
1!
1%
#605220000000
0!
0%
#605225000000
1!
1%
#605230000000
0!
0%
#605235000000
1!
1%
#605240000000
0!
0%
#605245000000
1!
1%
#605250000000
0!
0%
#605255000000
1!
1%
#605260000000
0!
0%
#605265000000
1!
1%
#605270000000
0!
0%
#605275000000
1!
1%
#605280000000
0!
0%
#605285000000
1!
1%
#605290000000
0!
0%
#605295000000
1!
1%
#605300000000
0!
0%
#605305000000
1!
1%
#605310000000
0!
0%
#605315000000
1!
1%
#605320000000
0!
0%
#605325000000
1!
1%
#605330000000
0!
0%
#605335000000
1!
1%
#605340000000
0!
0%
#605345000000
1!
1%
#605350000000
0!
0%
#605355000000
1!
1%
#605360000000
0!
0%
#605365000000
1!
1%
#605370000000
0!
0%
#605375000000
1!
1%
#605380000000
0!
0%
#605385000000
1!
1%
#605390000000
0!
0%
#605395000000
1!
1%
#605400000000
0!
0%
#605405000000
1!
1%
#605410000000
0!
0%
#605415000000
1!
1%
#605420000000
0!
0%
#605425000000
1!
1%
#605430000000
0!
0%
#605435000000
1!
1%
#605440000000
0!
0%
#605445000000
1!
1%
#605450000000
0!
0%
#605455000000
1!
1%
#605460000000
0!
0%
#605465000000
1!
1%
#605470000000
0!
0%
#605475000000
1!
1%
#605480000000
0!
0%
#605485000000
1!
1%
#605490000000
0!
0%
#605495000000
1!
1%
#605500000000
0!
0%
#605505000000
1!
1%
#605510000000
0!
0%
#605515000000
1!
1%
#605520000000
0!
0%
#605525000000
1!
1%
#605530000000
0!
0%
#605535000000
1!
1%
#605540000000
0!
0%
#605545000000
1!
1%
#605550000000
0!
0%
#605555000000
1!
1%
#605560000000
0!
0%
#605565000000
1!
1%
#605570000000
0!
0%
#605575000000
1!
1%
#605580000000
0!
0%
#605585000000
1!
1%
#605590000000
0!
0%
#605595000000
1!
1%
#605600000000
0!
0%
#605605000000
1!
1%
#605610000000
0!
0%
#605615000000
1!
1%
#605620000000
0!
0%
#605625000000
1!
1%
#605630000000
0!
0%
#605635000000
1!
1%
#605640000000
0!
0%
#605645000000
1!
1%
#605650000000
0!
0%
#605655000000
1!
1%
#605660000000
0!
0%
#605665000000
1!
1%
#605670000000
0!
0%
#605675000000
1!
1%
#605680000000
0!
0%
#605685000000
1!
1%
#605690000000
0!
0%
#605695000000
1!
1%
#605700000000
0!
0%
#605705000000
1!
1%
#605710000000
0!
0%
#605715000000
1!
1%
#605720000000
0!
0%
#605725000000
1!
1%
#605730000000
0!
0%
#605735000000
1!
1%
#605740000000
0!
0%
#605745000000
1!
1%
#605750000000
0!
0%
#605755000000
1!
1%
#605760000000
0!
0%
#605765000000
1!
1%
#605770000000
0!
0%
#605775000000
1!
1%
#605780000000
0!
0%
#605785000000
1!
1%
#605790000000
0!
0%
#605795000000
1!
1%
#605800000000
0!
0%
#605805000000
1!
1%
#605810000000
0!
0%
#605815000000
1!
1%
#605820000000
0!
0%
#605825000000
1!
1%
#605830000000
0!
0%
#605835000000
1!
1%
#605840000000
0!
0%
#605845000000
1!
1%
#605850000000
0!
0%
#605855000000
1!
1%
#605860000000
0!
0%
#605865000000
1!
1%
#605870000000
0!
0%
#605875000000
1!
1%
#605880000000
0!
0%
#605885000000
1!
1%
#605890000000
0!
0%
#605895000000
1!
1%
#605900000000
0!
0%
#605905000000
1!
1%
#605910000000
0!
0%
#605915000000
1!
1%
#605920000000
0!
0%
#605925000000
1!
1%
#605930000000
0!
0%
#605935000000
1!
1%
#605940000000
0!
0%
#605945000000
1!
1%
#605950000000
0!
0%
#605955000000
1!
1%
#605960000000
0!
0%
#605965000000
1!
1%
#605970000000
0!
0%
#605975000000
1!
1%
#605980000000
0!
0%
#605985000000
1!
1%
#605990000000
0!
0%
#605995000000
1!
1%
#606000000000
0!
0%
#606005000000
1!
1%
#606010000000
0!
0%
#606015000000
1!
1%
#606020000000
0!
0%
#606025000000
1!
1%
#606030000000
0!
0%
#606035000000
1!
1%
#606040000000
0!
0%
#606045000000
1!
1%
#606050000000
0!
0%
#606055000000
1!
1%
#606060000000
0!
0%
#606065000000
1!
1%
#606070000000
0!
0%
#606075000000
1!
1%
#606080000000
0!
0%
#606085000000
1!
1%
#606090000000
0!
0%
#606095000000
1!
1%
#606100000000
0!
0%
#606105000000
1!
1%
#606110000000
0!
0%
#606115000000
1!
1%
#606120000000
0!
0%
#606125000000
1!
1%
#606130000000
0!
0%
#606135000000
1!
1%
#606140000000
0!
0%
#606145000000
1!
1%
#606150000000
0!
0%
#606155000000
1!
1%
#606160000000
0!
0%
#606165000000
1!
1%
#606170000000
0!
0%
#606175000000
1!
1%
#606180000000
0!
0%
#606185000000
1!
1%
#606190000000
0!
0%
#606195000000
1!
1%
#606200000000
0!
0%
#606205000000
1!
1%
#606210000000
0!
0%
#606215000000
1!
1%
#606220000000
0!
0%
#606225000000
1!
1%
#606230000000
0!
0%
#606235000000
1!
1%
#606240000000
0!
0%
#606245000000
1!
1%
#606250000000
0!
0%
#606255000000
1!
1%
#606260000000
0!
0%
#606265000000
1!
1%
#606270000000
0!
0%
#606275000000
1!
1%
#606280000000
0!
0%
#606285000000
1!
1%
#606290000000
0!
0%
#606295000000
1!
1%
#606300000000
0!
0%
#606305000000
1!
1%
#606310000000
0!
0%
#606315000000
1!
1%
#606320000000
0!
0%
#606325000000
1!
1%
#606330000000
0!
0%
#606335000000
1!
1%
#606340000000
0!
0%
#606345000000
1!
1%
#606350000000
0!
0%
#606355000000
1!
1%
#606360000000
0!
0%
#606365000000
1!
1%
#606370000000
0!
0%
#606375000000
1!
1%
#606380000000
0!
0%
#606385000000
1!
1%
#606390000000
0!
0%
#606395000000
1!
1%
#606400000000
0!
0%
#606405000000
1!
1%
#606410000000
0!
0%
#606415000000
1!
1%
#606420000000
0!
0%
#606425000000
1!
1%
#606430000000
0!
0%
#606435000000
1!
1%
#606440000000
0!
0%
#606445000000
1!
1%
#606450000000
0!
0%
#606455000000
1!
1%
#606460000000
0!
0%
#606465000000
1!
1%
#606470000000
0!
0%
#606475000000
1!
1%
#606480000000
0!
0%
#606485000000
1!
1%
#606490000000
0!
0%
#606495000000
1!
1%
#606500000000
0!
0%
#606505000000
1!
1%
#606510000000
0!
0%
#606515000000
1!
1%
#606520000000
0!
0%
#606525000000
1!
1%
#606530000000
0!
0%
#606535000000
1!
1%
#606540000000
0!
0%
#606545000000
1!
1%
#606550000000
0!
0%
#606555000000
1!
1%
#606560000000
0!
0%
#606565000000
1!
1%
#606570000000
0!
0%
#606575000000
1!
1%
#606580000000
0!
0%
#606585000000
1!
1%
#606590000000
0!
0%
#606595000000
1!
1%
#606600000000
0!
0%
#606605000000
1!
1%
#606610000000
0!
0%
#606615000000
1!
1%
#606620000000
0!
0%
#606625000000
1!
1%
#606630000000
0!
0%
#606635000000
1!
1%
#606640000000
0!
0%
#606645000000
1!
1%
#606650000000
0!
0%
#606655000000
1!
1%
#606660000000
0!
0%
#606665000000
1!
1%
#606670000000
0!
0%
#606675000000
1!
1%
#606680000000
0!
0%
#606685000000
1!
1%
#606690000000
0!
0%
#606695000000
1!
1%
#606700000000
0!
0%
#606705000000
1!
1%
#606710000000
0!
0%
#606715000000
1!
1%
#606720000000
0!
0%
#606725000000
1!
1%
#606730000000
0!
0%
#606735000000
1!
1%
#606740000000
0!
0%
#606745000000
1!
1%
#606750000000
0!
0%
#606755000000
1!
1%
#606760000000
0!
0%
#606765000000
1!
1%
#606770000000
0!
0%
#606775000000
1!
1%
#606780000000
0!
0%
#606785000000
1!
1%
#606790000000
0!
0%
#606795000000
1!
1%
#606800000000
0!
0%
#606805000000
1!
1%
#606810000000
0!
0%
#606815000000
1!
1%
#606820000000
0!
0%
#606825000000
1!
1%
#606830000000
0!
0%
#606835000000
1!
1%
#606840000000
0!
0%
#606845000000
1!
1%
#606850000000
0!
0%
#606855000000
1!
1%
#606860000000
0!
0%
#606865000000
1!
1%
#606870000000
0!
0%
#606875000000
1!
1%
#606880000000
0!
0%
#606885000000
1!
1%
#606890000000
0!
0%
#606895000000
1!
1%
#606900000000
0!
0%
#606905000000
1!
1%
#606910000000
0!
0%
#606915000000
1!
1%
#606920000000
0!
0%
#606925000000
1!
1%
#606930000000
0!
0%
#606935000000
1!
1%
#606940000000
0!
0%
#606945000000
1!
1%
#606950000000
0!
0%
#606955000000
1!
1%
#606960000000
0!
0%
#606965000000
1!
1%
#606970000000
0!
0%
#606975000000
1!
1%
#606980000000
0!
0%
#606985000000
1!
1%
#606990000000
0!
0%
#606995000000
1!
1%
#607000000000
0!
0%
#607005000000
1!
1%
#607010000000
0!
0%
#607015000000
1!
1%
#607020000000
0!
0%
#607025000000
1!
1%
#607030000000
0!
0%
#607035000000
1!
1%
#607040000000
0!
0%
#607045000000
1!
1%
#607050000000
0!
0%
#607055000000
1!
1%
#607060000000
0!
0%
#607065000000
1!
1%
#607070000000
0!
0%
#607075000000
1!
1%
#607080000000
0!
0%
#607085000000
1!
1%
#607090000000
0!
0%
#607095000000
1!
1%
#607100000000
0!
0%
#607105000000
1!
1%
#607110000000
0!
0%
#607115000000
1!
1%
#607120000000
0!
0%
#607125000000
1!
1%
#607130000000
0!
0%
#607135000000
1!
1%
#607140000000
0!
0%
#607145000000
1!
1%
#607150000000
0!
0%
#607155000000
1!
1%
#607160000000
0!
0%
#607165000000
1!
1%
#607170000000
0!
0%
#607175000000
1!
1%
#607180000000
0!
0%
#607185000000
1!
1%
#607190000000
0!
0%
#607195000000
1!
1%
#607200000000
0!
0%
#607205000000
1!
1%
#607210000000
0!
0%
#607215000000
1!
1%
#607220000000
0!
0%
#607225000000
1!
1%
#607230000000
0!
0%
#607235000000
1!
1%
#607240000000
0!
0%
#607245000000
1!
1%
#607250000000
0!
0%
#607255000000
1!
1%
#607260000000
0!
0%
#607265000000
1!
1%
#607270000000
0!
0%
#607275000000
1!
1%
#607280000000
0!
0%
#607285000000
1!
1%
#607290000000
0!
0%
#607295000000
1!
1%
#607300000000
0!
0%
#607305000000
1!
1%
#607310000000
0!
0%
#607315000000
1!
1%
#607320000000
0!
0%
#607325000000
1!
1%
#607330000000
0!
0%
#607335000000
1!
1%
#607340000000
0!
0%
#607345000000
1!
1%
#607350000000
0!
0%
#607355000000
1!
1%
#607360000000
0!
0%
#607365000000
1!
1%
#607370000000
0!
0%
#607375000000
1!
1%
#607380000000
0!
0%
#607385000000
1!
1%
#607390000000
0!
0%
#607395000000
1!
1%
#607400000000
0!
0%
#607405000000
1!
1%
#607410000000
0!
0%
#607415000000
1!
1%
#607420000000
0!
0%
#607425000000
1!
1%
#607430000000
0!
0%
#607435000000
1!
1%
#607440000000
0!
0%
#607445000000
1!
1%
#607450000000
0!
0%
#607455000000
1!
1%
#607460000000
0!
0%
#607465000000
1!
1%
#607470000000
0!
0%
#607475000000
1!
1%
#607480000000
0!
0%
#607485000000
1!
1%
#607490000000
0!
0%
#607495000000
1!
1%
#607500000000
0!
0%
#607505000000
1!
1%
#607510000000
0!
0%
#607515000000
1!
1%
#607520000000
0!
0%
#607525000000
1!
1%
#607530000000
0!
0%
#607535000000
1!
1%
#607540000000
0!
0%
#607545000000
1!
1%
#607550000000
0!
0%
#607555000000
1!
1%
#607560000000
0!
0%
#607565000000
1!
1%
#607570000000
0!
0%
#607575000000
1!
1%
#607580000000
0!
0%
#607585000000
1!
1%
#607590000000
0!
0%
#607595000000
1!
1%
#607600000000
0!
0%
#607605000000
1!
1%
#607610000000
0!
0%
#607615000000
1!
1%
#607620000000
0!
0%
#607625000000
1!
1%
#607630000000
0!
0%
#607635000000
1!
1%
#607640000000
0!
0%
#607645000000
1!
1%
#607650000000
0!
0%
#607655000000
1!
1%
#607660000000
0!
0%
#607665000000
1!
1%
#607670000000
0!
0%
#607675000000
1!
1%
#607680000000
0!
0%
#607685000000
1!
1%
#607690000000
0!
0%
#607695000000
1!
1%
#607700000000
0!
0%
#607705000000
1!
1%
#607710000000
0!
0%
#607715000000
1!
1%
#607720000000
0!
0%
#607725000000
1!
1%
#607730000000
0!
0%
#607735000000
1!
1%
#607740000000
0!
0%
#607745000000
1!
1%
#607750000000
0!
0%
#607755000000
1!
1%
#607760000000
0!
0%
#607765000000
1!
1%
#607770000000
0!
0%
#607775000000
1!
1%
#607780000000
0!
0%
#607785000000
1!
1%
#607790000000
0!
0%
#607795000000
1!
1%
#607800000000
0!
0%
#607805000000
1!
1%
#607810000000
0!
0%
#607815000000
1!
1%
#607820000000
0!
0%
#607825000000
1!
1%
#607830000000
0!
0%
#607835000000
1!
1%
#607840000000
0!
0%
#607845000000
1!
1%
#607850000000
0!
0%
#607855000000
1!
1%
#607860000000
0!
0%
#607865000000
1!
1%
#607870000000
0!
0%
#607875000000
1!
1%
#607880000000
0!
0%
#607885000000
1!
1%
#607890000000
0!
0%
#607895000000
1!
1%
#607900000000
0!
0%
#607905000000
1!
1%
#607910000000
0!
0%
#607915000000
1!
1%
#607920000000
0!
0%
#607925000000
1!
1%
#607930000000
0!
0%
#607935000000
1!
1%
#607940000000
0!
0%
#607945000000
1!
1%
#607950000000
0!
0%
#607955000000
1!
1%
#607960000000
0!
0%
#607965000000
1!
1%
#607970000000
0!
0%
#607975000000
1!
1%
#607980000000
0!
0%
#607985000000
1!
1%
#607990000000
0!
0%
#607995000000
1!
1%
#608000000000
0!
0%
#608005000000
1!
1%
#608010000000
0!
0%
#608015000000
1!
1%
#608020000000
0!
0%
#608025000000
1!
1%
#608030000000
0!
0%
#608035000000
1!
1%
#608040000000
0!
0%
#608045000000
1!
1%
#608050000000
0!
0%
#608055000000
1!
1%
#608060000000
0!
0%
#608065000000
1!
1%
#608070000000
0!
0%
#608075000000
1!
1%
#608080000000
0!
0%
#608085000000
1!
1%
#608090000000
0!
0%
#608095000000
1!
1%
#608100000000
0!
0%
#608105000000
1!
1%
#608110000000
0!
0%
#608115000000
1!
1%
#608120000000
0!
0%
#608125000000
1!
1%
#608130000000
0!
0%
#608135000000
1!
1%
#608140000000
0!
0%
#608145000000
1!
1%
#608150000000
0!
0%
#608155000000
1!
1%
#608160000000
0!
0%
#608165000000
1!
1%
#608170000000
0!
0%
#608175000000
1!
1%
#608180000000
0!
0%
#608185000000
1!
1%
#608190000000
0!
0%
#608195000000
1!
1%
#608200000000
0!
0%
#608205000000
1!
1%
#608210000000
0!
0%
#608215000000
1!
1%
#608220000000
0!
0%
#608225000000
1!
1%
#608230000000
0!
0%
#608235000000
1!
1%
#608240000000
0!
0%
#608245000000
1!
1%
#608250000000
0!
0%
#608255000000
1!
1%
#608260000000
0!
0%
#608265000000
1!
1%
#608270000000
0!
0%
#608275000000
1!
1%
#608280000000
0!
0%
#608285000000
1!
1%
#608290000000
0!
0%
#608295000000
1!
1%
#608300000000
0!
0%
#608305000000
1!
1%
#608310000000
0!
0%
#608315000000
1!
1%
#608320000000
0!
0%
#608325000000
1!
1%
#608330000000
0!
0%
#608335000000
1!
1%
#608340000000
0!
0%
#608345000000
1!
1%
#608350000000
0!
0%
#608355000000
1!
1%
#608360000000
0!
0%
#608365000000
1!
1%
#608370000000
0!
0%
#608375000000
1!
1%
#608380000000
0!
0%
#608385000000
1!
1%
#608390000000
0!
0%
#608395000000
1!
1%
#608400000000
0!
0%
#608405000000
1!
1%
#608410000000
0!
0%
#608415000000
1!
1%
#608420000000
0!
0%
#608425000000
1!
1%
#608430000000
0!
0%
#608435000000
1!
1%
#608440000000
0!
0%
#608445000000
1!
1%
#608450000000
0!
0%
#608455000000
1!
1%
#608460000000
0!
0%
#608465000000
1!
1%
#608470000000
0!
0%
#608475000000
1!
1%
#608480000000
0!
0%
#608485000000
1!
1%
#608490000000
0!
0%
#608495000000
1!
1%
#608500000000
0!
0%
#608505000000
1!
1%
#608510000000
0!
0%
#608515000000
1!
1%
#608520000000
0!
0%
#608525000000
1!
1%
#608530000000
0!
0%
#608535000000
1!
1%
#608540000000
0!
0%
#608545000000
1!
1%
#608550000000
0!
0%
#608555000000
1!
1%
#608560000000
0!
0%
#608565000000
1!
1%
#608570000000
0!
0%
#608575000000
1!
1%
#608580000000
0!
0%
#608585000000
1!
1%
#608590000000
0!
0%
#608595000000
1!
1%
#608600000000
0!
0%
#608605000000
1!
1%
#608610000000
0!
0%
#608615000000
1!
1%
#608620000000
0!
0%
#608625000000
1!
1%
#608630000000
0!
0%
#608635000000
1!
1%
#608640000000
0!
0%
#608645000000
1!
1%
#608650000000
0!
0%
#608655000000
1!
1%
#608660000000
0!
0%
#608665000000
1!
1%
#608670000000
0!
0%
#608675000000
1!
1%
#608680000000
0!
0%
#608685000000
1!
1%
#608690000000
0!
0%
#608695000000
1!
1%
#608700000000
0!
0%
#608705000000
1!
1%
#608710000000
0!
0%
#608715000000
1!
1%
#608720000000
0!
0%
#608725000000
1!
1%
#608730000000
0!
0%
#608735000000
1!
1%
#608740000000
0!
0%
#608745000000
1!
1%
#608750000000
0!
0%
#608755000000
1!
1%
#608760000000
0!
0%
#608765000000
1!
1%
#608770000000
0!
0%
#608775000000
1!
1%
#608780000000
0!
0%
#608785000000
1!
1%
#608790000000
0!
0%
#608795000000
1!
1%
#608800000000
0!
0%
#608805000000
1!
1%
#608810000000
0!
0%
#608815000000
1!
1%
#608820000000
0!
0%
#608825000000
1!
1%
#608830000000
0!
0%
#608835000000
1!
1%
#608840000000
0!
0%
#608845000000
1!
1%
#608850000000
0!
0%
#608855000000
1!
1%
#608860000000
0!
0%
#608865000000
1!
1%
#608870000000
0!
0%
#608875000000
1!
1%
#608880000000
0!
0%
#608885000000
1!
1%
#608890000000
0!
0%
#608895000000
1!
1%
#608900000000
0!
0%
#608905000000
1!
1%
#608910000000
0!
0%
#608915000000
1!
1%
#608920000000
0!
0%
#608925000000
1!
1%
#608930000000
0!
0%
#608935000000
1!
1%
#608940000000
0!
0%
#608945000000
1!
1%
#608950000000
0!
0%
#608955000000
1!
1%
#608960000000
0!
0%
#608965000000
1!
1%
#608970000000
0!
0%
#608975000000
1!
1%
#608980000000
0!
0%
#608985000000
1!
1%
#608990000000
0!
0%
#608995000000
1!
1%
#609000000000
0!
0%
#609005000000
1!
1%
#609010000000
0!
0%
#609015000000
1!
1%
#609020000000
0!
0%
#609025000000
1!
1%
#609030000000
0!
0%
#609035000000
1!
1%
#609040000000
0!
0%
#609045000000
1!
1%
#609050000000
0!
0%
#609055000000
1!
1%
#609060000000
0!
0%
#609065000000
1!
1%
#609070000000
0!
0%
#609075000000
1!
1%
#609080000000
0!
0%
#609085000000
1!
1%
#609090000000
0!
0%
#609095000000
1!
1%
#609100000000
0!
0%
#609105000000
1!
1%
#609110000000
0!
0%
#609115000000
1!
1%
#609120000000
0!
0%
#609125000000
1!
1%
#609130000000
0!
0%
#609135000000
1!
1%
#609140000000
0!
0%
#609145000000
1!
1%
#609150000000
0!
0%
#609155000000
1!
1%
#609160000000
0!
0%
#609165000000
1!
1%
#609170000000
0!
0%
#609175000000
1!
1%
#609180000000
0!
0%
#609185000000
1!
1%
#609190000000
0!
0%
#609195000000
1!
1%
#609200000000
0!
0%
#609205000000
1!
1%
#609210000000
0!
0%
#609215000000
1!
1%
#609220000000
0!
0%
#609225000000
1!
1%
#609230000000
0!
0%
#609235000000
1!
1%
#609240000000
0!
0%
#609245000000
1!
1%
#609250000000
0!
0%
#609255000000
1!
1%
#609260000000
0!
0%
#609265000000
1!
1%
#609270000000
0!
0%
#609275000000
1!
1%
#609280000000
0!
0%
#609285000000
1!
1%
#609290000000
0!
0%
#609295000000
1!
1%
#609300000000
0!
0%
#609305000000
1!
1%
#609310000000
0!
0%
#609315000000
1!
1%
#609320000000
0!
0%
#609325000000
1!
1%
#609330000000
0!
0%
#609335000000
1!
1%
#609340000000
0!
0%
#609345000000
1!
1%
#609350000000
0!
0%
#609355000000
1!
1%
#609360000000
0!
0%
#609365000000
1!
1%
#609370000000
0!
0%
#609375000000
1!
1%
#609380000000
0!
0%
#609385000000
1!
1%
#609390000000
0!
0%
#609395000000
1!
1%
#609400000000
0!
0%
#609405000000
1!
1%
#609410000000
0!
0%
#609415000000
1!
1%
#609420000000
0!
0%
#609425000000
1!
1%
#609430000000
0!
0%
#609435000000
1!
1%
#609440000000
0!
0%
#609445000000
1!
1%
#609450000000
0!
0%
#609455000000
1!
1%
#609460000000
0!
0%
#609465000000
1!
1%
#609470000000
0!
0%
#609475000000
1!
1%
#609480000000
0!
0%
#609485000000
1!
1%
#609490000000
0!
0%
#609495000000
1!
1%
#609500000000
0!
0%
#609505000000
1!
1%
#609510000000
0!
0%
#609515000000
1!
1%
#609520000000
0!
0%
#609525000000
1!
1%
#609530000000
0!
0%
#609535000000
1!
1%
#609540000000
0!
0%
#609545000000
1!
1%
#609550000000
0!
0%
#609555000000
1!
1%
#609560000000
0!
0%
#609565000000
1!
1%
#609570000000
0!
0%
#609575000000
1!
1%
#609580000000
0!
0%
#609585000000
1!
1%
#609590000000
0!
0%
#609595000000
1!
1%
#609600000000
0!
0%
#609605000000
1!
1%
#609610000000
0!
0%
#609615000000
1!
1%
#609620000000
0!
0%
#609625000000
1!
1%
#609630000000
0!
0%
#609635000000
1!
1%
#609640000000
0!
0%
#609645000000
1!
1%
#609650000000
0!
0%
#609655000000
1!
1%
#609660000000
0!
0%
#609665000000
1!
1%
#609670000000
0!
0%
#609675000000
1!
1%
#609680000000
0!
0%
#609685000000
1!
1%
#609690000000
0!
0%
#609695000000
1!
1%
#609700000000
0!
0%
#609705000000
1!
1%
#609710000000
0!
0%
#609715000000
1!
1%
#609720000000
0!
0%
#609725000000
1!
1%
#609730000000
0!
0%
#609735000000
1!
1%
#609740000000
0!
0%
#609745000000
1!
1%
#609750000000
0!
0%
#609755000000
1!
1%
#609760000000
0!
0%
#609765000000
1!
1%
#609770000000
0!
0%
#609775000000
1!
1%
#609780000000
0!
0%
#609785000000
1!
1%
#609790000000
0!
0%
#609795000000
1!
1%
#609800000000
0!
0%
#609805000000
1!
1%
#609810000000
0!
0%
#609815000000
1!
1%
#609820000000
0!
0%
#609825000000
1!
1%
#609830000000
0!
0%
#609835000000
1!
1%
#609840000000
0!
0%
#609845000000
1!
1%
#609850000000
0!
0%
#609855000000
1!
1%
#609860000000
0!
0%
#609865000000
1!
1%
#609870000000
0!
0%
#609875000000
1!
1%
#609880000000
0!
0%
#609885000000
1!
1%
#609890000000
0!
0%
#609895000000
1!
1%
#609900000000
0!
0%
#609905000000
1!
1%
#609910000000
0!
0%
#609915000000
1!
1%
#609920000000
0!
0%
#609925000000
1!
1%
#609930000000
0!
0%
#609935000000
1!
1%
#609940000000
0!
0%
#609945000000
1!
1%
#609950000000
0!
0%
#609955000000
1!
1%
#609960000000
0!
0%
#609965000000
1!
1%
#609970000000
0!
0%
#609975000000
1!
1%
#609980000000
0!
0%
#609985000000
1!
1%
#609990000000
0!
0%
#609995000000
1!
1%
#610000000000
0!
0%
#610005000000
1!
1%
#610010000000
0!
0%
#610015000000
1!
1%
#610020000000
0!
0%
#610025000000
1!
1%
#610030000000
0!
0%
#610035000000
1!
1%
#610040000000
0!
0%
#610045000000
1!
1%
#610050000000
0!
0%
#610055000000
1!
1%
#610060000000
0!
0%
#610065000000
1!
1%
#610070000000
0!
0%
#610075000000
1!
1%
#610080000000
0!
0%
#610085000000
1!
1%
#610090000000
0!
0%
#610095000000
1!
1%
#610100000000
0!
0%
#610105000000
1!
1%
#610110000000
0!
0%
#610115000000
1!
1%
#610120000000
0!
0%
#610125000000
1!
1%
#610130000000
0!
0%
#610135000000
1!
1%
#610140000000
0!
0%
#610145000000
1!
1%
#610150000000
0!
0%
#610155000000
1!
1%
#610160000000
0!
0%
#610165000000
1!
1%
#610170000000
0!
0%
#610175000000
1!
1%
#610180000000
0!
0%
#610185000000
1!
1%
#610190000000
0!
0%
#610195000000
1!
1%
#610200000000
0!
0%
#610205000000
1!
1%
#610210000000
0!
0%
#610215000000
1!
1%
#610220000000
0!
0%
#610225000000
1!
1%
#610230000000
0!
0%
#610235000000
1!
1%
#610240000000
0!
0%
#610245000000
1!
1%
#610250000000
0!
0%
#610255000000
1!
1%
#610260000000
0!
0%
#610265000000
1!
1%
#610270000000
0!
0%
#610275000000
1!
1%
#610280000000
0!
0%
#610285000000
1!
1%
#610290000000
0!
0%
#610295000000
1!
1%
#610300000000
0!
0%
#610305000000
1!
1%
#610310000000
0!
0%
#610315000000
1!
1%
#610320000000
0!
0%
#610325000000
1!
1%
#610330000000
0!
0%
#610335000000
1!
1%
#610340000000
0!
0%
#610345000000
1!
1%
#610350000000
0!
0%
#610355000000
1!
1%
#610360000000
0!
0%
#610365000000
1!
1%
#610370000000
0!
0%
#610375000000
1!
1%
#610380000000
0!
0%
#610385000000
1!
1%
#610390000000
0!
0%
#610395000000
1!
1%
#610400000000
0!
0%
#610405000000
1!
1%
#610410000000
0!
0%
#610415000000
1!
1%
#610420000000
0!
0%
#610425000000
1!
1%
#610430000000
0!
0%
#610435000000
1!
1%
#610440000000
0!
0%
#610445000000
1!
1%
#610450000000
0!
0%
#610455000000
1!
1%
#610460000000
0!
0%
#610465000000
1!
1%
#610470000000
0!
0%
#610475000000
1!
1%
#610480000000
0!
0%
#610485000000
1!
1%
#610490000000
0!
0%
#610495000000
1!
1%
#610500000000
0!
0%
#610505000000
1!
1%
#610510000000
0!
0%
#610515000000
1!
1%
#610520000000
0!
0%
#610525000000
1!
1%
#610530000000
0!
0%
#610535000000
1!
1%
#610540000000
0!
0%
#610545000000
1!
1%
#610550000000
0!
0%
#610555000000
1!
1%
#610560000000
0!
0%
#610565000000
1!
1%
#610570000000
0!
0%
#610575000000
1!
1%
#610580000000
0!
0%
#610585000000
1!
1%
#610590000000
0!
0%
#610595000000
1!
1%
#610600000000
0!
0%
#610605000000
1!
1%
#610610000000
0!
0%
#610615000000
1!
1%
#610620000000
0!
0%
#610625000000
1!
1%
#610630000000
0!
0%
#610635000000
1!
1%
#610640000000
0!
0%
#610645000000
1!
1%
#610650000000
0!
0%
#610655000000
1!
1%
#610660000000
0!
0%
#610665000000
1!
1%
#610670000000
0!
0%
#610675000000
1!
1%
#610680000000
0!
0%
#610685000000
1!
1%
#610690000000
0!
0%
#610695000000
1!
1%
#610700000000
0!
0%
#610705000000
1!
1%
#610710000000
0!
0%
#610715000000
1!
1%
#610720000000
0!
0%
#610725000000
1!
1%
#610730000000
0!
0%
#610735000000
1!
1%
#610740000000
0!
0%
#610745000000
1!
1%
#610750000000
0!
0%
#610755000000
1!
1%
#610760000000
0!
0%
#610765000000
1!
1%
#610770000000
0!
0%
#610775000000
1!
1%
#610780000000
0!
0%
#610785000000
1!
1%
#610790000000
0!
0%
#610795000000
1!
1%
#610800000000
0!
0%
#610805000000
1!
1%
#610810000000
0!
0%
#610815000000
1!
1%
#610820000000
0!
0%
#610825000000
1!
1%
#610830000000
0!
0%
#610835000000
1!
1%
#610840000000
0!
0%
#610845000000
1!
1%
#610850000000
0!
0%
#610855000000
1!
1%
#610860000000
0!
0%
#610865000000
1!
1%
#610870000000
0!
0%
#610875000000
1!
1%
#610880000000
0!
0%
#610885000000
1!
1%
#610890000000
0!
0%
#610895000000
1!
1%
#610900000000
0!
0%
#610905000000
1!
1%
#610910000000
0!
0%
#610915000000
1!
1%
#610920000000
0!
0%
#610925000000
1!
1%
#610930000000
0!
0%
#610935000000
1!
1%
#610940000000
0!
0%
#610945000000
1!
1%
#610950000000
0!
0%
#610955000000
1!
1%
#610960000000
0!
0%
#610965000000
1!
1%
#610970000000
0!
0%
#610975000000
1!
1%
#610980000000
0!
0%
#610985000000
1!
1%
#610990000000
0!
0%
#610995000000
1!
1%
#611000000000
0!
0%
#611005000000
1!
1%
#611010000000
0!
0%
#611015000000
1!
1%
#611020000000
0!
0%
#611025000000
1!
1%
#611030000000
0!
0%
#611035000000
1!
1%
#611040000000
0!
0%
#611045000000
1!
1%
#611050000000
0!
0%
#611055000000
1!
1%
#611060000000
0!
0%
#611065000000
1!
1%
#611070000000
0!
0%
#611075000000
1!
1%
#611080000000
0!
0%
#611085000000
1!
1%
#611090000000
0!
0%
#611095000000
1!
1%
#611100000000
0!
0%
#611105000000
1!
1%
#611110000000
0!
0%
#611115000000
1!
1%
#611120000000
0!
0%
#611125000000
1!
1%
#611130000000
0!
0%
#611135000000
1!
1%
#611140000000
0!
0%
#611145000000
1!
1%
#611150000000
0!
0%
#611155000000
1!
1%
#611160000000
0!
0%
#611165000000
1!
1%
#611170000000
0!
0%
#611175000000
1!
1%
#611180000000
0!
0%
#611185000000
1!
1%
#611190000000
0!
0%
#611195000000
1!
1%
#611200000000
0!
0%
#611205000000
1!
1%
#611210000000
0!
0%
#611215000000
1!
1%
#611220000000
0!
0%
#611225000000
1!
1%
#611230000000
0!
0%
#611235000000
1!
1%
#611240000000
0!
0%
#611245000000
1!
1%
#611250000000
0!
0%
#611255000000
1!
1%
#611260000000
0!
0%
#611265000000
1!
1%
#611270000000
0!
0%
#611275000000
1!
1%
#611280000000
0!
0%
#611285000000
1!
1%
#611290000000
0!
0%
#611295000000
1!
1%
#611300000000
0!
0%
#611305000000
1!
1%
#611310000000
0!
0%
#611315000000
1!
1%
#611320000000
0!
0%
#611325000000
1!
1%
#611330000000
0!
0%
#611335000000
1!
1%
#611340000000
0!
0%
#611345000000
1!
1%
#611350000000
0!
0%
#611355000000
1!
1%
#611360000000
0!
0%
#611365000000
1!
1%
#611370000000
0!
0%
#611375000000
1!
1%
#611380000000
0!
0%
#611385000000
1!
1%
#611390000000
0!
0%
#611395000000
1!
1%
#611400000000
0!
0%
#611405000000
1!
1%
#611410000000
0!
0%
#611415000000
1!
1%
#611420000000
0!
0%
#611425000000
1!
1%
#611430000000
0!
0%
#611435000000
1!
1%
#611440000000
0!
0%
#611445000000
1!
1%
#611450000000
0!
0%
#611455000000
1!
1%
#611460000000
0!
0%
#611465000000
1!
1%
#611470000000
0!
0%
#611475000000
1!
1%
#611480000000
0!
0%
#611485000000
1!
1%
#611490000000
0!
0%
#611495000000
1!
1%
#611500000000
0!
0%
#611505000000
1!
1%
#611510000000
0!
0%
#611515000000
1!
1%
#611520000000
0!
0%
#611525000000
1!
1%
#611530000000
0!
0%
#611535000000
1!
1%
#611540000000
0!
0%
#611545000000
1!
1%
#611550000000
0!
0%
#611555000000
1!
1%
#611560000000
0!
0%
#611565000000
1!
1%
#611570000000
0!
0%
#611575000000
1!
1%
#611580000000
0!
0%
#611585000000
1!
1%
#611590000000
0!
0%
#611595000000
1!
1%
#611600000000
0!
0%
#611605000000
1!
1%
#611610000000
0!
0%
#611615000000
1!
1%
#611620000000
0!
0%
#611625000000
1!
1%
#611630000000
0!
0%
#611635000000
1!
1%
#611640000000
0!
0%
#611645000000
1!
1%
#611650000000
0!
0%
#611655000000
1!
1%
#611660000000
0!
0%
#611665000000
1!
1%
#611670000000
0!
0%
#611675000000
1!
1%
#611680000000
0!
0%
#611685000000
1!
1%
#611690000000
0!
0%
#611695000000
1!
1%
#611700000000
0!
0%
#611705000000
1!
1%
#611710000000
0!
0%
#611715000000
1!
1%
#611720000000
0!
0%
#611725000000
1!
1%
#611730000000
0!
0%
#611735000000
1!
1%
#611740000000
0!
0%
#611745000000
1!
1%
#611750000000
0!
0%
#611755000000
1!
1%
#611760000000
0!
0%
#611765000000
1!
1%
#611770000000
0!
0%
#611775000000
1!
1%
#611780000000
0!
0%
#611785000000
1!
1%
#611790000000
0!
0%
#611795000000
1!
1%
#611800000000
0!
0%
#611805000000
1!
1%
#611810000000
0!
0%
#611815000000
1!
1%
#611820000000
0!
0%
#611825000000
1!
1%
#611830000000
0!
0%
#611835000000
1!
1%
#611840000000
0!
0%
#611845000000
1!
1%
#611850000000
0!
0%
#611855000000
1!
1%
#611860000000
0!
0%
#611865000000
1!
1%
#611870000000
0!
0%
#611875000000
1!
1%
#611880000000
0!
0%
#611885000000
1!
1%
#611890000000
0!
0%
#611895000000
1!
1%
#611900000000
0!
0%
#611905000000
1!
1%
#611910000000
0!
0%
#611915000000
1!
1%
#611920000000
0!
0%
#611925000000
1!
1%
#611930000000
0!
0%
#611935000000
1!
1%
#611940000000
0!
0%
#611945000000
1!
1%
#611950000000
0!
0%
#611955000000
1!
1%
#611960000000
0!
0%
#611965000000
1!
1%
#611970000000
0!
0%
#611975000000
1!
1%
#611980000000
0!
0%
#611985000000
1!
1%
#611990000000
0!
0%
#611995000000
1!
1%
#612000000000
0!
0%
#612005000000
1!
1%
#612010000000
0!
0%
#612015000000
1!
1%
#612020000000
0!
0%
#612025000000
1!
1%
#612030000000
0!
0%
#612035000000
1!
1%
#612040000000
0!
0%
#612045000000
1!
1%
#612050000000
0!
0%
#612055000000
1!
1%
#612060000000
0!
0%
#612065000000
1!
1%
#612070000000
0!
0%
#612075000000
1!
1%
#612080000000
0!
0%
#612085000000
1!
1%
#612090000000
0!
0%
#612095000000
1!
1%
#612100000000
0!
0%
#612105000000
1!
1%
#612110000000
0!
0%
#612115000000
1!
1%
#612120000000
0!
0%
#612125000000
1!
1%
#612130000000
0!
0%
#612135000000
1!
1%
#612140000000
0!
0%
#612145000000
1!
1%
#612150000000
0!
0%
#612155000000
1!
1%
#612160000000
0!
0%
#612165000000
1!
1%
#612170000000
0!
0%
#612175000000
1!
1%
#612180000000
0!
0%
#612185000000
1!
1%
#612190000000
0!
0%
#612195000000
1!
1%
#612200000000
0!
0%
#612205000000
1!
1%
#612210000000
0!
0%
#612215000000
1!
1%
#612220000000
0!
0%
#612225000000
1!
1%
#612230000000
0!
0%
#612235000000
1!
1%
#612240000000
0!
0%
#612245000000
1!
1%
#612250000000
0!
0%
#612255000000
1!
1%
#612260000000
0!
0%
#612265000000
1!
1%
#612270000000
0!
0%
#612275000000
1!
1%
#612280000000
0!
0%
#612285000000
1!
1%
#612290000000
0!
0%
#612295000000
1!
1%
#612300000000
0!
0%
#612305000000
1!
1%
#612310000000
0!
0%
#612315000000
1!
1%
#612320000000
0!
0%
#612325000000
1!
1%
#612330000000
0!
0%
#612335000000
1!
1%
#612340000000
0!
0%
#612345000000
1!
1%
#612350000000
0!
0%
#612355000000
1!
1%
#612360000000
0!
0%
#612365000000
1!
1%
#612370000000
0!
0%
#612375000000
1!
1%
#612380000000
0!
0%
#612385000000
1!
1%
#612390000000
0!
0%
#612395000000
1!
1%
#612400000000
0!
0%
#612405000000
1!
1%
#612410000000
0!
0%
#612415000000
1!
1%
#612420000000
0!
0%
#612425000000
1!
1%
#612430000000
0!
0%
#612435000000
1!
1%
#612440000000
0!
0%
#612445000000
1!
1%
#612450000000
0!
0%
#612455000000
1!
1%
#612460000000
0!
0%
#612465000000
1!
1%
#612470000000
0!
0%
#612475000000
1!
1%
#612480000000
0!
0%
#612485000000
1!
1%
#612490000000
0!
0%
#612495000000
1!
1%
#612500000000
0!
0%
#612505000000
1!
1%
#612510000000
0!
0%
#612515000000
1!
1%
#612520000000
0!
0%
#612525000000
1!
1%
#612530000000
0!
0%
#612535000000
1!
1%
#612540000000
0!
0%
#612545000000
1!
1%
#612550000000
0!
0%
#612555000000
1!
1%
#612560000000
0!
0%
#612565000000
1!
1%
#612570000000
0!
0%
#612575000000
1!
1%
#612580000000
0!
0%
#612585000000
1!
1%
#612590000000
0!
0%
#612595000000
1!
1%
#612600000000
0!
0%
#612605000000
1!
1%
#612610000000
0!
0%
#612615000000
1!
1%
#612620000000
0!
0%
#612625000000
1!
1%
#612630000000
0!
0%
#612635000000
1!
1%
#612640000000
0!
0%
#612645000000
1!
1%
#612650000000
0!
0%
#612655000000
1!
1%
#612660000000
0!
0%
#612665000000
1!
1%
#612670000000
0!
0%
#612675000000
1!
1%
#612680000000
0!
0%
#612685000000
1!
1%
#612690000000
0!
0%
#612695000000
1!
1%
#612700000000
0!
0%
#612705000000
1!
1%
#612710000000
0!
0%
#612715000000
1!
1%
#612720000000
0!
0%
#612725000000
1!
1%
#612730000000
0!
0%
#612735000000
1!
1%
#612740000000
0!
0%
#612745000000
1!
1%
#612750000000
0!
0%
#612755000000
1!
1%
#612760000000
0!
0%
#612765000000
1!
1%
#612770000000
0!
0%
#612775000000
1!
1%
#612780000000
0!
0%
#612785000000
1!
1%
#612790000000
0!
0%
#612795000000
1!
1%
#612800000000
0!
0%
#612805000000
1!
1%
#612810000000
0!
0%
#612815000000
1!
1%
#612820000000
0!
0%
#612825000000
1!
1%
#612830000000
0!
0%
#612835000000
1!
1%
#612840000000
0!
0%
#612845000000
1!
1%
#612850000000
0!
0%
#612855000000
1!
1%
#612860000000
0!
0%
#612865000000
1!
1%
#612870000000
0!
0%
#612875000000
1!
1%
#612880000000
0!
0%
#612885000000
1!
1%
#612890000000
0!
0%
#612895000000
1!
1%
#612900000000
0!
0%
#612905000000
1!
1%
#612910000000
0!
0%
#612915000000
1!
1%
#612920000000
0!
0%
#612925000000
1!
1%
#612930000000
0!
0%
#612935000000
1!
1%
#612940000000
0!
0%
#612945000000
1!
1%
#612950000000
0!
0%
#612955000000
1!
1%
#612960000000
0!
0%
#612965000000
1!
1%
#612970000000
0!
0%
#612975000000
1!
1%
#612980000000
0!
0%
#612985000000
1!
1%
#612990000000
0!
0%
#612995000000
1!
1%
#613000000000
0!
0%
#613005000000
1!
1%
#613010000000
0!
0%
#613015000000
1!
1%
#613020000000
0!
0%
#613025000000
1!
1%
#613030000000
0!
0%
#613035000000
1!
1%
#613040000000
0!
0%
#613045000000
1!
1%
#613050000000
0!
0%
#613055000000
1!
1%
#613060000000
0!
0%
#613065000000
1!
1%
#613070000000
0!
0%
#613075000000
1!
1%
#613080000000
0!
0%
#613085000000
1!
1%
#613090000000
0!
0%
#613095000000
1!
1%
#613100000000
0!
0%
#613105000000
1!
1%
#613110000000
0!
0%
#613115000000
1!
1%
#613120000000
0!
0%
#613125000000
1!
1%
#613130000000
0!
0%
#613135000000
1!
1%
#613140000000
0!
0%
#613145000000
1!
1%
#613150000000
0!
0%
#613155000000
1!
1%
#613160000000
0!
0%
#613165000000
1!
1%
#613170000000
0!
0%
#613175000000
1!
1%
#613180000000
0!
0%
#613185000000
1!
1%
#613190000000
0!
0%
#613195000000
1!
1%
#613200000000
0!
0%
#613205000000
1!
1%
#613210000000
0!
0%
#613215000000
1!
1%
#613220000000
0!
0%
#613225000000
1!
1%
#613230000000
0!
0%
#613235000000
1!
1%
#613240000000
0!
0%
#613245000000
1!
1%
#613250000000
0!
0%
#613255000000
1!
1%
#613260000000
0!
0%
#613265000000
1!
1%
#613270000000
0!
0%
#613275000000
1!
1%
#613280000000
0!
0%
#613285000000
1!
1%
#613290000000
0!
0%
#613295000000
1!
1%
#613300000000
0!
0%
#613305000000
1!
1%
#613310000000
0!
0%
#613315000000
1!
1%
#613320000000
0!
0%
#613325000000
1!
1%
#613330000000
0!
0%
#613335000000
1!
1%
#613340000000
0!
0%
#613345000000
1!
1%
#613350000000
0!
0%
#613355000000
1!
1%
#613360000000
0!
0%
#613365000000
1!
1%
#613370000000
0!
0%
#613375000000
1!
1%
#613380000000
0!
0%
#613385000000
1!
1%
#613390000000
0!
0%
#613395000000
1!
1%
#613400000000
0!
0%
#613405000000
1!
1%
#613410000000
0!
0%
#613415000000
1!
1%
#613420000000
0!
0%
#613425000000
1!
1%
#613430000000
0!
0%
#613435000000
1!
1%
#613440000000
0!
0%
#613445000000
1!
1%
#613450000000
0!
0%
#613455000000
1!
1%
#613460000000
0!
0%
#613465000000
1!
1%
#613470000000
0!
0%
#613475000000
1!
1%
#613480000000
0!
0%
#613485000000
1!
1%
#613490000000
0!
0%
#613495000000
1!
1%
#613500000000
0!
0%
#613505000000
1!
1%
#613510000000
0!
0%
#613515000000
1!
1%
#613520000000
0!
0%
#613525000000
1!
1%
#613530000000
0!
0%
#613535000000
1!
1%
#613540000000
0!
0%
#613545000000
1!
1%
#613550000000
0!
0%
#613555000000
1!
1%
#613560000000
0!
0%
#613565000000
1!
1%
#613570000000
0!
0%
#613575000000
1!
1%
#613580000000
0!
0%
#613585000000
1!
1%
#613590000000
0!
0%
#613595000000
1!
1%
#613600000000
0!
0%
#613605000000
1!
1%
#613610000000
0!
0%
#613615000000
1!
1%
#613620000000
0!
0%
#613625000000
1!
1%
#613630000000
0!
0%
#613635000000
1!
1%
#613640000000
0!
0%
#613645000000
1!
1%
#613650000000
0!
0%
#613655000000
1!
1%
#613660000000
0!
0%
#613665000000
1!
1%
#613670000000
0!
0%
#613675000000
1!
1%
#613680000000
0!
0%
#613685000000
1!
1%
#613690000000
0!
0%
#613695000000
1!
1%
#613700000000
0!
0%
#613705000000
1!
1%
#613710000000
0!
0%
#613715000000
1!
1%
#613720000000
0!
0%
#613725000000
1!
1%
#613730000000
0!
0%
#613735000000
1!
1%
#613740000000
0!
0%
#613745000000
1!
1%
#613750000000
0!
0%
#613755000000
1!
1%
#613760000000
0!
0%
#613765000000
1!
1%
#613770000000
0!
0%
#613775000000
1!
1%
#613780000000
0!
0%
#613785000000
1!
1%
#613790000000
0!
0%
#613795000000
1!
1%
#613800000000
0!
0%
#613805000000
1!
1%
#613810000000
0!
0%
#613815000000
1!
1%
#613820000000
0!
0%
#613825000000
1!
1%
#613830000000
0!
0%
#613835000000
1!
1%
#613840000000
0!
0%
#613845000000
1!
1%
#613850000000
0!
0%
#613855000000
1!
1%
#613860000000
0!
0%
#613865000000
1!
1%
#613870000000
0!
0%
#613875000000
1!
1%
#613880000000
0!
0%
#613885000000
1!
1%
#613890000000
0!
0%
#613895000000
1!
1%
#613900000000
0!
0%
#613905000000
1!
1%
#613910000000
0!
0%
#613915000000
1!
1%
#613920000000
0!
0%
#613925000000
1!
1%
#613930000000
0!
0%
#613935000000
1!
1%
#613940000000
0!
0%
#613945000000
1!
1%
#613950000000
0!
0%
#613955000000
1!
1%
#613960000000
0!
0%
#613965000000
1!
1%
#613970000000
0!
0%
#613975000000
1!
1%
#613980000000
0!
0%
#613985000000
1!
1%
#613990000000
0!
0%
#613995000000
1!
1%
#614000000000
0!
0%
#614005000000
1!
1%
#614010000000
0!
0%
#614015000000
1!
1%
#614020000000
0!
0%
#614025000000
1!
1%
#614030000000
0!
0%
#614035000000
1!
1%
#614040000000
0!
0%
#614045000000
1!
1%
#614050000000
0!
0%
#614055000000
1!
1%
#614060000000
0!
0%
#614065000000
1!
1%
#614070000000
0!
0%
#614075000000
1!
1%
#614080000000
0!
0%
#614085000000
1!
1%
#614090000000
0!
0%
#614095000000
1!
1%
#614100000000
0!
0%
#614105000000
1!
1%
#614110000000
0!
0%
#614115000000
1!
1%
#614120000000
0!
0%
#614125000000
1!
1%
#614130000000
0!
0%
#614135000000
1!
1%
#614140000000
0!
0%
#614145000000
1!
1%
#614150000000
0!
0%
#614155000000
1!
1%
#614160000000
0!
0%
#614165000000
1!
1%
#614170000000
0!
0%
#614175000000
1!
1%
#614180000000
0!
0%
#614185000000
1!
1%
#614190000000
0!
0%
#614195000000
1!
1%
#614200000000
0!
0%
#614205000000
1!
1%
#614210000000
0!
0%
#614215000000
1!
1%
#614220000000
0!
0%
#614225000000
1!
1%
#614230000000
0!
0%
#614235000000
1!
1%
#614240000000
0!
0%
#614245000000
1!
1%
#614250000000
0!
0%
#614255000000
1!
1%
#614260000000
0!
0%
#614265000000
1!
1%
#614270000000
0!
0%
#614275000000
1!
1%
#614280000000
0!
0%
#614285000000
1!
1%
#614290000000
0!
0%
#614295000000
1!
1%
#614300000000
0!
0%
#614305000000
1!
1%
#614310000000
0!
0%
#614315000000
1!
1%
#614320000000
0!
0%
#614325000000
1!
1%
#614330000000
0!
0%
#614335000000
1!
1%
#614340000000
0!
0%
#614345000000
1!
1%
#614350000000
0!
0%
#614355000000
1!
1%
#614360000000
0!
0%
#614365000000
1!
1%
#614370000000
0!
0%
#614375000000
1!
1%
#614380000000
0!
0%
#614385000000
1!
1%
#614390000000
0!
0%
#614395000000
1!
1%
#614400000000
0!
0%
#614405000000
1!
1%
#614410000000
0!
0%
#614415000000
1!
1%
#614420000000
0!
0%
#614425000000
1!
1%
#614430000000
0!
0%
#614435000000
1!
1%
#614440000000
0!
0%
#614445000000
1!
1%
#614450000000
0!
0%
#614455000000
1!
1%
#614460000000
0!
0%
#614465000000
1!
1%
#614470000000
0!
0%
#614475000000
1!
1%
#614480000000
0!
0%
#614485000000
1!
1%
#614490000000
0!
0%
#614495000000
1!
1%
#614500000000
0!
0%
#614505000000
1!
1%
#614510000000
0!
0%
#614515000000
1!
1%
#614520000000
0!
0%
#614525000000
1!
1%
#614530000000
0!
0%
#614535000000
1!
1%
#614540000000
0!
0%
#614545000000
1!
1%
#614550000000
0!
0%
#614555000000
1!
1%
#614560000000
0!
0%
#614565000000
1!
1%
#614570000000
0!
0%
#614575000000
1!
1%
#614580000000
0!
0%
#614585000000
1!
1%
#614590000000
0!
0%
#614595000000
1!
1%
#614600000000
0!
0%
#614605000000
1!
1%
#614610000000
0!
0%
#614615000000
1!
1%
#614620000000
0!
0%
#614625000000
1!
1%
#614630000000
0!
0%
#614635000000
1!
1%
#614640000000
0!
0%
#614645000000
1!
1%
#614650000000
0!
0%
#614655000000
1!
1%
#614660000000
0!
0%
#614665000000
1!
1%
#614670000000
0!
0%
#614675000000
1!
1%
#614680000000
0!
0%
#614685000000
1!
1%
#614690000000
0!
0%
#614695000000
1!
1%
#614700000000
0!
0%
#614705000000
1!
1%
#614710000000
0!
0%
#614715000000
1!
1%
#614720000000
0!
0%
#614725000000
1!
1%
#614730000000
0!
0%
#614735000000
1!
1%
#614740000000
0!
0%
#614745000000
1!
1%
#614750000000
0!
0%
#614755000000
1!
1%
#614760000000
0!
0%
#614765000000
1!
1%
#614770000000
0!
0%
#614775000000
1!
1%
#614780000000
0!
0%
#614785000000
1!
1%
#614790000000
0!
0%
#614795000000
1!
1%
#614800000000
0!
0%
#614805000000
1!
1%
#614810000000
0!
0%
#614815000000
1!
1%
#614820000000
0!
0%
#614825000000
1!
1%
#614830000000
0!
0%
#614835000000
1!
1%
#614840000000
0!
0%
#614845000000
1!
1%
#614850000000
0!
0%
#614855000000
1!
1%
#614860000000
0!
0%
#614865000000
1!
1%
#614870000000
0!
0%
#614875000000
1!
1%
#614880000000
0!
0%
#614885000000
1!
1%
#614890000000
0!
0%
#614895000000
1!
1%
#614900000000
0!
0%
#614905000000
1!
1%
#614910000000
0!
0%
#614915000000
1!
1%
#614920000000
0!
0%
#614925000000
1!
1%
#614930000000
0!
0%
#614935000000
1!
1%
#614940000000
0!
0%
#614945000000
1!
1%
#614950000000
0!
0%
#614955000000
1!
1%
#614960000000
0!
0%
#614965000000
1!
1%
#614970000000
0!
0%
#614975000000
1!
1%
#614980000000
0!
0%
#614985000000
1!
1%
#614990000000
0!
0%
#614995000000
1!
1%
#615000000000
0!
0%
#615005000000
1!
1%
#615010000000
0!
0%
#615015000000
1!
1%
#615020000000
0!
0%
#615025000000
1!
1%
#615030000000
0!
0%
#615035000000
1!
1%
#615040000000
0!
0%
#615045000000
1!
1%
#615050000000
0!
0%
#615055000000
1!
1%
#615060000000
0!
0%
#615065000000
1!
1%
#615070000000
0!
0%
#615075000000
1!
1%
#615080000000
0!
0%
#615085000000
1!
1%
#615090000000
0!
0%
#615095000000
1!
1%
#615100000000
0!
0%
#615105000000
1!
1%
#615110000000
0!
0%
#615115000000
1!
1%
#615120000000
0!
0%
#615125000000
1!
1%
#615130000000
0!
0%
#615135000000
1!
1%
#615140000000
0!
0%
#615145000000
1!
1%
#615150000000
0!
0%
#615155000000
1!
1%
#615160000000
0!
0%
#615165000000
1!
1%
#615170000000
0!
0%
#615175000000
1!
1%
#615180000000
0!
0%
#615185000000
1!
1%
#615190000000
0!
0%
#615195000000
1!
1%
#615200000000
0!
0%
#615205000000
1!
1%
#615210000000
0!
0%
#615215000000
1!
1%
#615220000000
0!
0%
#615225000000
1!
1%
#615230000000
0!
0%
#615235000000
1!
1%
#615240000000
0!
0%
#615245000000
1!
1%
#615250000000
0!
0%
#615255000000
1!
1%
#615260000000
0!
0%
#615265000000
1!
1%
#615270000000
0!
0%
#615275000000
1!
1%
#615280000000
0!
0%
#615285000000
1!
1%
#615290000000
0!
0%
#615295000000
1!
1%
#615300000000
0!
0%
#615305000000
1!
1%
#615310000000
0!
0%
#615315000000
1!
1%
#615320000000
0!
0%
#615325000000
1!
1%
#615330000000
0!
0%
#615335000000
1!
1%
#615340000000
0!
0%
#615345000000
1!
1%
#615350000000
0!
0%
#615355000000
1!
1%
#615360000000
0!
0%
#615365000000
1!
1%
#615370000000
0!
0%
#615375000000
1!
1%
#615380000000
0!
0%
#615385000000
1!
1%
#615390000000
0!
0%
#615395000000
1!
1%
#615400000000
0!
0%
#615405000000
1!
1%
#615410000000
0!
0%
#615415000000
1!
1%
#615420000000
0!
0%
#615425000000
1!
1%
#615430000000
0!
0%
#615435000000
1!
1%
#615440000000
0!
0%
#615445000000
1!
1%
#615450000000
0!
0%
#615455000000
1!
1%
#615460000000
0!
0%
#615465000000
1!
1%
#615470000000
0!
0%
#615475000000
1!
1%
#615480000000
0!
0%
#615485000000
1!
1%
#615490000000
0!
0%
#615495000000
1!
1%
#615500000000
0!
0%
#615505000000
1!
1%
#615510000000
0!
0%
#615515000000
1!
1%
#615520000000
0!
0%
#615525000000
1!
1%
#615530000000
0!
0%
#615535000000
1!
1%
#615540000000
0!
0%
#615545000000
1!
1%
#615550000000
0!
0%
#615555000000
1!
1%
#615560000000
0!
0%
#615565000000
1!
1%
#615570000000
0!
0%
#615575000000
1!
1%
#615580000000
0!
0%
#615585000000
1!
1%
#615590000000
0!
0%
#615595000000
1!
1%
#615600000000
0!
0%
#615605000000
1!
1%
#615610000000
0!
0%
#615615000000
1!
1%
#615620000000
0!
0%
#615625000000
1!
1%
#615630000000
0!
0%
#615635000000
1!
1%
#615640000000
0!
0%
#615645000000
1!
1%
#615650000000
0!
0%
#615655000000
1!
1%
#615660000000
0!
0%
#615665000000
1!
1%
#615670000000
0!
0%
#615675000000
1!
1%
#615680000000
0!
0%
#615685000000
1!
1%
#615690000000
0!
0%
#615695000000
1!
1%
#615700000000
0!
0%
#615705000000
1!
1%
#615710000000
0!
0%
#615715000000
1!
1%
#615720000000
0!
0%
#615725000000
1!
1%
#615730000000
0!
0%
#615735000000
1!
1%
#615740000000
0!
0%
#615745000000
1!
1%
#615750000000
0!
0%
#615755000000
1!
1%
#615760000000
0!
0%
#615765000000
1!
1%
#615770000000
0!
0%
#615775000000
1!
1%
#615780000000
0!
0%
#615785000000
1!
1%
#615790000000
0!
0%
#615795000000
1!
1%
#615800000000
0!
0%
#615805000000
1!
1%
#615810000000
0!
0%
#615815000000
1!
1%
#615820000000
0!
0%
#615825000000
1!
1%
#615830000000
0!
0%
#615835000000
1!
1%
#615840000000
0!
0%
#615845000000
1!
1%
#615850000000
0!
0%
#615855000000
1!
1%
#615860000000
0!
0%
#615865000000
1!
1%
#615870000000
0!
0%
#615875000000
1!
1%
#615880000000
0!
0%
#615885000000
1!
1%
#615890000000
0!
0%
#615895000000
1!
1%
#615900000000
0!
0%
#615905000000
1!
1%
#615910000000
0!
0%
#615915000000
1!
1%
#615920000000
0!
0%
#615925000000
1!
1%
#615930000000
0!
0%
#615935000000
1!
1%
#615940000000
0!
0%
#615945000000
1!
1%
#615950000000
0!
0%
#615955000000
1!
1%
#615960000000
0!
0%
#615965000000
1!
1%
#615970000000
0!
0%
#615975000000
1!
1%
#615980000000
0!
0%
#615985000000
1!
1%
#615990000000
0!
0%
#615995000000
1!
1%
#616000000000
0!
0%
#616005000000
1!
1%
#616010000000
0!
0%
#616015000000
1!
1%
#616020000000
0!
0%
#616025000000
1!
1%
#616030000000
0!
0%
#616035000000
1!
1%
#616040000000
0!
0%
#616045000000
1!
1%
#616050000000
0!
0%
#616055000000
1!
1%
#616060000000
0!
0%
#616065000000
1!
1%
#616070000000
0!
0%
#616075000000
1!
1%
#616080000000
0!
0%
#616085000000
1!
1%
#616090000000
0!
0%
#616095000000
1!
1%
#616100000000
0!
0%
#616105000000
1!
1%
#616110000000
0!
0%
#616115000000
1!
1%
#616120000000
0!
0%
#616125000000
1!
1%
#616130000000
0!
0%
#616135000000
1!
1%
#616140000000
0!
0%
#616145000000
1!
1%
#616150000000
0!
0%
#616155000000
1!
1%
#616160000000
0!
0%
#616165000000
1!
1%
#616170000000
0!
0%
#616175000000
1!
1%
#616180000000
0!
0%
#616185000000
1!
1%
#616190000000
0!
0%
#616195000000
1!
1%
#616200000000
0!
0%
#616205000000
1!
1%
#616210000000
0!
0%
#616215000000
1!
1%
#616220000000
0!
0%
#616225000000
1!
1%
#616230000000
0!
0%
#616235000000
1!
1%
#616240000000
0!
0%
#616245000000
1!
1%
#616250000000
0!
0%
#616255000000
1!
1%
#616260000000
0!
0%
#616265000000
1!
1%
#616270000000
0!
0%
#616275000000
1!
1%
#616280000000
0!
0%
#616285000000
1!
1%
#616290000000
0!
0%
#616295000000
1!
1%
#616300000000
0!
0%
#616305000000
1!
1%
#616310000000
0!
0%
#616315000000
1!
1%
#616320000000
0!
0%
#616325000000
1!
1%
#616330000000
0!
0%
#616335000000
1!
1%
#616340000000
0!
0%
#616345000000
1!
1%
#616350000000
0!
0%
#616355000000
1!
1%
#616360000000
0!
0%
#616365000000
1!
1%
#616370000000
0!
0%
#616375000000
1!
1%
#616380000000
0!
0%
#616385000000
1!
1%
#616390000000
0!
0%
#616395000000
1!
1%
#616400000000
0!
0%
#616405000000
1!
1%
#616410000000
0!
0%
#616415000000
1!
1%
#616420000000
0!
0%
#616425000000
1!
1%
#616430000000
0!
0%
#616435000000
1!
1%
#616440000000
0!
0%
#616445000000
1!
1%
#616450000000
0!
0%
#616455000000
1!
1%
#616460000000
0!
0%
#616465000000
1!
1%
#616470000000
0!
0%
#616475000000
1!
1%
#616480000000
0!
0%
#616485000000
1!
1%
#616490000000
0!
0%
#616495000000
1!
1%
#616500000000
0!
0%
#616505000000
1!
1%
#616510000000
0!
0%
#616515000000
1!
1%
#616520000000
0!
0%
#616525000000
1!
1%
#616530000000
0!
0%
#616535000000
1!
1%
#616540000000
0!
0%
#616545000000
1!
1%
#616550000000
0!
0%
#616555000000
1!
1%
#616560000000
0!
0%
#616565000000
1!
1%
#616570000000
0!
0%
#616575000000
1!
1%
#616580000000
0!
0%
#616585000000
1!
1%
#616590000000
0!
0%
#616595000000
1!
1%
#616600000000
0!
0%
#616605000000
1!
1%
#616610000000
0!
0%
#616615000000
1!
1%
#616620000000
0!
0%
#616625000000
1!
1%
#616630000000
0!
0%
#616635000000
1!
1%
#616640000000
0!
0%
#616645000000
1!
1%
#616650000000
0!
0%
#616655000000
1!
1%
#616660000000
0!
0%
#616665000000
1!
1%
#616670000000
0!
0%
#616675000000
1!
1%
#616680000000
0!
0%
#616685000000
1!
1%
#616690000000
0!
0%
#616695000000
1!
1%
#616700000000
0!
0%
#616705000000
1!
1%
#616710000000
0!
0%
#616715000000
1!
1%
#616720000000
0!
0%
#616725000000
1!
1%
#616730000000
0!
0%
#616735000000
1!
1%
#616740000000
0!
0%
#616745000000
1!
1%
#616750000000
0!
0%
#616755000000
1!
1%
#616760000000
0!
0%
#616765000000
1!
1%
#616770000000
0!
0%
#616775000000
1!
1%
#616780000000
0!
0%
#616785000000
1!
1%
#616790000000
0!
0%
#616795000000
1!
1%
#616800000000
0!
0%
#616805000000
1!
1%
#616810000000
0!
0%
#616815000000
1!
1%
#616820000000
0!
0%
#616825000000
1!
1%
#616830000000
0!
0%
#616835000000
1!
1%
#616840000000
0!
0%
#616845000000
1!
1%
#616850000000
0!
0%
#616855000000
1!
1%
#616860000000
0!
0%
#616865000000
1!
1%
#616870000000
0!
0%
#616875000000
1!
1%
#616880000000
0!
0%
#616885000000
1!
1%
#616890000000
0!
0%
#616895000000
1!
1%
#616900000000
0!
0%
#616905000000
1!
1%
#616910000000
0!
0%
#616915000000
1!
1%
#616920000000
0!
0%
#616925000000
1!
1%
#616930000000
0!
0%
#616935000000
1!
1%
#616940000000
0!
0%
#616945000000
1!
1%
#616950000000
0!
0%
#616955000000
1!
1%
#616960000000
0!
0%
#616965000000
1!
1%
#616970000000
0!
0%
#616975000000
1!
1%
#616980000000
0!
0%
#616985000000
1!
1%
#616990000000
0!
0%
#616995000000
1!
1%
#617000000000
0!
0%
#617005000000
1!
1%
#617010000000
0!
0%
#617015000000
1!
1%
#617020000000
0!
0%
#617025000000
1!
1%
#617030000000
0!
0%
#617035000000
1!
1%
#617040000000
0!
0%
#617045000000
1!
1%
#617050000000
0!
0%
#617055000000
1!
1%
#617060000000
0!
0%
#617065000000
1!
1%
#617070000000
0!
0%
#617075000000
1!
1%
#617080000000
0!
0%
#617085000000
1!
1%
#617090000000
0!
0%
#617095000000
1!
1%
#617100000000
0!
0%
#617105000000
1!
1%
#617110000000
0!
0%
#617115000000
1!
1%
#617120000000
0!
0%
#617125000000
1!
1%
#617130000000
0!
0%
#617135000000
1!
1%
#617140000000
0!
0%
#617145000000
1!
1%
#617150000000
0!
0%
#617155000000
1!
1%
#617160000000
0!
0%
#617165000000
1!
1%
#617170000000
0!
0%
#617175000000
1!
1%
#617180000000
0!
0%
#617185000000
1!
1%
#617190000000
0!
0%
#617195000000
1!
1%
#617200000000
0!
0%
#617205000000
1!
1%
#617210000000
0!
0%
#617215000000
1!
1%
#617220000000
0!
0%
#617225000000
1!
1%
#617230000000
0!
0%
#617235000000
1!
1%
#617240000000
0!
0%
#617245000000
1!
1%
#617250000000
0!
0%
#617255000000
1!
1%
#617260000000
0!
0%
#617265000000
1!
1%
#617270000000
0!
0%
#617275000000
1!
1%
#617280000000
0!
0%
#617285000000
1!
1%
#617290000000
0!
0%
#617295000000
1!
1%
#617300000000
0!
0%
#617305000000
1!
1%
#617310000000
0!
0%
#617315000000
1!
1%
#617320000000
0!
0%
#617325000000
1!
1%
#617330000000
0!
0%
#617335000000
1!
1%
#617340000000
0!
0%
#617345000000
1!
1%
#617350000000
0!
0%
#617355000000
1!
1%
#617360000000
0!
0%
#617365000000
1!
1%
#617370000000
0!
0%
#617375000000
1!
1%
#617380000000
0!
0%
#617385000000
1!
1%
#617390000000
0!
0%
#617395000000
1!
1%
#617400000000
0!
0%
#617405000000
1!
1%
#617410000000
0!
0%
#617415000000
1!
1%
#617420000000
0!
0%
#617425000000
1!
1%
#617430000000
0!
0%
#617435000000
1!
1%
#617440000000
0!
0%
#617445000000
1!
1%
#617450000000
0!
0%
#617455000000
1!
1%
#617460000000
0!
0%
#617465000000
1!
1%
#617470000000
0!
0%
#617475000000
1!
1%
#617480000000
0!
0%
#617485000000
1!
1%
#617490000000
0!
0%
#617495000000
1!
1%
#617500000000
0!
0%
#617505000000
1!
1%
#617510000000
0!
0%
#617515000000
1!
1%
#617520000000
0!
0%
#617525000000
1!
1%
#617530000000
0!
0%
#617535000000
1!
1%
#617540000000
0!
0%
#617545000000
1!
1%
#617550000000
0!
0%
#617555000000
1!
1%
#617560000000
0!
0%
#617565000000
1!
1%
#617570000000
0!
0%
#617575000000
1!
1%
#617580000000
0!
0%
#617585000000
1!
1%
#617590000000
0!
0%
#617595000000
1!
1%
#617600000000
0!
0%
#617605000000
1!
1%
#617610000000
0!
0%
#617615000000
1!
1%
#617620000000
0!
0%
#617625000000
1!
1%
#617630000000
0!
0%
#617635000000
1!
1%
#617640000000
0!
0%
#617645000000
1!
1%
#617650000000
0!
0%
#617655000000
1!
1%
#617660000000
0!
0%
#617665000000
1!
1%
#617670000000
0!
0%
#617675000000
1!
1%
#617680000000
0!
0%
#617685000000
1!
1%
#617690000000
0!
0%
#617695000000
1!
1%
#617700000000
0!
0%
#617705000000
1!
1%
#617710000000
0!
0%
#617715000000
1!
1%
#617720000000
0!
0%
#617725000000
1!
1%
#617730000000
0!
0%
#617735000000
1!
1%
#617740000000
0!
0%
#617745000000
1!
1%
#617750000000
0!
0%
#617755000000
1!
1%
#617760000000
0!
0%
#617765000000
1!
1%
#617770000000
0!
0%
#617775000000
1!
1%
#617780000000
0!
0%
#617785000000
1!
1%
#617790000000
0!
0%
#617795000000
1!
1%
#617800000000
0!
0%
#617805000000
1!
1%
#617810000000
0!
0%
#617815000000
1!
1%
#617820000000
0!
0%
#617825000000
1!
1%
#617830000000
0!
0%
#617835000000
1!
1%
#617840000000
0!
0%
#617845000000
1!
1%
#617850000000
0!
0%
#617855000000
1!
1%
#617860000000
0!
0%
#617865000000
1!
1%
#617870000000
0!
0%
#617875000000
1!
1%
#617880000000
0!
0%
#617885000000
1!
1%
#617890000000
0!
0%
#617895000000
1!
1%
#617900000000
0!
0%
#617905000000
1!
1%
#617910000000
0!
0%
#617915000000
1!
1%
#617920000000
0!
0%
#617925000000
1!
1%
#617930000000
0!
0%
#617935000000
1!
1%
#617940000000
0!
0%
#617945000000
1!
1%
#617950000000
0!
0%
#617955000000
1!
1%
#617960000000
0!
0%
#617965000000
1!
1%
#617970000000
0!
0%
#617975000000
1!
1%
#617980000000
0!
0%
#617985000000
1!
1%
#617990000000
0!
0%
#617995000000
1!
1%
#618000000000
0!
0%
#618005000000
1!
1%
#618010000000
0!
0%
#618015000000
1!
1%
#618020000000
0!
0%
#618025000000
1!
1%
#618030000000
0!
0%
#618035000000
1!
1%
#618040000000
0!
0%
#618045000000
1!
1%
#618050000000
0!
0%
#618055000000
1!
1%
#618060000000
0!
0%
#618065000000
1!
1%
#618070000000
0!
0%
#618075000000
1!
1%
#618080000000
0!
0%
#618085000000
1!
1%
#618090000000
0!
0%
#618095000000
1!
1%
#618100000000
0!
0%
#618105000000
1!
1%
#618110000000
0!
0%
#618115000000
1!
1%
#618120000000
0!
0%
#618125000000
1!
1%
#618130000000
0!
0%
#618135000000
1!
1%
#618140000000
0!
0%
#618145000000
1!
1%
#618150000000
0!
0%
#618155000000
1!
1%
#618160000000
0!
0%
#618165000000
1!
1%
#618170000000
0!
0%
#618175000000
1!
1%
#618180000000
0!
0%
#618185000000
1!
1%
#618190000000
0!
0%
#618195000000
1!
1%
#618200000000
0!
0%
#618205000000
1!
1%
#618210000000
0!
0%
#618215000000
1!
1%
#618220000000
0!
0%
#618225000000
1!
1%
#618230000000
0!
0%
#618235000000
1!
1%
#618240000000
0!
0%
#618245000000
1!
1%
#618250000000
0!
0%
#618255000000
1!
1%
#618260000000
0!
0%
#618265000000
1!
1%
#618270000000
0!
0%
#618275000000
1!
1%
#618280000000
0!
0%
#618285000000
1!
1%
#618290000000
0!
0%
#618295000000
1!
1%
#618300000000
0!
0%
#618305000000
1!
1%
#618310000000
0!
0%
#618315000000
1!
1%
#618320000000
0!
0%
#618325000000
1!
1%
#618330000000
0!
0%
#618335000000
1!
1%
#618340000000
0!
0%
#618345000000
1!
1%
#618350000000
0!
0%
#618355000000
1!
1%
#618360000000
0!
0%
#618365000000
1!
1%
#618370000000
0!
0%
#618375000000
1!
1%
#618380000000
0!
0%
#618385000000
1!
1%
#618390000000
0!
0%
#618395000000
1!
1%
#618400000000
0!
0%
#618405000000
1!
1%
#618410000000
0!
0%
#618415000000
1!
1%
#618420000000
0!
0%
#618425000000
1!
1%
#618430000000
0!
0%
#618435000000
1!
1%
#618440000000
0!
0%
#618445000000
1!
1%
#618450000000
0!
0%
#618455000000
1!
1%
#618460000000
0!
0%
#618465000000
1!
1%
#618470000000
0!
0%
#618475000000
1!
1%
#618480000000
0!
0%
#618485000000
1!
1%
#618490000000
0!
0%
#618495000000
1!
1%
#618500000000
0!
0%
#618505000000
1!
1%
#618510000000
0!
0%
#618515000000
1!
1%
#618520000000
0!
0%
#618525000000
1!
1%
#618530000000
0!
0%
#618535000000
1!
1%
#618540000000
0!
0%
#618545000000
1!
1%
#618550000000
0!
0%
#618555000000
1!
1%
#618560000000
0!
0%
#618565000000
1!
1%
#618570000000
0!
0%
#618575000000
1!
1%
#618580000000
0!
0%
#618585000000
1!
1%
#618590000000
0!
0%
#618595000000
1!
1%
#618600000000
0!
0%
#618605000000
1!
1%
#618610000000
0!
0%
#618615000000
1!
1%
#618620000000
0!
0%
#618625000000
1!
1%
#618630000000
0!
0%
#618635000000
1!
1%
#618640000000
0!
0%
#618645000000
1!
1%
#618650000000
0!
0%
#618655000000
1!
1%
#618660000000
0!
0%
#618665000000
1!
1%
#618670000000
0!
0%
#618675000000
1!
1%
#618680000000
0!
0%
#618685000000
1!
1%
#618690000000
0!
0%
#618695000000
1!
1%
#618700000000
0!
0%
#618705000000
1!
1%
#618710000000
0!
0%
#618715000000
1!
1%
#618720000000
0!
0%
#618725000000
1!
1%
#618730000000
0!
0%
#618735000000
1!
1%
#618740000000
0!
0%
#618745000000
1!
1%
#618750000000
0!
0%
#618755000000
1!
1%
#618760000000
0!
0%
#618765000000
1!
1%
#618770000000
0!
0%
#618775000000
1!
1%
#618780000000
0!
0%
#618785000000
1!
1%
#618790000000
0!
0%
#618795000000
1!
1%
#618800000000
0!
0%
#618805000000
1!
1%
#618810000000
0!
0%
#618815000000
1!
1%
#618820000000
0!
0%
#618825000000
1!
1%
#618830000000
0!
0%
#618835000000
1!
1%
#618840000000
0!
0%
#618845000000
1!
1%
#618850000000
0!
0%
#618855000000
1!
1%
#618860000000
0!
0%
#618865000000
1!
1%
#618870000000
0!
0%
#618875000000
1!
1%
#618880000000
0!
0%
#618885000000
1!
1%
#618890000000
0!
0%
#618895000000
1!
1%
#618900000000
0!
0%
#618905000000
1!
1%
#618910000000
0!
0%
#618915000000
1!
1%
#618920000000
0!
0%
#618925000000
1!
1%
#618930000000
0!
0%
#618935000000
1!
1%
#618940000000
0!
0%
#618945000000
1!
1%
#618950000000
0!
0%
#618955000000
1!
1%
#618960000000
0!
0%
#618965000000
1!
1%
#618970000000
0!
0%
#618975000000
1!
1%
#618980000000
0!
0%
#618985000000
1!
1%
#618990000000
0!
0%
#618995000000
1!
1%
#619000000000
0!
0%
#619005000000
1!
1%
#619010000000
0!
0%
#619015000000
1!
1%
#619020000000
0!
0%
#619025000000
1!
1%
#619030000000
0!
0%
#619035000000
1!
1%
#619040000000
0!
0%
#619045000000
1!
1%
#619050000000
0!
0%
#619055000000
1!
1%
#619060000000
0!
0%
#619065000000
1!
1%
#619070000000
0!
0%
#619075000000
1!
1%
#619080000000
0!
0%
#619085000000
1!
1%
#619090000000
0!
0%
#619095000000
1!
1%
#619100000000
0!
0%
#619105000000
1!
1%
#619110000000
0!
0%
#619115000000
1!
1%
#619120000000
0!
0%
#619125000000
1!
1%
#619130000000
0!
0%
#619135000000
1!
1%
#619140000000
0!
0%
#619145000000
1!
1%
#619150000000
0!
0%
#619155000000
1!
1%
#619160000000
0!
0%
#619165000000
1!
1%
#619170000000
0!
0%
#619175000000
1!
1%
#619180000000
0!
0%
#619185000000
1!
1%
#619190000000
0!
0%
#619195000000
1!
1%
#619200000000
0!
0%
#619205000000
1!
1%
#619210000000
0!
0%
#619215000000
1!
1%
#619220000000
0!
0%
#619225000000
1!
1%
#619230000000
0!
0%
#619235000000
1!
1%
#619240000000
0!
0%
#619245000000
1!
1%
#619250000000
0!
0%
#619255000000
1!
1%
#619260000000
0!
0%
#619265000000
1!
1%
#619270000000
0!
0%
#619275000000
1!
1%
#619280000000
0!
0%
#619285000000
1!
1%
#619290000000
0!
0%
#619295000000
1!
1%
#619300000000
0!
0%
#619305000000
1!
1%
#619310000000
0!
0%
#619315000000
1!
1%
#619320000000
0!
0%
#619325000000
1!
1%
#619330000000
0!
0%
#619335000000
1!
1%
#619340000000
0!
0%
#619345000000
1!
1%
#619350000000
0!
0%
#619355000000
1!
1%
#619360000000
0!
0%
#619365000000
1!
1%
#619370000000
0!
0%
#619375000000
1!
1%
#619380000000
0!
0%
#619385000000
1!
1%
#619390000000
0!
0%
#619395000000
1!
1%
#619400000000
0!
0%
#619405000000
1!
1%
#619410000000
0!
0%
#619415000000
1!
1%
#619420000000
0!
0%
#619425000000
1!
1%
#619430000000
0!
0%
#619435000000
1!
1%
#619440000000
0!
0%
#619445000000
1!
1%
#619450000000
0!
0%
#619455000000
1!
1%
#619460000000
0!
0%
#619465000000
1!
1%
#619470000000
0!
0%
#619475000000
1!
1%
#619480000000
0!
0%
#619485000000
1!
1%
#619490000000
0!
0%
#619495000000
1!
1%
#619500000000
0!
0%
#619505000000
1!
1%
#619510000000
0!
0%
#619515000000
1!
1%
#619520000000
0!
0%
#619525000000
1!
1%
#619530000000
0!
0%
#619535000000
1!
1%
#619540000000
0!
0%
#619545000000
1!
1%
#619550000000
0!
0%
#619555000000
1!
1%
#619560000000
0!
0%
#619565000000
1!
1%
#619570000000
0!
0%
#619575000000
1!
1%
#619580000000
0!
0%
#619585000000
1!
1%
#619590000000
0!
0%
#619595000000
1!
1%
#619600000000
0!
0%
#619605000000
1!
1%
#619610000000
0!
0%
#619615000000
1!
1%
#619620000000
0!
0%
#619625000000
1!
1%
#619630000000
0!
0%
#619635000000
1!
1%
#619640000000
0!
0%
#619645000000
1!
1%
#619650000000
0!
0%
#619655000000
1!
1%
#619660000000
0!
0%
#619665000000
1!
1%
#619670000000
0!
0%
#619675000000
1!
1%
#619680000000
0!
0%
#619685000000
1!
1%
#619690000000
0!
0%
#619695000000
1!
1%
#619700000000
0!
0%
#619705000000
1!
1%
#619710000000
0!
0%
#619715000000
1!
1%
#619720000000
0!
0%
#619725000000
1!
1%
#619730000000
0!
0%
#619735000000
1!
1%
#619740000000
0!
0%
#619745000000
1!
1%
#619750000000
0!
0%
#619755000000
1!
1%
#619760000000
0!
0%
#619765000000
1!
1%
#619770000000
0!
0%
#619775000000
1!
1%
#619780000000
0!
0%
#619785000000
1!
1%
#619790000000
0!
0%
#619795000000
1!
1%
#619800000000
0!
0%
#619805000000
1!
1%
#619810000000
0!
0%
#619815000000
1!
1%
#619820000000
0!
0%
#619825000000
1!
1%
#619830000000
0!
0%
#619835000000
1!
1%
#619840000000
0!
0%
#619845000000
1!
1%
#619850000000
0!
0%
#619855000000
1!
1%
#619860000000
0!
0%
#619865000000
1!
1%
#619870000000
0!
0%
#619875000000
1!
1%
#619880000000
0!
0%
#619885000000
1!
1%
#619890000000
0!
0%
#619895000000
1!
1%
#619900000000
0!
0%
#619905000000
1!
1%
#619910000000
0!
0%
#619915000000
1!
1%
#619920000000
0!
0%
#619925000000
1!
1%
#619930000000
0!
0%
#619935000000
1!
1%
#619940000000
0!
0%
#619945000000
1!
1%
#619950000000
0!
0%
#619955000000
1!
1%
#619960000000
0!
0%
#619965000000
1!
1%
#619970000000
0!
0%
#619975000000
1!
1%
#619980000000
0!
0%
#619985000000
1!
1%
#619990000000
0!
0%
#619995000000
1!
1%
#620000000000
0!
0%
#620005000000
1!
1%
#620010000000
0!
0%
#620015000000
1!
1%
#620020000000
0!
0%
#620025000000
1!
1%
#620030000000
0!
0%
#620035000000
1!
1%
#620040000000
0!
0%
#620045000000
1!
1%
#620050000000
0!
0%
#620055000000
1!
1%
#620060000000
0!
0%
#620065000000
1!
1%
#620070000000
0!
0%
#620075000000
1!
1%
#620080000000
0!
0%
#620085000000
1!
1%
#620090000000
0!
0%
#620095000000
1!
1%
#620100000000
0!
0%
#620105000000
1!
1%
#620110000000
0!
0%
#620115000000
1!
1%
#620120000000
0!
0%
#620125000000
1!
1%
#620130000000
0!
0%
#620135000000
1!
1%
#620140000000
0!
0%
#620145000000
1!
1%
#620150000000
0!
0%
#620155000000
1!
1%
#620160000000
0!
0%
#620165000000
1!
1%
#620170000000
0!
0%
#620175000000
1!
1%
#620180000000
0!
0%
#620185000000
1!
1%
#620190000000
0!
0%
#620195000000
1!
1%
#620200000000
0!
0%
#620205000000
1!
1%
#620210000000
0!
0%
#620215000000
1!
1%
#620220000000
0!
0%
#620225000000
1!
1%
#620230000000
0!
0%
#620235000000
1!
1%
#620240000000
0!
0%
#620245000000
1!
1%
#620250000000
0!
0%
#620255000000
1!
1%
#620260000000
0!
0%
#620265000000
1!
1%
#620270000000
0!
0%
#620275000000
1!
1%
#620280000000
0!
0%
#620285000000
1!
1%
#620290000000
0!
0%
#620295000000
1!
1%
#620300000000
0!
0%
#620305000000
1!
1%
#620310000000
0!
0%
#620315000000
1!
1%
#620320000000
0!
0%
#620325000000
1!
1%
#620330000000
0!
0%
#620335000000
1!
1%
#620340000000
0!
0%
#620345000000
1!
1%
#620350000000
0!
0%
#620355000000
1!
1%
#620360000000
0!
0%
#620365000000
1!
1%
#620370000000
0!
0%
#620375000000
1!
1%
#620380000000
0!
0%
#620385000000
1!
1%
#620390000000
0!
0%
#620395000000
1!
1%
#620400000000
0!
0%
#620405000000
1!
1%
#620410000000
0!
0%
#620415000000
1!
1%
#620420000000
0!
0%
#620425000000
1!
1%
#620430000000
0!
0%
#620435000000
1!
1%
#620440000000
0!
0%
#620445000000
1!
1%
#620450000000
0!
0%
#620455000000
1!
1%
#620460000000
0!
0%
#620465000000
1!
1%
#620470000000
0!
0%
#620475000000
1!
1%
#620480000000
0!
0%
#620485000000
1!
1%
#620490000000
0!
0%
#620495000000
1!
1%
#620500000000
0!
0%
#620505000000
1!
1%
#620510000000
0!
0%
#620515000000
1!
1%
#620520000000
0!
0%
#620525000000
1!
1%
#620530000000
0!
0%
#620535000000
1!
1%
#620540000000
0!
0%
#620545000000
1!
1%
#620550000000
0!
0%
#620555000000
1!
1%
#620560000000
0!
0%
#620565000000
1!
1%
#620570000000
0!
0%
#620575000000
1!
1%
#620580000000
0!
0%
#620585000000
1!
1%
#620590000000
0!
0%
#620595000000
1!
1%
#620600000000
0!
0%
#620605000000
1!
1%
#620610000000
0!
0%
#620615000000
1!
1%
#620620000000
0!
0%
#620625000000
1!
1%
#620630000000
0!
0%
#620635000000
1!
1%
#620640000000
0!
0%
#620645000000
1!
1%
#620650000000
0!
0%
#620655000000
1!
1%
#620660000000
0!
0%
#620665000000
1!
1%
#620670000000
0!
0%
#620675000000
1!
1%
#620680000000
0!
0%
#620685000000
1!
1%
#620690000000
0!
0%
#620695000000
1!
1%
#620700000000
0!
0%
#620705000000
1!
1%
#620710000000
0!
0%
#620715000000
1!
1%
#620720000000
0!
0%
#620725000000
1!
1%
#620730000000
0!
0%
#620735000000
1!
1%
#620740000000
0!
0%
#620745000000
1!
1%
#620750000000
0!
0%
#620755000000
1!
1%
#620760000000
0!
0%
#620765000000
1!
1%
#620770000000
0!
0%
#620775000000
1!
1%
#620780000000
0!
0%
#620785000000
1!
1%
#620790000000
0!
0%
#620795000000
1!
1%
#620800000000
0!
0%
#620805000000
1!
1%
#620810000000
0!
0%
#620815000000
1!
1%
#620820000000
0!
0%
#620825000000
1!
1%
#620830000000
0!
0%
#620835000000
1!
1%
#620840000000
0!
0%
#620845000000
1!
1%
#620850000000
0!
0%
#620855000000
1!
1%
#620860000000
0!
0%
#620865000000
1!
1%
#620870000000
0!
0%
#620875000000
1!
1%
#620880000000
0!
0%
#620885000000
1!
1%
#620890000000
0!
0%
#620895000000
1!
1%
#620900000000
0!
0%
#620905000000
1!
1%
#620910000000
0!
0%
#620915000000
1!
1%
#620920000000
0!
0%
#620925000000
1!
1%
#620930000000
0!
0%
#620935000000
1!
1%
#620940000000
0!
0%
#620945000000
1!
1%
#620950000000
0!
0%
#620955000000
1!
1%
#620960000000
0!
0%
#620965000000
1!
1%
#620970000000
0!
0%
#620975000000
1!
1%
#620980000000
0!
0%
#620985000000
1!
1%
#620990000000
0!
0%
#620995000000
1!
1%
#621000000000
0!
0%
#621005000000
1!
1%
#621010000000
0!
0%
#621015000000
1!
1%
#621020000000
0!
0%
#621025000000
1!
1%
#621030000000
0!
0%
#621035000000
1!
1%
#621040000000
0!
0%
#621045000000
1!
1%
#621050000000
0!
0%
#621055000000
1!
1%
#621060000000
0!
0%
#621065000000
1!
1%
#621070000000
0!
0%
#621075000000
1!
1%
#621080000000
0!
0%
#621085000000
1!
1%
#621090000000
0!
0%
#621095000000
1!
1%
#621100000000
0!
0%
#621105000000
1!
1%
#621110000000
0!
0%
#621115000000
1!
1%
#621120000000
0!
0%
#621125000000
1!
1%
#621130000000
0!
0%
#621135000000
1!
1%
#621140000000
0!
0%
#621145000000
1!
1%
#621150000000
0!
0%
#621155000000
1!
1%
#621160000000
0!
0%
#621165000000
1!
1%
#621170000000
0!
0%
#621175000000
1!
1%
#621180000000
0!
0%
#621185000000
1!
1%
#621190000000
0!
0%
#621195000000
1!
1%
#621200000000
0!
0%
#621205000000
1!
1%
#621210000000
0!
0%
#621215000000
1!
1%
#621220000000
0!
0%
#621225000000
1!
1%
#621230000000
0!
0%
#621235000000
1!
1%
#621240000000
0!
0%
#621245000000
1!
1%
#621250000000
0!
0%
#621255000000
1!
1%
#621260000000
0!
0%
#621265000000
1!
1%
#621270000000
0!
0%
#621275000000
1!
1%
#621280000000
0!
0%
#621285000000
1!
1%
#621290000000
0!
0%
#621295000000
1!
1%
#621300000000
0!
0%
#621305000000
1!
1%
#621310000000
0!
0%
#621315000000
1!
1%
#621320000000
0!
0%
#621325000000
1!
1%
#621330000000
0!
0%
#621335000000
1!
1%
#621340000000
0!
0%
#621345000000
1!
1%
#621350000000
0!
0%
#621355000000
1!
1%
#621360000000
0!
0%
#621365000000
1!
1%
#621370000000
0!
0%
#621375000000
1!
1%
#621380000000
0!
0%
#621385000000
1!
1%
#621390000000
0!
0%
#621395000000
1!
1%
#621400000000
0!
0%
#621405000000
1!
1%
#621410000000
0!
0%
#621415000000
1!
1%
#621420000000
0!
0%
#621425000000
1!
1%
#621430000000
0!
0%
#621435000000
1!
1%
#621440000000
0!
0%
#621445000000
1!
1%
#621450000000
0!
0%
#621455000000
1!
1%
#621460000000
0!
0%
#621465000000
1!
1%
#621470000000
0!
0%
#621475000000
1!
1%
#621480000000
0!
0%
#621485000000
1!
1%
#621490000000
0!
0%
#621495000000
1!
1%
#621500000000
0!
0%
#621505000000
1!
1%
#621510000000
0!
0%
#621515000000
1!
1%
#621520000000
0!
0%
#621525000000
1!
1%
#621530000000
0!
0%
#621535000000
1!
1%
#621540000000
0!
0%
#621545000000
1!
1%
#621550000000
0!
0%
#621555000000
1!
1%
#621560000000
0!
0%
#621565000000
1!
1%
#621570000000
0!
0%
#621575000000
1!
1%
#621580000000
0!
0%
#621585000000
1!
1%
#621590000000
0!
0%
#621595000000
1!
1%
#621600000000
0!
0%
#621605000000
1!
1%
#621610000000
0!
0%
#621615000000
1!
1%
#621620000000
0!
0%
#621625000000
1!
1%
#621630000000
0!
0%
#621635000000
1!
1%
#621640000000
0!
0%
#621645000000
1!
1%
#621650000000
0!
0%
#621655000000
1!
1%
#621660000000
0!
0%
#621665000000
1!
1%
#621670000000
0!
0%
#621675000000
1!
1%
#621680000000
0!
0%
#621685000000
1!
1%
#621690000000
0!
0%
#621695000000
1!
1%
#621700000000
0!
0%
#621705000000
1!
1%
#621710000000
0!
0%
#621715000000
1!
1%
#621720000000
0!
0%
#621725000000
1!
1%
#621730000000
0!
0%
#621735000000
1!
1%
#621740000000
0!
0%
#621745000000
1!
1%
#621750000000
0!
0%
#621755000000
1!
1%
#621760000000
0!
0%
#621765000000
1!
1%
#621770000000
0!
0%
#621775000000
1!
1%
#621780000000
0!
0%
#621785000000
1!
1%
#621790000000
0!
0%
#621795000000
1!
1%
#621800000000
0!
0%
#621805000000
1!
1%
#621810000000
0!
0%
#621815000000
1!
1%
#621820000000
0!
0%
#621825000000
1!
1%
#621830000000
0!
0%
#621835000000
1!
1%
#621840000000
0!
0%
#621845000000
1!
1%
#621850000000
0!
0%
#621855000000
1!
1%
#621860000000
0!
0%
#621865000000
1!
1%
#621870000000
0!
0%
#621875000000
1!
1%
#621880000000
0!
0%
#621885000000
1!
1%
#621890000000
0!
0%
#621895000000
1!
1%
#621900000000
0!
0%
#621905000000
1!
1%
#621910000000
0!
0%
#621915000000
1!
1%
#621920000000
0!
0%
#621925000000
1!
1%
#621930000000
0!
0%
#621935000000
1!
1%
#621940000000
0!
0%
#621945000000
1!
1%
#621950000000
0!
0%
#621955000000
1!
1%
#621960000000
0!
0%
#621965000000
1!
1%
#621970000000
0!
0%
#621975000000
1!
1%
#621980000000
0!
0%
#621985000000
1!
1%
#621990000000
0!
0%
#621995000000
1!
1%
#622000000000
0!
0%
#622005000000
1!
1%
#622010000000
0!
0%
#622015000000
1!
1%
#622020000000
0!
0%
#622025000000
1!
1%
#622030000000
0!
0%
#622035000000
1!
1%
#622040000000
0!
0%
#622045000000
1!
1%
#622050000000
0!
0%
#622055000000
1!
1%
#622060000000
0!
0%
#622065000000
1!
1%
#622070000000
0!
0%
#622075000000
1!
1%
#622080000000
0!
0%
#622085000000
1!
1%
#622090000000
0!
0%
#622095000000
1!
1%
#622100000000
0!
0%
#622105000000
1!
1%
#622110000000
0!
0%
#622115000000
1!
1%
#622120000000
0!
0%
#622125000000
1!
1%
#622130000000
0!
0%
#622135000000
1!
1%
#622140000000
0!
0%
#622145000000
1!
1%
#622150000000
0!
0%
#622155000000
1!
1%
#622160000000
0!
0%
#622165000000
1!
1%
#622170000000
0!
0%
#622175000000
1!
1%
#622180000000
0!
0%
#622185000000
1!
1%
#622190000000
0!
0%
#622195000000
1!
1%
#622200000000
0!
0%
#622205000000
1!
1%
#622210000000
0!
0%
#622215000000
1!
1%
#622220000000
0!
0%
#622225000000
1!
1%
#622230000000
0!
0%
#622235000000
1!
1%
#622240000000
0!
0%
#622245000000
1!
1%
#622250000000
0!
0%
#622255000000
1!
1%
#622260000000
0!
0%
#622265000000
1!
1%
#622270000000
0!
0%
#622275000000
1!
1%
#622280000000
0!
0%
#622285000000
1!
1%
#622290000000
0!
0%
#622295000000
1!
1%
#622300000000
0!
0%
#622305000000
1!
1%
#622310000000
0!
0%
#622315000000
1!
1%
#622320000000
0!
0%
#622325000000
1!
1%
#622330000000
0!
0%
#622335000000
1!
1%
#622340000000
0!
0%
#622345000000
1!
1%
#622350000000
0!
0%
#622355000000
1!
1%
#622360000000
0!
0%
#622365000000
1!
1%
#622370000000
0!
0%
#622375000000
1!
1%
#622380000000
0!
0%
#622385000000
1!
1%
#622390000000
0!
0%
#622395000000
1!
1%
#622400000000
0!
0%
#622405000000
1!
1%
#622410000000
0!
0%
#622415000000
1!
1%
#622420000000
0!
0%
#622425000000
1!
1%
#622430000000
0!
0%
#622435000000
1!
1%
#622440000000
0!
0%
#622445000000
1!
1%
#622450000000
0!
0%
#622455000000
1!
1%
#622460000000
0!
0%
#622465000000
1!
1%
#622470000000
0!
0%
#622475000000
1!
1%
#622480000000
0!
0%
#622485000000
1!
1%
#622490000000
0!
0%
#622495000000
1!
1%
#622500000000
0!
0%
#622505000000
1!
1%
#622510000000
0!
0%
#622515000000
1!
1%
#622520000000
0!
0%
#622525000000
1!
1%
#622530000000
0!
0%
#622535000000
1!
1%
#622540000000
0!
0%
#622545000000
1!
1%
#622550000000
0!
0%
#622555000000
1!
1%
#622560000000
0!
0%
#622565000000
1!
1%
#622570000000
0!
0%
#622575000000
1!
1%
#622580000000
0!
0%
#622585000000
1!
1%
#622590000000
0!
0%
#622595000000
1!
1%
#622600000000
0!
0%
#622605000000
1!
1%
#622610000000
0!
0%
#622615000000
1!
1%
#622620000000
0!
0%
#622625000000
1!
1%
#622630000000
0!
0%
#622635000000
1!
1%
#622640000000
0!
0%
#622645000000
1!
1%
#622650000000
0!
0%
#622655000000
1!
1%
#622660000000
0!
0%
#622665000000
1!
1%
#622670000000
0!
0%
#622675000000
1!
1%
#622680000000
0!
0%
#622685000000
1!
1%
#622690000000
0!
0%
#622695000000
1!
1%
#622700000000
0!
0%
#622705000000
1!
1%
#622710000000
0!
0%
#622715000000
1!
1%
#622720000000
0!
0%
#622725000000
1!
1%
#622730000000
0!
0%
#622735000000
1!
1%
#622740000000
0!
0%
#622745000000
1!
1%
#622750000000
0!
0%
#622755000000
1!
1%
#622760000000
0!
0%
#622765000000
1!
1%
#622770000000
0!
0%
#622775000000
1!
1%
#622780000000
0!
0%
#622785000000
1!
1%
#622790000000
0!
0%
#622795000000
1!
1%
#622800000000
0!
0%
#622805000000
1!
1%
#622810000000
0!
0%
#622815000000
1!
1%
#622820000000
0!
0%
#622825000000
1!
1%
#622830000000
0!
0%
#622835000000
1!
1%
#622840000000
0!
0%
#622845000000
1!
1%
#622850000000
0!
0%
#622855000000
1!
1%
#622860000000
0!
0%
#622865000000
1!
1%
#622870000000
0!
0%
#622875000000
1!
1%
#622880000000
0!
0%
#622885000000
1!
1%
#622890000000
0!
0%
#622895000000
1!
1%
#622900000000
0!
0%
#622905000000
1!
1%
#622910000000
0!
0%
#622915000000
1!
1%
#622920000000
0!
0%
#622925000000
1!
1%
#622930000000
0!
0%
#622935000000
1!
1%
#622940000000
0!
0%
#622945000000
1!
1%
#622950000000
0!
0%
#622955000000
1!
1%
#622960000000
0!
0%
#622965000000
1!
1%
#622970000000
0!
0%
#622975000000
1!
1%
#622980000000
0!
0%
#622985000000
1!
1%
#622990000000
0!
0%
#622995000000
1!
1%
#623000000000
0!
0%
#623005000000
1!
1%
#623010000000
0!
0%
#623015000000
1!
1%
#623020000000
0!
0%
#623025000000
1!
1%
#623030000000
0!
0%
#623035000000
1!
1%
#623040000000
0!
0%
#623045000000
1!
1%
#623050000000
0!
0%
#623055000000
1!
1%
#623060000000
0!
0%
#623065000000
1!
1%
#623070000000
0!
0%
#623075000000
1!
1%
#623080000000
0!
0%
#623085000000
1!
1%
#623090000000
0!
0%
#623095000000
1!
1%
#623100000000
0!
0%
#623105000000
1!
1%
#623110000000
0!
0%
#623115000000
1!
1%
#623120000000
0!
0%
#623125000000
1!
1%
#623130000000
0!
0%
#623135000000
1!
1%
#623140000000
0!
0%
#623145000000
1!
1%
#623150000000
0!
0%
#623155000000
1!
1%
#623160000000
0!
0%
#623165000000
1!
1%
#623170000000
0!
0%
#623175000000
1!
1%
#623180000000
0!
0%
#623185000000
1!
1%
#623190000000
0!
0%
#623195000000
1!
1%
#623200000000
0!
0%
#623205000000
1!
1%
#623210000000
0!
0%
#623215000000
1!
1%
#623220000000
0!
0%
#623225000000
1!
1%
#623230000000
0!
0%
#623235000000
1!
1%
#623240000000
0!
0%
#623245000000
1!
1%
#623250000000
0!
0%
#623255000000
1!
1%
#623260000000
0!
0%
#623265000000
1!
1%
#623270000000
0!
0%
#623275000000
1!
1%
#623280000000
0!
0%
#623285000000
1!
1%
#623290000000
0!
0%
#623295000000
1!
1%
#623300000000
0!
0%
#623305000000
1!
1%
#623310000000
0!
0%
#623315000000
1!
1%
#623320000000
0!
0%
#623325000000
1!
1%
#623330000000
0!
0%
#623335000000
1!
1%
#623340000000
0!
0%
#623345000000
1!
1%
#623350000000
0!
0%
#623355000000
1!
1%
#623360000000
0!
0%
#623365000000
1!
1%
#623370000000
0!
0%
#623375000000
1!
1%
#623380000000
0!
0%
#623385000000
1!
1%
#623390000000
0!
0%
#623395000000
1!
1%
#623400000000
0!
0%
#623405000000
1!
1%
#623410000000
0!
0%
#623415000000
1!
1%
#623420000000
0!
0%
#623425000000
1!
1%
#623430000000
0!
0%
#623435000000
1!
1%
#623440000000
0!
0%
#623445000000
1!
1%
#623450000000
0!
0%
#623455000000
1!
1%
#623460000000
0!
0%
#623465000000
1!
1%
#623470000000
0!
0%
#623475000000
1!
1%
#623480000000
0!
0%
#623485000000
1!
1%
#623490000000
0!
0%
#623495000000
1!
1%
#623500000000
0!
0%
#623505000000
1!
1%
#623510000000
0!
0%
#623515000000
1!
1%
#623520000000
0!
0%
#623525000000
1!
1%
#623530000000
0!
0%
#623535000000
1!
1%
#623540000000
0!
0%
#623545000000
1!
1%
#623550000000
0!
0%
#623555000000
1!
1%
#623560000000
0!
0%
#623565000000
1!
1%
#623570000000
0!
0%
#623575000000
1!
1%
#623580000000
0!
0%
#623585000000
1!
1%
#623590000000
0!
0%
#623595000000
1!
1%
#623600000000
0!
0%
#623605000000
1!
1%
#623610000000
0!
0%
#623615000000
1!
1%
#623620000000
0!
0%
#623625000000
1!
1%
#623630000000
0!
0%
#623635000000
1!
1%
#623640000000
0!
0%
#623645000000
1!
1%
#623650000000
0!
0%
#623655000000
1!
1%
#623660000000
0!
0%
#623665000000
1!
1%
#623670000000
0!
0%
#623675000000
1!
1%
#623680000000
0!
0%
#623685000000
1!
1%
#623690000000
0!
0%
#623695000000
1!
1%
#623700000000
0!
0%
#623705000000
1!
1%
#623710000000
0!
0%
#623715000000
1!
1%
#623720000000
0!
0%
#623725000000
1!
1%
#623730000000
0!
0%
#623735000000
1!
1%
#623740000000
0!
0%
#623745000000
1!
1%
#623750000000
0!
0%
#623755000000
1!
1%
#623760000000
0!
0%
#623765000000
1!
1%
#623770000000
0!
0%
#623775000000
1!
1%
#623780000000
0!
0%
#623785000000
1!
1%
#623790000000
0!
0%
#623795000000
1!
1%
#623800000000
0!
0%
#623805000000
1!
1%
#623810000000
0!
0%
#623815000000
1!
1%
#623820000000
0!
0%
#623825000000
1!
1%
#623830000000
0!
0%
#623835000000
1!
1%
#623840000000
0!
0%
#623845000000
1!
1%
#623850000000
0!
0%
#623855000000
1!
1%
#623860000000
0!
0%
#623865000000
1!
1%
#623870000000
0!
0%
#623875000000
1!
1%
#623880000000
0!
0%
#623885000000
1!
1%
#623890000000
0!
0%
#623895000000
1!
1%
#623900000000
0!
0%
#623905000000
1!
1%
#623910000000
0!
0%
#623915000000
1!
1%
#623920000000
0!
0%
#623925000000
1!
1%
#623930000000
0!
0%
#623935000000
1!
1%
#623940000000
0!
0%
#623945000000
1!
1%
#623950000000
0!
0%
#623955000000
1!
1%
#623960000000
0!
0%
#623965000000
1!
1%
#623970000000
0!
0%
#623975000000
1!
1%
#623980000000
0!
0%
#623985000000
1!
1%
#623990000000
0!
0%
#623995000000
1!
1%
#624000000000
0!
0%
#624005000000
1!
1%
#624010000000
0!
0%
#624015000000
1!
1%
#624020000000
0!
0%
#624025000000
1!
1%
#624030000000
0!
0%
#624035000000
1!
1%
#624040000000
0!
0%
#624045000000
1!
1%
#624050000000
0!
0%
#624055000000
1!
1%
#624060000000
0!
0%
#624065000000
1!
1%
#624070000000
0!
0%
#624075000000
1!
1%
#624080000000
0!
0%
#624085000000
1!
1%
#624090000000
0!
0%
#624095000000
1!
1%
#624100000000
0!
0%
#624105000000
1!
1%
#624110000000
0!
0%
#624115000000
1!
1%
#624120000000
0!
0%
#624125000000
1!
1%
#624130000000
0!
0%
#624135000000
1!
1%
#624140000000
0!
0%
#624145000000
1!
1%
#624150000000
0!
0%
#624155000000
1!
1%
#624160000000
0!
0%
#624165000000
1!
1%
#624170000000
0!
0%
#624175000000
1!
1%
#624180000000
0!
0%
#624185000000
1!
1%
#624190000000
0!
0%
#624195000000
1!
1%
#624200000000
0!
0%
#624205000000
1!
1%
#624210000000
0!
0%
#624215000000
1!
1%
#624220000000
0!
0%
#624225000000
1!
1%
#624230000000
0!
0%
#624235000000
1!
1%
#624240000000
0!
0%
#624245000000
1!
1%
#624250000000
0!
0%
#624255000000
1!
1%
#624260000000
0!
0%
#624265000000
1!
1%
#624270000000
0!
0%
#624275000000
1!
1%
#624280000000
0!
0%
#624285000000
1!
1%
#624290000000
0!
0%
#624295000000
1!
1%
#624300000000
0!
0%
#624305000000
1!
1%
#624310000000
0!
0%
#624315000000
1!
1%
#624320000000
0!
0%
#624325000000
1!
1%
#624330000000
0!
0%
#624335000000
1!
1%
#624340000000
0!
0%
#624345000000
1!
1%
#624350000000
0!
0%
#624355000000
1!
1%
#624360000000
0!
0%
#624365000000
1!
1%
#624370000000
0!
0%
#624375000000
1!
1%
#624380000000
0!
0%
#624385000000
1!
1%
#624390000000
0!
0%
#624395000000
1!
1%
#624400000000
0!
0%
#624405000000
1!
1%
#624410000000
0!
0%
#624415000000
1!
1%
#624420000000
0!
0%
#624425000000
1!
1%
#624430000000
0!
0%
#624435000000
1!
1%
#624440000000
0!
0%
#624445000000
1!
1%
#624450000000
0!
0%
#624455000000
1!
1%
#624460000000
0!
0%
#624465000000
1!
1%
#624470000000
0!
0%
#624475000000
1!
1%
#624480000000
0!
0%
#624485000000
1!
1%
#624490000000
0!
0%
#624495000000
1!
1%
#624500000000
0!
0%
#624505000000
1!
1%
#624510000000
0!
0%
#624515000000
1!
1%
#624520000000
0!
0%
#624525000000
1!
1%
#624530000000
0!
0%
#624535000000
1!
1%
#624540000000
0!
0%
#624545000000
1!
1%
#624550000000
0!
0%
#624555000000
1!
1%
#624560000000
0!
0%
#624565000000
1!
1%
#624570000000
0!
0%
#624575000000
1!
1%
#624580000000
0!
0%
#624585000000
1!
1%
#624590000000
0!
0%
#624595000000
1!
1%
#624600000000
0!
0%
#624605000000
1!
1%
#624610000000
0!
0%
#624615000000
1!
1%
#624620000000
0!
0%
#624625000000
1!
1%
#624630000000
0!
0%
#624635000000
1!
1%
#624640000000
0!
0%
#624645000000
1!
1%
#624650000000
0!
0%
#624655000000
1!
1%
#624660000000
0!
0%
#624665000000
1!
1%
#624670000000
0!
0%
#624675000000
1!
1%
#624680000000
0!
0%
#624685000000
1!
1%
#624690000000
0!
0%
#624695000000
1!
1%
#624700000000
0!
0%
#624705000000
1!
1%
#624710000000
0!
0%
#624715000000
1!
1%
#624720000000
0!
0%
#624725000000
1!
1%
#624730000000
0!
0%
#624735000000
1!
1%
#624740000000
0!
0%
#624745000000
1!
1%
#624750000000
0!
0%
#624755000000
1!
1%
#624760000000
0!
0%
#624765000000
1!
1%
#624770000000
0!
0%
#624775000000
1!
1%
#624780000000
0!
0%
#624785000000
1!
1%
#624790000000
0!
0%
#624795000000
1!
1%
#624800000000
0!
0%
#624805000000
1!
1%
#624810000000
0!
0%
#624815000000
1!
1%
#624820000000
0!
0%
#624825000000
1!
1%
#624830000000
0!
0%
#624835000000
1!
1%
#624840000000
0!
0%
#624845000000
1!
1%
#624850000000
0!
0%
#624855000000
1!
1%
#624860000000
0!
0%
#624865000000
1!
1%
#624870000000
0!
0%
#624875000000
1!
1%
#624880000000
0!
0%
#624885000000
1!
1%
#624890000000
0!
0%
#624895000000
1!
1%
#624900000000
0!
0%
#624905000000
1!
1%
#624910000000
0!
0%
#624915000000
1!
1%
#624920000000
0!
0%
#624925000000
1!
1%
#624930000000
0!
0%
#624935000000
1!
1%
#624940000000
0!
0%
#624945000000
1!
1%
#624950000000
0!
0%
#624955000000
1!
1%
#624960000000
0!
0%
#624965000000
1!
1%
#624970000000
0!
0%
#624975000000
1!
1%
#624980000000
0!
0%
#624985000000
1!
1%
#624990000000
0!
0%
#624995000000
1!
1%
#625000000000
0!
0%
#625005000000
1!
1%
#625010000000
0!
0%
#625015000000
1!
1%
#625020000000
0!
0%
#625025000000
1!
1%
#625030000000
0!
0%
#625035000000
1!
1%
#625040000000
0!
0%
#625045000000
1!
1%
#625050000000
0!
0%
#625055000000
1!
1%
#625060000000
0!
0%
#625065000000
1!
1%
#625070000000
0!
0%
#625075000000
1!
1%
#625080000000
0!
0%
#625085000000
1!
1%
#625090000000
0!
0%
#625095000000
1!
1%
#625100000000
0!
0%
#625105000000
1!
1%
#625110000000
0!
0%
#625115000000
1!
1%
#625120000000
0!
0%
#625125000000
1!
1%
#625130000000
0!
0%
#625135000000
1!
1%
#625140000000
0!
0%
#625145000000
1!
1%
#625150000000
0!
0%
#625155000000
1!
1%
#625160000000
0!
0%
#625165000000
1!
1%
#625170000000
0!
0%
#625175000000
1!
1%
#625180000000
0!
0%
#625185000000
1!
1%
#625190000000
0!
0%
#625195000000
1!
1%
#625200000000
0!
0%
#625205000000
1!
1%
#625210000000
0!
0%
#625215000000
1!
1%
#625220000000
0!
0%
#625225000000
1!
1%
#625230000000
0!
0%
#625235000000
1!
1%
#625240000000
0!
0%
#625245000000
1!
1%
#625250000000
0!
0%
#625255000000
1!
1%
#625260000000
0!
0%
#625265000000
1!
1%
#625270000000
0!
0%
#625275000000
1!
1%
#625280000000
0!
0%
#625285000000
1!
1%
#625290000000
0!
0%
#625295000000
1!
1%
#625300000000
0!
0%
#625305000000
1!
1%
#625310000000
0!
0%
#625315000000
1!
1%
#625320000000
0!
0%
#625325000000
1!
1%
#625330000000
0!
0%
#625335000000
1!
1%
#625340000000
0!
0%
#625345000000
1!
1%
#625350000000
0!
0%
#625355000000
1!
1%
#625360000000
0!
0%
#625365000000
1!
1%
#625370000000
0!
0%
#625375000000
1!
1%
#625380000000
0!
0%
#625385000000
1!
1%
#625390000000
0!
0%
#625395000000
1!
1%
#625400000000
0!
0%
#625405000000
1!
1%
#625410000000
0!
0%
#625415000000
1!
1%
#625420000000
0!
0%
#625425000000
1!
1%
#625430000000
0!
0%
#625435000000
1!
1%
#625440000000
0!
0%
#625445000000
1!
1%
#625450000000
0!
0%
#625455000000
1!
1%
#625460000000
0!
0%
#625465000000
1!
1%
#625470000000
0!
0%
#625475000000
1!
1%
#625480000000
0!
0%
#625485000000
1!
1%
#625490000000
0!
0%
#625495000000
1!
1%
#625500000000
0!
0%
#625505000000
1!
1%
#625510000000
0!
0%
#625515000000
1!
1%
#625520000000
0!
0%
#625525000000
1!
1%
#625530000000
0!
0%
#625535000000
1!
1%
#625540000000
0!
0%
#625545000000
1!
1%
#625550000000
0!
0%
#625555000000
1!
1%
#625560000000
0!
0%
#625565000000
1!
1%
#625570000000
0!
0%
#625575000000
1!
1%
#625580000000
0!
0%
#625585000000
1!
1%
#625590000000
0!
0%
#625595000000
1!
1%
#625600000000
0!
0%
#625605000000
1!
1%
#625610000000
0!
0%
#625615000000
1!
1%
#625620000000
0!
0%
#625625000000
1!
1%
#625630000000
0!
0%
#625635000000
1!
1%
#625640000000
0!
0%
#625645000000
1!
1%
#625650000000
0!
0%
#625655000000
1!
1%
#625660000000
0!
0%
#625665000000
1!
1%
#625670000000
0!
0%
#625675000000
1!
1%
#625680000000
0!
0%
#625685000000
1!
1%
#625690000000
0!
0%
#625695000000
1!
1%
#625700000000
0!
0%
#625705000000
1!
1%
#625710000000
0!
0%
#625715000000
1!
1%
#625720000000
0!
0%
#625725000000
1!
1%
#625730000000
0!
0%
#625735000000
1!
1%
#625740000000
0!
0%
#625745000000
1!
1%
#625750000000
0!
0%
#625755000000
1!
1%
#625760000000
0!
0%
#625765000000
1!
1%
#625770000000
0!
0%
#625775000000
1!
1%
#625780000000
0!
0%
#625785000000
1!
1%
#625790000000
0!
0%
#625795000000
1!
1%
#625800000000
0!
0%
#625805000000
1!
1%
#625810000000
0!
0%
#625815000000
1!
1%
#625820000000
0!
0%
#625825000000
1!
1%
#625830000000
0!
0%
#625835000000
1!
1%
#625840000000
0!
0%
#625845000000
1!
1%
#625850000000
0!
0%
#625855000000
1!
1%
#625860000000
0!
0%
#625865000000
1!
1%
#625870000000
0!
0%
#625875000000
1!
1%
#625880000000
0!
0%
#625885000000
1!
1%
#625890000000
0!
0%
#625895000000
1!
1%
#625900000000
0!
0%
#625905000000
1!
1%
#625910000000
0!
0%
#625915000000
1!
1%
#625920000000
0!
0%
#625925000000
1!
1%
#625930000000
0!
0%
#625935000000
1!
1%
#625940000000
0!
0%
#625945000000
1!
1%
#625950000000
0!
0%
#625955000000
1!
1%
#625960000000
0!
0%
#625965000000
1!
1%
#625970000000
0!
0%
#625975000000
1!
1%
#625980000000
0!
0%
#625985000000
1!
1%
#625990000000
0!
0%
#625995000000
1!
1%
#626000000000
0!
0%
#626005000000
1!
1%
#626010000000
0!
0%
#626015000000
1!
1%
#626020000000
0!
0%
#626025000000
1!
1%
#626030000000
0!
0%
#626035000000
1!
1%
#626040000000
0!
0%
#626045000000
1!
1%
#626050000000
0!
0%
#626055000000
1!
1%
#626060000000
0!
0%
#626065000000
1!
1%
#626070000000
0!
0%
#626075000000
1!
1%
#626080000000
0!
0%
#626085000000
1!
1%
#626090000000
0!
0%
#626095000000
1!
1%
#626100000000
0!
0%
#626105000000
1!
1%
#626110000000
0!
0%
#626115000000
1!
1%
#626120000000
0!
0%
#626125000000
1!
1%
#626130000000
0!
0%
#626135000000
1!
1%
#626140000000
0!
0%
#626145000000
1!
1%
#626150000000
0!
0%
#626155000000
1!
1%
#626160000000
0!
0%
#626165000000
1!
1%
#626170000000
0!
0%
#626175000000
1!
1%
#626180000000
0!
0%
#626185000000
1!
1%
#626190000000
0!
0%
#626195000000
1!
1%
#626200000000
0!
0%
#626205000000
1!
1%
#626210000000
0!
0%
#626215000000
1!
1%
#626220000000
0!
0%
#626225000000
1!
1%
#626230000000
0!
0%
#626235000000
1!
1%
#626240000000
0!
0%
#626245000000
1!
1%
#626250000000
0!
0%
#626255000000
1!
1%
#626260000000
0!
0%
#626265000000
1!
1%
#626270000000
0!
0%
#626275000000
1!
1%
#626280000000
0!
0%
#626285000000
1!
1%
#626290000000
0!
0%
#626295000000
1!
1%
#626300000000
0!
0%
#626305000000
1!
1%
#626310000000
0!
0%
#626315000000
1!
1%
#626320000000
0!
0%
#626325000000
1!
1%
#626330000000
0!
0%
#626335000000
1!
1%
#626340000000
0!
0%
#626345000000
1!
1%
#626350000000
0!
0%
#626355000000
1!
1%
#626360000000
0!
0%
#626365000000
1!
1%
#626370000000
0!
0%
#626375000000
1!
1%
#626380000000
0!
0%
#626385000000
1!
1%
#626390000000
0!
0%
#626395000000
1!
1%
#626400000000
0!
0%
#626405000000
1!
1%
#626410000000
0!
0%
#626415000000
1!
1%
#626420000000
0!
0%
#626425000000
1!
1%
#626430000000
0!
0%
#626435000000
1!
1%
#626440000000
0!
0%
#626445000000
1!
1%
#626450000000
0!
0%
#626455000000
1!
1%
#626460000000
0!
0%
#626465000000
1!
1%
#626470000000
0!
0%
#626475000000
1!
1%
#626480000000
0!
0%
#626485000000
1!
1%
#626490000000
0!
0%
#626495000000
1!
1%
#626500000000
0!
0%
#626505000000
1!
1%
#626510000000
0!
0%
#626515000000
1!
1%
#626520000000
0!
0%
#626525000000
1!
1%
#626530000000
0!
0%
#626535000000
1!
1%
#626540000000
0!
0%
#626545000000
1!
1%
#626550000000
0!
0%
#626555000000
1!
1%
#626560000000
0!
0%
#626565000000
1!
1%
#626570000000
0!
0%
#626575000000
1!
1%
#626580000000
0!
0%
#626585000000
1!
1%
#626590000000
0!
0%
#626595000000
1!
1%
#626600000000
0!
0%
#626605000000
1!
1%
#626610000000
0!
0%
#626615000000
1!
1%
#626620000000
0!
0%
#626625000000
1!
1%
#626630000000
0!
0%
#626635000000
1!
1%
#626640000000
0!
0%
#626645000000
1!
1%
#626650000000
0!
0%
#626655000000
1!
1%
#626660000000
0!
0%
#626665000000
1!
1%
#626670000000
0!
0%
#626675000000
1!
1%
#626680000000
0!
0%
#626685000000
1!
1%
#626690000000
0!
0%
#626695000000
1!
1%
#626700000000
0!
0%
#626705000000
1!
1%
#626710000000
0!
0%
#626715000000
1!
1%
#626720000000
0!
0%
#626725000000
1!
1%
#626730000000
0!
0%
#626735000000
1!
1%
#626740000000
0!
0%
#626745000000
1!
1%
#626750000000
0!
0%
#626755000000
1!
1%
#626760000000
0!
0%
#626765000000
1!
1%
#626770000000
0!
0%
#626775000000
1!
1%
#626780000000
0!
0%
#626785000000
1!
1%
#626790000000
0!
0%
#626795000000
1!
1%
#626800000000
0!
0%
#626805000000
1!
1%
#626810000000
0!
0%
#626815000000
1!
1%
#626820000000
0!
0%
#626825000000
1!
1%
#626830000000
0!
0%
#626835000000
1!
1%
#626840000000
0!
0%
#626845000000
1!
1%
#626850000000
0!
0%
#626855000000
1!
1%
#626860000000
0!
0%
#626865000000
1!
1%
#626870000000
0!
0%
#626875000000
1!
1%
#626880000000
0!
0%
#626885000000
1!
1%
#626890000000
0!
0%
#626895000000
1!
1%
#626900000000
0!
0%
#626905000000
1!
1%
#626910000000
0!
0%
#626915000000
1!
1%
#626920000000
0!
0%
#626925000000
1!
1%
#626930000000
0!
0%
#626935000000
1!
1%
#626940000000
0!
0%
#626945000000
1!
1%
#626950000000
0!
0%
#626955000000
1!
1%
#626960000000
0!
0%
#626965000000
1!
1%
#626970000000
0!
0%
#626975000000
1!
1%
#626980000000
0!
0%
#626985000000
1!
1%
#626990000000
0!
0%
#626995000000
1!
1%
#627000000000
0!
0%
#627005000000
1!
1%
#627010000000
0!
0%
#627015000000
1!
1%
#627020000000
0!
0%
#627025000000
1!
1%
#627030000000
0!
0%
#627035000000
1!
1%
#627040000000
0!
0%
#627045000000
1!
1%
#627050000000
0!
0%
#627055000000
1!
1%
#627060000000
0!
0%
#627065000000
1!
1%
#627070000000
0!
0%
#627075000000
1!
1%
#627080000000
0!
0%
#627085000000
1!
1%
#627090000000
0!
0%
#627095000000
1!
1%
#627100000000
0!
0%
#627105000000
1!
1%
#627110000000
0!
0%
#627115000000
1!
1%
#627120000000
0!
0%
#627125000000
1!
1%
#627130000000
0!
0%
#627135000000
1!
1%
#627140000000
0!
0%
#627145000000
1!
1%
#627150000000
0!
0%
#627155000000
1!
1%
#627160000000
0!
0%
#627165000000
1!
1%
#627170000000
0!
0%
#627175000000
1!
1%
#627180000000
0!
0%
#627185000000
1!
1%
#627190000000
0!
0%
#627195000000
1!
1%
#627200000000
0!
0%
#627205000000
1!
1%
#627210000000
0!
0%
#627215000000
1!
1%
#627220000000
0!
0%
#627225000000
1!
1%
#627230000000
0!
0%
#627235000000
1!
1%
#627240000000
0!
0%
#627245000000
1!
1%
#627250000000
0!
0%
#627255000000
1!
1%
#627260000000
0!
0%
#627265000000
1!
1%
#627270000000
0!
0%
#627275000000
1!
1%
#627280000000
0!
0%
#627285000000
1!
1%
#627290000000
0!
0%
#627295000000
1!
1%
#627300000000
0!
0%
#627305000000
1!
1%
#627310000000
0!
0%
#627315000000
1!
1%
#627320000000
0!
0%
#627325000000
1!
1%
#627330000000
0!
0%
#627335000000
1!
1%
#627340000000
0!
0%
#627345000000
1!
1%
#627350000000
0!
0%
#627355000000
1!
1%
#627360000000
0!
0%
#627365000000
1!
1%
#627370000000
0!
0%
#627375000000
1!
1%
#627380000000
0!
0%
#627385000000
1!
1%
#627390000000
0!
0%
#627395000000
1!
1%
#627400000000
0!
0%
#627405000000
1!
1%
#627410000000
0!
0%
#627415000000
1!
1%
#627420000000
0!
0%
#627425000000
1!
1%
#627430000000
0!
0%
#627435000000
1!
1%
#627440000000
0!
0%
#627445000000
1!
1%
#627450000000
0!
0%
#627455000000
1!
1%
#627460000000
0!
0%
#627465000000
1!
1%
#627470000000
0!
0%
#627475000000
1!
1%
#627480000000
0!
0%
#627485000000
1!
1%
#627490000000
0!
0%
#627495000000
1!
1%
#627500000000
0!
0%
#627505000000
1!
1%
#627510000000
0!
0%
#627515000000
1!
1%
#627520000000
0!
0%
#627525000000
1!
1%
#627530000000
0!
0%
#627535000000
1!
1%
#627540000000
0!
0%
#627545000000
1!
1%
#627550000000
0!
0%
#627555000000
1!
1%
#627560000000
0!
0%
#627565000000
1!
1%
#627570000000
0!
0%
#627575000000
1!
1%
#627580000000
0!
0%
#627585000000
1!
1%
#627590000000
0!
0%
#627595000000
1!
1%
#627600000000
0!
0%
#627605000000
1!
1%
#627610000000
0!
0%
#627615000000
1!
1%
#627620000000
0!
0%
#627625000000
1!
1%
#627630000000
0!
0%
#627635000000
1!
1%
#627640000000
0!
0%
#627645000000
1!
1%
#627650000000
0!
0%
#627655000000
1!
1%
#627660000000
0!
0%
#627665000000
1!
1%
#627670000000
0!
0%
#627675000000
1!
1%
#627680000000
0!
0%
#627685000000
1!
1%
#627690000000
0!
0%
#627695000000
1!
1%
#627700000000
0!
0%
#627705000000
1!
1%
#627710000000
0!
0%
#627715000000
1!
1%
#627720000000
0!
0%
#627725000000
1!
1%
#627730000000
0!
0%
#627735000000
1!
1%
#627740000000
0!
0%
#627745000000
1!
1%
#627750000000
0!
0%
#627755000000
1!
1%
#627760000000
0!
0%
#627765000000
1!
1%
#627770000000
0!
0%
#627775000000
1!
1%
#627780000000
0!
0%
#627785000000
1!
1%
#627790000000
0!
0%
#627795000000
1!
1%
#627800000000
0!
0%
#627805000000
1!
1%
#627810000000
0!
0%
#627815000000
1!
1%
#627820000000
0!
0%
#627825000000
1!
1%
#627830000000
0!
0%
#627835000000
1!
1%
#627840000000
0!
0%
#627845000000
1!
1%
#627850000000
0!
0%
#627855000000
1!
1%
#627860000000
0!
0%
#627865000000
1!
1%
#627870000000
0!
0%
#627875000000
1!
1%
#627880000000
0!
0%
#627885000000
1!
1%
#627890000000
0!
0%
#627895000000
1!
1%
#627900000000
0!
0%
#627905000000
1!
1%
#627910000000
0!
0%
#627915000000
1!
1%
#627920000000
0!
0%
#627925000000
1!
1%
#627930000000
0!
0%
#627935000000
1!
1%
#627940000000
0!
0%
#627945000000
1!
1%
#627950000000
0!
0%
#627955000000
1!
1%
#627960000000
0!
0%
#627965000000
1!
1%
#627970000000
0!
0%
#627975000000
1!
1%
#627980000000
0!
0%
#627985000000
1!
1%
#627990000000
0!
0%
#627995000000
1!
1%
#628000000000
0!
0%
#628005000000
1!
1%
#628010000000
0!
0%
#628015000000
1!
1%
#628020000000
0!
0%
#628025000000
1!
1%
#628030000000
0!
0%
#628035000000
1!
1%
#628040000000
0!
0%
#628045000000
1!
1%
#628050000000
0!
0%
#628055000000
1!
1%
#628060000000
0!
0%
#628065000000
1!
1%
#628070000000
0!
0%
#628075000000
1!
1%
#628080000000
0!
0%
#628085000000
1!
1%
#628090000000
0!
0%
#628095000000
1!
1%
#628100000000
0!
0%
#628105000000
1!
1%
#628110000000
0!
0%
#628115000000
1!
1%
#628120000000
0!
0%
#628125000000
1!
1%
#628130000000
0!
0%
#628135000000
1!
1%
#628140000000
0!
0%
#628145000000
1!
1%
#628150000000
0!
0%
#628155000000
1!
1%
#628160000000
0!
0%
#628165000000
1!
1%
#628170000000
0!
0%
#628175000000
1!
1%
#628180000000
0!
0%
#628185000000
1!
1%
#628190000000
0!
0%
#628195000000
1!
1%
#628200000000
0!
0%
#628205000000
1!
1%
#628210000000
0!
0%
#628215000000
1!
1%
#628220000000
0!
0%
#628225000000
1!
1%
#628230000000
0!
0%
#628235000000
1!
1%
#628240000000
0!
0%
#628245000000
1!
1%
#628250000000
0!
0%
#628255000000
1!
1%
#628260000000
0!
0%
#628265000000
1!
1%
#628270000000
0!
0%
#628275000000
1!
1%
#628280000000
0!
0%
#628285000000
1!
1%
#628290000000
0!
0%
#628295000000
1!
1%
#628300000000
0!
0%
#628305000000
1!
1%
#628310000000
0!
0%
#628315000000
1!
1%
#628320000000
0!
0%
#628325000000
1!
1%
#628330000000
0!
0%
#628335000000
1!
1%
#628340000000
0!
0%
#628345000000
1!
1%
#628350000000
0!
0%
#628355000000
1!
1%
#628360000000
0!
0%
#628365000000
1!
1%
#628370000000
0!
0%
#628375000000
1!
1%
#628380000000
0!
0%
#628385000000
1!
1%
#628390000000
0!
0%
#628395000000
1!
1%
#628400000000
0!
0%
#628405000000
1!
1%
#628410000000
0!
0%
#628415000000
1!
1%
#628420000000
0!
0%
#628425000000
1!
1%
#628430000000
0!
0%
#628435000000
1!
1%
#628440000000
0!
0%
#628445000000
1!
1%
#628450000000
0!
0%
#628455000000
1!
1%
#628460000000
0!
0%
#628465000000
1!
1%
#628470000000
0!
0%
#628475000000
1!
1%
#628480000000
0!
0%
#628485000000
1!
1%
#628490000000
0!
0%
#628495000000
1!
1%
#628500000000
0!
0%
#628505000000
1!
1%
#628510000000
0!
0%
#628515000000
1!
1%
#628520000000
0!
0%
#628525000000
1!
1%
#628530000000
0!
0%
#628535000000
1!
1%
#628540000000
0!
0%
#628545000000
1!
1%
#628550000000
0!
0%
#628555000000
1!
1%
#628560000000
0!
0%
#628565000000
1!
1%
#628570000000
0!
0%
#628575000000
1!
1%
#628580000000
0!
0%
#628585000000
1!
1%
#628590000000
0!
0%
#628595000000
1!
1%
#628600000000
0!
0%
#628605000000
1!
1%
#628610000000
0!
0%
#628615000000
1!
1%
#628620000000
0!
0%
#628625000000
1!
1%
#628630000000
0!
0%
#628635000000
1!
1%
#628640000000
0!
0%
#628645000000
1!
1%
#628650000000
0!
0%
#628655000000
1!
1%
#628660000000
0!
0%
#628665000000
1!
1%
#628670000000
0!
0%
#628675000000
1!
1%
#628680000000
0!
0%
#628685000000
1!
1%
#628690000000
0!
0%
#628695000000
1!
1%
#628700000000
0!
0%
#628705000000
1!
1%
#628710000000
0!
0%
#628715000000
1!
1%
#628720000000
0!
0%
#628725000000
1!
1%
#628730000000
0!
0%
#628735000000
1!
1%
#628740000000
0!
0%
#628745000000
1!
1%
#628750000000
0!
0%
#628755000000
1!
1%
#628760000000
0!
0%
#628765000000
1!
1%
#628770000000
0!
0%
#628775000000
1!
1%
#628780000000
0!
0%
#628785000000
1!
1%
#628790000000
0!
0%
#628795000000
1!
1%
#628800000000
0!
0%
#628805000000
1!
1%
#628810000000
0!
0%
#628815000000
1!
1%
#628820000000
0!
0%
#628825000000
1!
1%
#628830000000
0!
0%
#628835000000
1!
1%
#628840000000
0!
0%
#628845000000
1!
1%
#628850000000
0!
0%
#628855000000
1!
1%
#628860000000
0!
0%
#628865000000
1!
1%
#628870000000
0!
0%
#628875000000
1!
1%
#628880000000
0!
0%
#628885000000
1!
1%
#628890000000
0!
0%
#628895000000
1!
1%
#628900000000
0!
0%
#628905000000
1!
1%
#628910000000
0!
0%
#628915000000
1!
1%
#628920000000
0!
0%
#628925000000
1!
1%
#628930000000
0!
0%
#628935000000
1!
1%
#628940000000
0!
0%
#628945000000
1!
1%
#628950000000
0!
0%
#628955000000
1!
1%
#628960000000
0!
0%
#628965000000
1!
1%
#628970000000
0!
0%
#628975000000
1!
1%
#628980000000
0!
0%
#628985000000
1!
1%
#628990000000
0!
0%
#628995000000
1!
1%
#629000000000
0!
0%
#629005000000
1!
1%
#629010000000
0!
0%
#629015000000
1!
1%
#629020000000
0!
0%
#629025000000
1!
1%
#629030000000
0!
0%
#629035000000
1!
1%
#629040000000
0!
0%
#629045000000
1!
1%
#629050000000
0!
0%
#629055000000
1!
1%
#629060000000
0!
0%
#629065000000
1!
1%
#629070000000
0!
0%
#629075000000
1!
1%
#629080000000
0!
0%
#629085000000
1!
1%
#629090000000
0!
0%
#629095000000
1!
1%
#629100000000
0!
0%
#629105000000
1!
1%
#629110000000
0!
0%
#629115000000
1!
1%
#629120000000
0!
0%
#629125000000
1!
1%
#629130000000
0!
0%
#629135000000
1!
1%
#629140000000
0!
0%
#629145000000
1!
1%
#629150000000
0!
0%
#629155000000
1!
1%
#629160000000
0!
0%
#629165000000
1!
1%
#629170000000
0!
0%
#629175000000
1!
1%
#629180000000
0!
0%
#629185000000
1!
1%
#629190000000
0!
0%
#629195000000
1!
1%
#629200000000
0!
0%
#629205000000
1!
1%
#629210000000
0!
0%
#629215000000
1!
1%
#629220000000
0!
0%
#629225000000
1!
1%
#629230000000
0!
0%
#629235000000
1!
1%
#629240000000
0!
0%
#629245000000
1!
1%
#629250000000
0!
0%
#629255000000
1!
1%
#629260000000
0!
0%
#629265000000
1!
1%
#629270000000
0!
0%
#629275000000
1!
1%
#629280000000
0!
0%
#629285000000
1!
1%
#629290000000
0!
0%
#629295000000
1!
1%
#629300000000
0!
0%
#629305000000
1!
1%
#629310000000
0!
0%
#629315000000
1!
1%
#629320000000
0!
0%
#629325000000
1!
1%
#629330000000
0!
0%
#629335000000
1!
1%
#629340000000
0!
0%
#629345000000
1!
1%
#629350000000
0!
0%
#629355000000
1!
1%
#629360000000
0!
0%
#629365000000
1!
1%
#629370000000
0!
0%
#629375000000
1!
1%
#629380000000
0!
0%
#629385000000
1!
1%
#629390000000
0!
0%
#629395000000
1!
1%
#629400000000
0!
0%
#629405000000
1!
1%
#629410000000
0!
0%
#629415000000
1!
1%
#629420000000
0!
0%
#629425000000
1!
1%
#629430000000
0!
0%
#629435000000
1!
1%
#629440000000
0!
0%
#629445000000
1!
1%
#629450000000
0!
0%
#629455000000
1!
1%
#629460000000
0!
0%
#629465000000
1!
1%
#629470000000
0!
0%
#629475000000
1!
1%
#629480000000
0!
0%
#629485000000
1!
1%
#629490000000
0!
0%
#629495000000
1!
1%
#629500000000
0!
0%
#629505000000
1!
1%
#629510000000
0!
0%
#629515000000
1!
1%
#629520000000
0!
0%
#629525000000
1!
1%
#629530000000
0!
0%
#629535000000
1!
1%
#629540000000
0!
0%
#629545000000
1!
1%
#629550000000
0!
0%
#629555000000
1!
1%
#629560000000
0!
0%
#629565000000
1!
1%
#629570000000
0!
0%
#629575000000
1!
1%
#629580000000
0!
0%
#629585000000
1!
1%
#629590000000
0!
0%
#629595000000
1!
1%
#629600000000
0!
0%
#629605000000
1!
1%
#629610000000
0!
0%
#629615000000
1!
1%
#629620000000
0!
0%
#629625000000
1!
1%
#629630000000
0!
0%
#629635000000
1!
1%
#629640000000
0!
0%
#629645000000
1!
1%
#629650000000
0!
0%
#629655000000
1!
1%
#629660000000
0!
0%
#629665000000
1!
1%
#629670000000
0!
0%
#629675000000
1!
1%
#629680000000
0!
0%
#629685000000
1!
1%
#629690000000
0!
0%
#629695000000
1!
1%
#629700000000
0!
0%
#629705000000
1!
1%
#629710000000
0!
0%
#629715000000
1!
1%
#629720000000
0!
0%
#629725000000
1!
1%
#629730000000
0!
0%
#629735000000
1!
1%
#629740000000
0!
0%
#629745000000
1!
1%
#629750000000
0!
0%
#629755000000
1!
1%
#629760000000
0!
0%
#629765000000
1!
1%
#629770000000
0!
0%
#629775000000
1!
1%
#629780000000
0!
0%
#629785000000
1!
1%
#629790000000
0!
0%
#629795000000
1!
1%
#629800000000
0!
0%
#629805000000
1!
1%
#629810000000
0!
0%
#629815000000
1!
1%
#629820000000
0!
0%
#629825000000
1!
1%
#629830000000
0!
0%
#629835000000
1!
1%
#629840000000
0!
0%
#629845000000
1!
1%
#629850000000
0!
0%
#629855000000
1!
1%
#629860000000
0!
0%
#629865000000
1!
1%
#629870000000
0!
0%
#629875000000
1!
1%
#629880000000
0!
0%
#629885000000
1!
1%
#629890000000
0!
0%
#629895000000
1!
1%
#629900000000
0!
0%
#629905000000
1!
1%
#629910000000
0!
0%
#629915000000
1!
1%
#629920000000
0!
0%
#629925000000
1!
1%
#629930000000
0!
0%
#629935000000
1!
1%
#629940000000
0!
0%
#629945000000
1!
1%
#629950000000
0!
0%
#629955000000
1!
1%
#629960000000
0!
0%
#629965000000
1!
1%
#629970000000
0!
0%
#629975000000
1!
1%
#629980000000
0!
0%
#629985000000
1!
1%
#629990000000
0!
0%
#629995000000
1!
1%
#630000000000
0!
0%
#630005000000
1!
1%
#630010000000
0!
0%
#630015000000
1!
1%
#630020000000
0!
0%
#630025000000
1!
1%
#630030000000
0!
0%
#630035000000
1!
1%
#630040000000
0!
0%
#630045000000
1!
1%
#630050000000
0!
0%
#630055000000
1!
1%
#630060000000
0!
0%
#630065000000
1!
1%
#630070000000
0!
0%
#630075000000
1!
1%
#630080000000
0!
0%
#630085000000
1!
1%
#630090000000
0!
0%
#630095000000
1!
1%
#630100000000
0!
0%
#630105000000
1!
1%
#630110000000
0!
0%
#630115000000
1!
1%
#630120000000
0!
0%
#630125000000
1!
1%
#630130000000
0!
0%
#630135000000
1!
1%
#630140000000
0!
0%
#630145000000
1!
1%
#630150000000
0!
0%
#630155000000
1!
1%
#630160000000
0!
0%
#630165000000
1!
1%
#630170000000
0!
0%
#630175000000
1!
1%
#630180000000
0!
0%
#630185000000
1!
1%
#630190000000
0!
0%
#630195000000
1!
1%
#630200000000
0!
0%
#630205000000
1!
1%
#630210000000
0!
0%
#630215000000
1!
1%
#630220000000
0!
0%
#630225000000
1!
1%
#630230000000
0!
0%
#630235000000
1!
1%
#630240000000
0!
0%
#630245000000
1!
1%
#630250000000
0!
0%
#630255000000
1!
1%
#630260000000
0!
0%
#630265000000
1!
1%
#630270000000
0!
0%
#630275000000
1!
1%
#630280000000
0!
0%
#630285000000
1!
1%
#630290000000
0!
0%
#630295000000
1!
1%
#630300000000
0!
0%
#630305000000
1!
1%
#630310000000
0!
0%
#630315000000
1!
1%
#630320000000
0!
0%
#630325000000
1!
1%
#630330000000
0!
0%
#630335000000
1!
1%
#630340000000
0!
0%
#630345000000
1!
1%
#630350000000
0!
0%
#630355000000
1!
1%
#630360000000
0!
0%
#630365000000
1!
1%
#630370000000
0!
0%
#630375000000
1!
1%
#630380000000
0!
0%
#630385000000
1!
1%
#630390000000
0!
0%
#630395000000
1!
1%
#630400000000
0!
0%
#630405000000
1!
1%
#630410000000
0!
0%
#630415000000
1!
1%
#630420000000
0!
0%
#630425000000
1!
1%
#630430000000
0!
0%
#630435000000
1!
1%
#630440000000
0!
0%
#630445000000
1!
1%
#630450000000
0!
0%
#630455000000
1!
1%
#630460000000
0!
0%
#630465000000
1!
1%
#630470000000
0!
0%
#630475000000
1!
1%
#630480000000
0!
0%
#630485000000
1!
1%
#630490000000
0!
0%
#630495000000
1!
1%
#630500000000
0!
0%
#630505000000
1!
1%
#630510000000
0!
0%
#630515000000
1!
1%
#630520000000
0!
0%
#630525000000
1!
1%
#630530000000
0!
0%
#630535000000
1!
1%
#630540000000
0!
0%
#630545000000
1!
1%
#630550000000
0!
0%
#630555000000
1!
1%
#630560000000
0!
0%
#630565000000
1!
1%
#630570000000
0!
0%
#630575000000
1!
1%
#630580000000
0!
0%
#630585000000
1!
1%
#630590000000
0!
0%
#630595000000
1!
1%
#630600000000
0!
0%
#630605000000
1!
1%
#630610000000
0!
0%
#630615000000
1!
1%
#630620000000
0!
0%
#630625000000
1!
1%
#630630000000
0!
0%
#630635000000
1!
1%
#630640000000
0!
0%
#630645000000
1!
1%
#630650000000
0!
0%
#630655000000
1!
1%
#630660000000
0!
0%
#630665000000
1!
1%
#630670000000
0!
0%
#630675000000
1!
1%
#630680000000
0!
0%
#630685000000
1!
1%
#630690000000
0!
0%
#630695000000
1!
1%
#630700000000
0!
0%
#630705000000
1!
1%
#630710000000
0!
0%
#630715000000
1!
1%
#630720000000
0!
0%
#630725000000
1!
1%
#630730000000
0!
0%
#630735000000
1!
1%
#630740000000
0!
0%
#630745000000
1!
1%
#630750000000
0!
0%
#630755000000
1!
1%
#630760000000
0!
0%
#630765000000
1!
1%
#630770000000
0!
0%
#630775000000
1!
1%
#630780000000
0!
0%
#630785000000
1!
1%
#630790000000
0!
0%
#630795000000
1!
1%
#630800000000
0!
0%
#630805000000
1!
1%
#630810000000
0!
0%
#630815000000
1!
1%
#630820000000
0!
0%
#630825000000
1!
1%
#630830000000
0!
0%
#630835000000
1!
1%
#630840000000
0!
0%
#630845000000
1!
1%
#630850000000
0!
0%
#630855000000
1!
1%
#630860000000
0!
0%
#630865000000
1!
1%
#630870000000
0!
0%
#630875000000
1!
1%
#630880000000
0!
0%
#630885000000
1!
1%
#630890000000
0!
0%
#630895000000
1!
1%
#630900000000
0!
0%
#630905000000
1!
1%
#630910000000
0!
0%
#630915000000
1!
1%
#630920000000
0!
0%
#630925000000
1!
1%
#630930000000
0!
0%
#630935000000
1!
1%
#630940000000
0!
0%
#630945000000
1!
1%
#630950000000
0!
0%
#630955000000
1!
1%
#630960000000
0!
0%
#630965000000
1!
1%
#630970000000
0!
0%
#630975000000
1!
1%
#630980000000
0!
0%
#630985000000
1!
1%
#630990000000
0!
0%
#630995000000
1!
1%
#631000000000
0!
0%
#631005000000
1!
1%
#631010000000
0!
0%
#631015000000
1!
1%
#631020000000
0!
0%
#631025000000
1!
1%
#631030000000
0!
0%
#631035000000
1!
1%
#631040000000
0!
0%
#631045000000
1!
1%
#631050000000
0!
0%
#631055000000
1!
1%
#631060000000
0!
0%
#631065000000
1!
1%
#631070000000
0!
0%
#631075000000
1!
1%
#631080000000
0!
0%
#631085000000
1!
1%
#631090000000
0!
0%
#631095000000
1!
1%
#631100000000
0!
0%
#631105000000
1!
1%
#631110000000
0!
0%
#631115000000
1!
1%
#631120000000
0!
0%
#631125000000
1!
1%
#631130000000
0!
0%
#631135000000
1!
1%
#631140000000
0!
0%
#631145000000
1!
1%
#631150000000
0!
0%
#631155000000
1!
1%
#631160000000
0!
0%
#631165000000
1!
1%
#631170000000
0!
0%
#631175000000
1!
1%
#631180000000
0!
0%
#631185000000
1!
1%
#631190000000
0!
0%
#631195000000
1!
1%
#631200000000
0!
0%
#631205000000
1!
1%
#631210000000
0!
0%
#631215000000
1!
1%
#631220000000
0!
0%
#631225000000
1!
1%
#631230000000
0!
0%
#631235000000
1!
1%
#631240000000
0!
0%
#631245000000
1!
1%
#631250000000
0!
0%
#631255000000
1!
1%
#631260000000
0!
0%
#631265000000
1!
1%
#631270000000
0!
0%
#631275000000
1!
1%
#631280000000
0!
0%
#631285000000
1!
1%
#631290000000
0!
0%
#631295000000
1!
1%
#631300000000
0!
0%
#631305000000
1!
1%
#631310000000
0!
0%
#631315000000
1!
1%
#631320000000
0!
0%
#631325000000
1!
1%
#631330000000
0!
0%
#631335000000
1!
1%
#631340000000
0!
0%
#631345000000
1!
1%
#631350000000
0!
0%
#631355000000
1!
1%
#631360000000
0!
0%
#631365000000
1!
1%
#631370000000
0!
0%
#631375000000
1!
1%
#631380000000
0!
0%
#631385000000
1!
1%
#631390000000
0!
0%
#631395000000
1!
1%
#631400000000
0!
0%
#631405000000
1!
1%
#631410000000
0!
0%
#631415000000
1!
1%
#631420000000
0!
0%
#631425000000
1!
1%
#631430000000
0!
0%
#631435000000
1!
1%
#631440000000
0!
0%
#631445000000
1!
1%
#631450000000
0!
0%
#631455000000
1!
1%
#631460000000
0!
0%
#631465000000
1!
1%
#631470000000
0!
0%
#631475000000
1!
1%
#631480000000
0!
0%
#631485000000
1!
1%
#631490000000
0!
0%
#631495000000
1!
1%
#631500000000
0!
0%
#631505000000
1!
1%
#631510000000
0!
0%
#631515000000
1!
1%
#631520000000
0!
0%
#631525000000
1!
1%
#631530000000
0!
0%
#631535000000
1!
1%
#631540000000
0!
0%
#631545000000
1!
1%
#631550000000
0!
0%
#631555000000
1!
1%
#631560000000
0!
0%
#631565000000
1!
1%
#631570000000
0!
0%
#631575000000
1!
1%
#631580000000
0!
0%
#631585000000
1!
1%
#631590000000
0!
0%
#631595000000
1!
1%
#631600000000
0!
0%
#631605000000
1!
1%
#631610000000
0!
0%
#631615000000
1!
1%
#631620000000
0!
0%
#631625000000
1!
1%
#631630000000
0!
0%
#631635000000
1!
1%
#631640000000
0!
0%
#631645000000
1!
1%
#631650000000
0!
0%
#631655000000
1!
1%
#631660000000
0!
0%
#631665000000
1!
1%
#631670000000
0!
0%
#631675000000
1!
1%
#631680000000
0!
0%
#631685000000
1!
1%
#631690000000
0!
0%
#631695000000
1!
1%
#631700000000
0!
0%
#631705000000
1!
1%
#631710000000
0!
0%
#631715000000
1!
1%
#631720000000
0!
0%
#631725000000
1!
1%
#631730000000
0!
0%
#631735000000
1!
1%
#631740000000
0!
0%
#631745000000
1!
1%
#631750000000
0!
0%
#631755000000
1!
1%
#631760000000
0!
0%
#631765000000
1!
1%
#631770000000
0!
0%
#631775000000
1!
1%
#631780000000
0!
0%
#631785000000
1!
1%
#631790000000
0!
0%
#631795000000
1!
1%
#631800000000
0!
0%
#631805000000
1!
1%
#631810000000
0!
0%
#631815000000
1!
1%
#631820000000
0!
0%
#631825000000
1!
1%
#631830000000
0!
0%
#631835000000
1!
1%
#631840000000
0!
0%
#631845000000
1!
1%
#631850000000
0!
0%
#631855000000
1!
1%
#631860000000
0!
0%
#631865000000
1!
1%
#631870000000
0!
0%
#631875000000
1!
1%
#631880000000
0!
0%
#631885000000
1!
1%
#631890000000
0!
0%
#631895000000
1!
1%
#631900000000
0!
0%
#631905000000
1!
1%
#631910000000
0!
0%
#631915000000
1!
1%
#631920000000
0!
0%
#631925000000
1!
1%
#631930000000
0!
0%
#631935000000
1!
1%
#631940000000
0!
0%
#631945000000
1!
1%
#631950000000
0!
0%
#631955000000
1!
1%
#631960000000
0!
0%
#631965000000
1!
1%
#631970000000
0!
0%
#631975000000
1!
1%
#631980000000
0!
0%
#631985000000
1!
1%
#631990000000
0!
0%
#631995000000
1!
1%
#632000000000
0!
0%
#632005000000
1!
1%
#632010000000
0!
0%
#632015000000
1!
1%
#632020000000
0!
0%
#632025000000
1!
1%
#632030000000
0!
0%
#632035000000
1!
1%
#632040000000
0!
0%
#632045000000
1!
1%
#632050000000
0!
0%
#632055000000
1!
1%
#632060000000
0!
0%
#632065000000
1!
1%
#632070000000
0!
0%
#632075000000
1!
1%
#632080000000
0!
0%
#632085000000
1!
1%
#632090000000
0!
0%
#632095000000
1!
1%
#632100000000
0!
0%
#632105000000
1!
1%
#632110000000
0!
0%
#632115000000
1!
1%
#632120000000
0!
0%
#632125000000
1!
1%
#632130000000
0!
0%
#632135000000
1!
1%
#632140000000
0!
0%
#632145000000
1!
1%
#632150000000
0!
0%
#632155000000
1!
1%
#632160000000
0!
0%
#632165000000
1!
1%
#632170000000
0!
0%
#632175000000
1!
1%
#632180000000
0!
0%
#632185000000
1!
1%
#632190000000
0!
0%
#632195000000
1!
1%
#632200000000
0!
0%
#632205000000
1!
1%
#632210000000
0!
0%
#632215000000
1!
1%
#632220000000
0!
0%
#632225000000
1!
1%
#632230000000
0!
0%
#632235000000
1!
1%
#632240000000
0!
0%
#632245000000
1!
1%
#632250000000
0!
0%
#632255000000
1!
1%
#632260000000
0!
0%
#632265000000
1!
1%
#632270000000
0!
0%
#632275000000
1!
1%
#632280000000
0!
0%
#632285000000
1!
1%
#632290000000
0!
0%
#632295000000
1!
1%
#632300000000
0!
0%
#632305000000
1!
1%
#632310000000
0!
0%
#632315000000
1!
1%
#632320000000
0!
0%
#632325000000
1!
1%
#632330000000
0!
0%
#632335000000
1!
1%
#632340000000
0!
0%
#632345000000
1!
1%
#632350000000
0!
0%
#632355000000
1!
1%
#632360000000
0!
0%
#632365000000
1!
1%
#632370000000
0!
0%
#632375000000
1!
1%
#632380000000
0!
0%
#632385000000
1!
1%
#632390000000
0!
0%
#632395000000
1!
1%
#632400000000
0!
0%
#632405000000
1!
1%
#632410000000
0!
0%
#632415000000
1!
1%
#632420000000
0!
0%
#632425000000
1!
1%
#632430000000
0!
0%
#632435000000
1!
1%
#632440000000
0!
0%
#632445000000
1!
1%
#632450000000
0!
0%
#632455000000
1!
1%
#632460000000
0!
0%
#632465000000
1!
1%
#632470000000
0!
0%
#632475000000
1!
1%
#632480000000
0!
0%
#632485000000
1!
1%
#632490000000
0!
0%
#632495000000
1!
1%
#632500000000
0!
0%
#632505000000
1!
1%
#632510000000
0!
0%
#632515000000
1!
1%
#632520000000
0!
0%
#632525000000
1!
1%
#632530000000
0!
0%
#632535000000
1!
1%
#632540000000
0!
0%
#632545000000
1!
1%
#632550000000
0!
0%
#632555000000
1!
1%
#632560000000
0!
0%
#632565000000
1!
1%
#632570000000
0!
0%
#632575000000
1!
1%
#632580000000
0!
0%
#632585000000
1!
1%
#632590000000
0!
0%
#632595000000
1!
1%
#632600000000
0!
0%
#632605000000
1!
1%
#632610000000
0!
0%
#632615000000
1!
1%
#632620000000
0!
0%
#632625000000
1!
1%
#632630000000
0!
0%
#632635000000
1!
1%
#632640000000
0!
0%
#632645000000
1!
1%
#632650000000
0!
0%
#632655000000
1!
1%
#632660000000
0!
0%
#632665000000
1!
1%
#632670000000
0!
0%
#632675000000
1!
1%
#632680000000
0!
0%
#632685000000
1!
1%
#632690000000
0!
0%
#632695000000
1!
1%
#632700000000
0!
0%
#632705000000
1!
1%
#632710000000
0!
0%
#632715000000
1!
1%
#632720000000
0!
0%
#632725000000
1!
1%
#632730000000
0!
0%
#632735000000
1!
1%
#632740000000
0!
0%
#632745000000
1!
1%
#632750000000
0!
0%
#632755000000
1!
1%
#632760000000
0!
0%
#632765000000
1!
1%
#632770000000
0!
0%
#632775000000
1!
1%
#632780000000
0!
0%
#632785000000
1!
1%
#632790000000
0!
0%
#632795000000
1!
1%
#632800000000
0!
0%
#632805000000
1!
1%
#632810000000
0!
0%
#632815000000
1!
1%
#632820000000
0!
0%
#632825000000
1!
1%
#632830000000
0!
0%
#632835000000
1!
1%
#632840000000
0!
0%
#632845000000
1!
1%
#632850000000
0!
0%
#632855000000
1!
1%
#632860000000
0!
0%
#632865000000
1!
1%
#632870000000
0!
0%
#632875000000
1!
1%
#632880000000
0!
0%
#632885000000
1!
1%
#632890000000
0!
0%
#632895000000
1!
1%
#632900000000
0!
0%
#632905000000
1!
1%
#632910000000
0!
0%
#632915000000
1!
1%
#632920000000
0!
0%
#632925000000
1!
1%
#632930000000
0!
0%
#632935000000
1!
1%
#632940000000
0!
0%
#632945000000
1!
1%
#632950000000
0!
0%
#632955000000
1!
1%
#632960000000
0!
0%
#632965000000
1!
1%
#632970000000
0!
0%
#632975000000
1!
1%
#632980000000
0!
0%
#632985000000
1!
1%
#632990000000
0!
0%
#632995000000
1!
1%
#633000000000
0!
0%
#633005000000
1!
1%
#633010000000
0!
0%
#633015000000
1!
1%
#633020000000
0!
0%
#633025000000
1!
1%
#633030000000
0!
0%
#633035000000
1!
1%
#633040000000
0!
0%
#633045000000
1!
1%
#633050000000
0!
0%
#633055000000
1!
1%
#633060000000
0!
0%
#633065000000
1!
1%
#633070000000
0!
0%
#633075000000
1!
1%
#633080000000
0!
0%
#633085000000
1!
1%
#633090000000
0!
0%
#633095000000
1!
1%
#633100000000
0!
0%
#633105000000
1!
1%
#633110000000
0!
0%
#633115000000
1!
1%
#633120000000
0!
0%
#633125000000
1!
1%
#633130000000
0!
0%
#633135000000
1!
1%
#633140000000
0!
0%
#633145000000
1!
1%
#633150000000
0!
0%
#633155000000
1!
1%
#633160000000
0!
0%
#633165000000
1!
1%
#633170000000
0!
0%
#633175000000
1!
1%
#633180000000
0!
0%
#633185000000
1!
1%
#633190000000
0!
0%
#633195000000
1!
1%
#633200000000
0!
0%
#633205000000
1!
1%
#633210000000
0!
0%
#633215000000
1!
1%
#633220000000
0!
0%
#633225000000
1!
1%
#633230000000
0!
0%
#633235000000
1!
1%
#633240000000
0!
0%
#633245000000
1!
1%
#633250000000
0!
0%
#633255000000
1!
1%
#633260000000
0!
0%
#633265000000
1!
1%
#633270000000
0!
0%
#633275000000
1!
1%
#633280000000
0!
0%
#633285000000
1!
1%
#633290000000
0!
0%
#633295000000
1!
1%
#633300000000
0!
0%
#633305000000
1!
1%
#633310000000
0!
0%
#633315000000
1!
1%
#633320000000
0!
0%
#633325000000
1!
1%
#633330000000
0!
0%
#633335000000
1!
1%
#633340000000
0!
0%
#633345000000
1!
1%
#633350000000
0!
0%
#633355000000
1!
1%
#633360000000
0!
0%
#633365000000
1!
1%
#633370000000
0!
0%
#633375000000
1!
1%
#633380000000
0!
0%
#633385000000
1!
1%
#633390000000
0!
0%
#633395000000
1!
1%
#633400000000
0!
0%
#633405000000
1!
1%
#633410000000
0!
0%
#633415000000
1!
1%
#633420000000
0!
0%
#633425000000
1!
1%
#633430000000
0!
0%
#633435000000
1!
1%
#633440000000
0!
0%
#633445000000
1!
1%
#633450000000
0!
0%
#633455000000
1!
1%
#633460000000
0!
0%
#633465000000
1!
1%
#633470000000
0!
0%
#633475000000
1!
1%
#633480000000
0!
0%
#633485000000
1!
1%
#633490000000
0!
0%
#633495000000
1!
1%
#633500000000
0!
0%
#633505000000
1!
1%
#633510000000
0!
0%
#633515000000
1!
1%
#633520000000
0!
0%
#633525000000
1!
1%
#633530000000
0!
0%
#633535000000
1!
1%
#633540000000
0!
0%
#633545000000
1!
1%
#633550000000
0!
0%
#633555000000
1!
1%
#633560000000
0!
0%
#633565000000
1!
1%
#633570000000
0!
0%
#633575000000
1!
1%
#633580000000
0!
0%
#633585000000
1!
1%
#633590000000
0!
0%
#633595000000
1!
1%
#633600000000
0!
0%
#633605000000
1!
1%
#633610000000
0!
0%
#633615000000
1!
1%
#633620000000
0!
0%
#633625000000
1!
1%
#633630000000
0!
0%
#633635000000
1!
1%
#633640000000
0!
0%
#633645000000
1!
1%
#633650000000
0!
0%
#633655000000
1!
1%
#633660000000
0!
0%
#633665000000
1!
1%
#633670000000
0!
0%
#633675000000
1!
1%
#633680000000
0!
0%
#633685000000
1!
1%
#633690000000
0!
0%
#633695000000
1!
1%
#633700000000
0!
0%
#633705000000
1!
1%
#633710000000
0!
0%
#633715000000
1!
1%
#633720000000
0!
0%
#633725000000
1!
1%
#633730000000
0!
0%
#633735000000
1!
1%
#633740000000
0!
0%
#633745000000
1!
1%
#633750000000
0!
0%
#633755000000
1!
1%
#633760000000
0!
0%
#633765000000
1!
1%
#633770000000
0!
0%
#633775000000
1!
1%
#633780000000
0!
0%
#633785000000
1!
1%
#633790000000
0!
0%
#633795000000
1!
1%
#633800000000
0!
0%
#633805000000
1!
1%
#633810000000
0!
0%
#633815000000
1!
1%
#633820000000
0!
0%
#633825000000
1!
1%
#633830000000
0!
0%
#633835000000
1!
1%
#633840000000
0!
0%
#633845000000
1!
1%
#633850000000
0!
0%
#633855000000
1!
1%
#633860000000
0!
0%
#633865000000
1!
1%
#633870000000
0!
0%
#633875000000
1!
1%
#633880000000
0!
0%
#633885000000
1!
1%
#633890000000
0!
0%
#633895000000
1!
1%
#633900000000
0!
0%
#633905000000
1!
1%
#633910000000
0!
0%
#633915000000
1!
1%
#633920000000
0!
0%
#633925000000
1!
1%
#633930000000
0!
0%
#633935000000
1!
1%
#633940000000
0!
0%
#633945000000
1!
1%
#633950000000
0!
0%
#633955000000
1!
1%
#633960000000
0!
0%
#633965000000
1!
1%
#633970000000
0!
0%
#633975000000
1!
1%
#633980000000
0!
0%
#633985000000
1!
1%
#633990000000
0!
0%
#633995000000
1!
1%
#634000000000
0!
0%
#634005000000
1!
1%
#634010000000
0!
0%
#634015000000
1!
1%
#634020000000
0!
0%
#634025000000
1!
1%
#634030000000
0!
0%
#634035000000
1!
1%
#634040000000
0!
0%
#634045000000
1!
1%
#634050000000
0!
0%
#634055000000
1!
1%
#634060000000
0!
0%
#634065000000
1!
1%
#634070000000
0!
0%
#634075000000
1!
1%
#634080000000
0!
0%
#634085000000
1!
1%
#634090000000
0!
0%
#634095000000
1!
1%
#634100000000
0!
0%
#634105000000
1!
1%
#634110000000
0!
0%
#634115000000
1!
1%
#634120000000
0!
0%
#634125000000
1!
1%
#634130000000
0!
0%
#634135000000
1!
1%
#634140000000
0!
0%
#634145000000
1!
1%
#634150000000
0!
0%
#634155000000
1!
1%
#634160000000
0!
0%
#634165000000
1!
1%
#634170000000
0!
0%
#634175000000
1!
1%
#634180000000
0!
0%
#634185000000
1!
1%
#634190000000
0!
0%
#634195000000
1!
1%
#634200000000
0!
0%
#634205000000
1!
1%
#634210000000
0!
0%
#634215000000
1!
1%
#634220000000
0!
0%
#634225000000
1!
1%
#634230000000
0!
0%
#634235000000
1!
1%
#634240000000
0!
0%
#634245000000
1!
1%
#634250000000
0!
0%
#634255000000
1!
1%
#634260000000
0!
0%
#634265000000
1!
1%
#634270000000
0!
0%
#634275000000
1!
1%
#634280000000
0!
0%
#634285000000
1!
1%
#634290000000
0!
0%
#634295000000
1!
1%
#634300000000
0!
0%
#634305000000
1!
1%
#634310000000
0!
0%
#634315000000
1!
1%
#634320000000
0!
0%
#634325000000
1!
1%
#634330000000
0!
0%
#634335000000
1!
1%
#634340000000
0!
0%
#634345000000
1!
1%
#634350000000
0!
0%
#634355000000
1!
1%
#634360000000
0!
0%
#634365000000
1!
1%
#634370000000
0!
0%
#634375000000
1!
1%
#634380000000
0!
0%
#634385000000
1!
1%
#634390000000
0!
0%
#634395000000
1!
1%
#634400000000
0!
0%
#634405000000
1!
1%
#634410000000
0!
0%
#634415000000
1!
1%
#634420000000
0!
0%
#634425000000
1!
1%
#634430000000
0!
0%
#634435000000
1!
1%
#634440000000
0!
0%
#634445000000
1!
1%
#634450000000
0!
0%
#634455000000
1!
1%
#634460000000
0!
0%
#634465000000
1!
1%
#634470000000
0!
0%
#634475000000
1!
1%
#634480000000
0!
0%
#634485000000
1!
1%
#634490000000
0!
0%
#634495000000
1!
1%
#634500000000
0!
0%
#634505000000
1!
1%
#634510000000
0!
0%
#634515000000
1!
1%
#634520000000
0!
0%
#634525000000
1!
1%
#634530000000
0!
0%
#634535000000
1!
1%
#634540000000
0!
0%
#634545000000
1!
1%
#634550000000
0!
0%
#634555000000
1!
1%
#634560000000
0!
0%
#634565000000
1!
1%
#634570000000
0!
0%
#634575000000
1!
1%
#634580000000
0!
0%
#634585000000
1!
1%
#634590000000
0!
0%
#634595000000
1!
1%
#634600000000
0!
0%
#634605000000
1!
1%
#634610000000
0!
0%
#634615000000
1!
1%
#634620000000
0!
0%
#634625000000
1!
1%
#634630000000
0!
0%
#634635000000
1!
1%
#634640000000
0!
0%
#634645000000
1!
1%
#634650000000
0!
0%
#634655000000
1!
1%
#634660000000
0!
0%
#634665000000
1!
1%
#634670000000
0!
0%
#634675000000
1!
1%
#634680000000
0!
0%
#634685000000
1!
1%
#634690000000
0!
0%
#634695000000
1!
1%
#634700000000
0!
0%
#634705000000
1!
1%
#634710000000
0!
0%
#634715000000
1!
1%
#634720000000
0!
0%
#634725000000
1!
1%
#634730000000
0!
0%
#634735000000
1!
1%
#634740000000
0!
0%
#634745000000
1!
1%
#634750000000
0!
0%
#634755000000
1!
1%
#634760000000
0!
0%
#634765000000
1!
1%
#634770000000
0!
0%
#634775000000
1!
1%
#634780000000
0!
0%
#634785000000
1!
1%
#634790000000
0!
0%
#634795000000
1!
1%
#634800000000
0!
0%
#634805000000
1!
1%
#634810000000
0!
0%
#634815000000
1!
1%
#634820000000
0!
0%
#634825000000
1!
1%
#634830000000
0!
0%
#634835000000
1!
1%
#634840000000
0!
0%
#634845000000
1!
1%
#634850000000
0!
0%
#634855000000
1!
1%
#634860000000
0!
0%
#634865000000
1!
1%
#634870000000
0!
0%
#634875000000
1!
1%
#634880000000
0!
0%
#634885000000
1!
1%
#634890000000
0!
0%
#634895000000
1!
1%
#634900000000
0!
0%
#634905000000
1!
1%
#634910000000
0!
0%
#634915000000
1!
1%
#634920000000
0!
0%
#634925000000
1!
1%
#634930000000
0!
0%
#634935000000
1!
1%
#634940000000
0!
0%
#634945000000
1!
1%
#634950000000
0!
0%
#634955000000
1!
1%
#634960000000
0!
0%
#634965000000
1!
1%
#634970000000
0!
0%
#634975000000
1!
1%
#634980000000
0!
0%
#634985000000
1!
1%
#634990000000
0!
0%
#634995000000
1!
1%
#635000000000
0!
0%
#635005000000
1!
1%
#635010000000
0!
0%
#635015000000
1!
1%
#635020000000
0!
0%
#635025000000
1!
1%
#635030000000
0!
0%
#635035000000
1!
1%
#635040000000
0!
0%
#635045000000
1!
1%
#635050000000
0!
0%
#635055000000
1!
1%
#635060000000
0!
0%
#635065000000
1!
1%
#635070000000
0!
0%
#635075000000
1!
1%
#635080000000
0!
0%
#635085000000
1!
1%
#635090000000
0!
0%
#635095000000
1!
1%
#635100000000
0!
0%
#635105000000
1!
1%
#635110000000
0!
0%
#635115000000
1!
1%
#635120000000
0!
0%
#635125000000
1!
1%
#635130000000
0!
0%
#635135000000
1!
1%
#635140000000
0!
0%
#635145000000
1!
1%
#635150000000
0!
0%
#635155000000
1!
1%
#635160000000
0!
0%
#635165000000
1!
1%
#635170000000
0!
0%
#635175000000
1!
1%
#635180000000
0!
0%
#635185000000
1!
1%
#635190000000
0!
0%
#635195000000
1!
1%
#635200000000
0!
0%
#635205000000
1!
1%
#635210000000
0!
0%
#635215000000
1!
1%
#635220000000
0!
0%
#635225000000
1!
1%
#635230000000
0!
0%
#635235000000
1!
1%
#635240000000
0!
0%
#635245000000
1!
1%
#635250000000
0!
0%
#635255000000
1!
1%
#635260000000
0!
0%
#635265000000
1!
1%
#635270000000
0!
0%
#635275000000
1!
1%
#635280000000
0!
0%
#635285000000
1!
1%
#635290000000
0!
0%
#635295000000
1!
1%
#635300000000
0!
0%
#635305000000
1!
1%
#635310000000
0!
0%
#635315000000
1!
1%
#635320000000
0!
0%
#635325000000
1!
1%
#635330000000
0!
0%
#635335000000
1!
1%
#635340000000
0!
0%
#635345000000
1!
1%
#635350000000
0!
0%
#635355000000
1!
1%
#635360000000
0!
0%
#635365000000
1!
1%
#635370000000
0!
0%
#635375000000
1!
1%
#635380000000
0!
0%
#635385000000
1!
1%
#635390000000
0!
0%
#635395000000
1!
1%
#635400000000
0!
0%
#635405000000
1!
1%
#635410000000
0!
0%
#635415000000
1!
1%
#635420000000
0!
0%
#635425000000
1!
1%
#635430000000
0!
0%
#635435000000
1!
1%
#635440000000
0!
0%
#635445000000
1!
1%
#635450000000
0!
0%
#635455000000
1!
1%
#635460000000
0!
0%
#635465000000
1!
1%
#635470000000
0!
0%
#635475000000
1!
1%
#635480000000
0!
0%
#635485000000
1!
1%
#635490000000
0!
0%
#635495000000
1!
1%
#635500000000
0!
0%
#635505000000
1!
1%
#635510000000
0!
0%
#635515000000
1!
1%
#635520000000
0!
0%
#635525000000
1!
1%
#635530000000
0!
0%
#635535000000
1!
1%
#635540000000
0!
0%
#635545000000
1!
1%
#635550000000
0!
0%
#635555000000
1!
1%
#635560000000
0!
0%
#635565000000
1!
1%
#635570000000
0!
0%
#635575000000
1!
1%
#635580000000
0!
0%
#635585000000
1!
1%
#635590000000
0!
0%
#635595000000
1!
1%
#635600000000
0!
0%
#635605000000
1!
1%
#635610000000
0!
0%
#635615000000
1!
1%
#635620000000
0!
0%
#635625000000
1!
1%
#635630000000
0!
0%
#635635000000
1!
1%
#635640000000
0!
0%
#635645000000
1!
1%
#635650000000
0!
0%
#635655000000
1!
1%
#635660000000
0!
0%
#635665000000
1!
1%
#635670000000
0!
0%
#635675000000
1!
1%
#635680000000
0!
0%
#635685000000
1!
1%
#635690000000
0!
0%
#635695000000
1!
1%
#635700000000
0!
0%
#635705000000
1!
1%
#635710000000
0!
0%
#635715000000
1!
1%
#635720000000
0!
0%
#635725000000
1!
1%
#635730000000
0!
0%
#635735000000
1!
1%
#635740000000
0!
0%
#635745000000
1!
1%
#635750000000
0!
0%
#635755000000
1!
1%
#635760000000
0!
0%
#635765000000
1!
1%
#635770000000
0!
0%
#635775000000
1!
1%
#635780000000
0!
0%
#635785000000
1!
1%
#635790000000
0!
0%
#635795000000
1!
1%
#635800000000
0!
0%
#635805000000
1!
1%
#635810000000
0!
0%
#635815000000
1!
1%
#635820000000
0!
0%
#635825000000
1!
1%
#635830000000
0!
0%
#635835000000
1!
1%
#635840000000
0!
0%
#635845000000
1!
1%
#635850000000
0!
0%
#635855000000
1!
1%
#635860000000
0!
0%
#635865000000
1!
1%
#635870000000
0!
0%
#635875000000
1!
1%
#635880000000
0!
0%
#635885000000
1!
1%
#635890000000
0!
0%
#635895000000
1!
1%
#635900000000
0!
0%
#635905000000
1!
1%
#635910000000
0!
0%
#635915000000
1!
1%
#635920000000
0!
0%
#635925000000
1!
1%
#635930000000
0!
0%
#635935000000
1!
1%
#635940000000
0!
0%
#635945000000
1!
1%
#635950000000
0!
0%
#635955000000
1!
1%
#635960000000
0!
0%
#635965000000
1!
1%
#635970000000
0!
0%
#635975000000
1!
1%
#635980000000
0!
0%
#635985000000
1!
1%
#635990000000
0!
0%
#635995000000
1!
1%
#636000000000
0!
0%
#636005000000
1!
1%
#636010000000
0!
0%
#636015000000
1!
1%
#636020000000
0!
0%
#636025000000
1!
1%
#636030000000
0!
0%
#636035000000
1!
1%
#636040000000
0!
0%
#636045000000
1!
1%
#636050000000
0!
0%
#636055000000
1!
1%
#636060000000
0!
0%
#636065000000
1!
1%
#636070000000
0!
0%
#636075000000
1!
1%
#636080000000
0!
0%
#636085000000
1!
1%
#636090000000
0!
0%
#636095000000
1!
1%
#636100000000
0!
0%
#636105000000
1!
1%
#636110000000
0!
0%
#636115000000
1!
1%
#636120000000
0!
0%
#636125000000
1!
1%
#636130000000
0!
0%
#636135000000
1!
1%
#636140000000
0!
0%
#636145000000
1!
1%
#636150000000
0!
0%
#636155000000
1!
1%
#636160000000
0!
0%
#636165000000
1!
1%
#636170000000
0!
0%
#636175000000
1!
1%
#636180000000
0!
0%
#636185000000
1!
1%
#636190000000
0!
0%
#636195000000
1!
1%
#636200000000
0!
0%
#636205000000
1!
1%
#636210000000
0!
0%
#636215000000
1!
1%
#636220000000
0!
0%
#636225000000
1!
1%
#636230000000
0!
0%
#636235000000
1!
1%
#636240000000
0!
0%
#636245000000
1!
1%
#636250000000
0!
0%
#636255000000
1!
1%
#636260000000
0!
0%
#636265000000
1!
1%
#636270000000
0!
0%
#636275000000
1!
1%
#636280000000
0!
0%
#636285000000
1!
1%
#636290000000
0!
0%
#636295000000
1!
1%
#636300000000
0!
0%
#636305000000
1!
1%
#636310000000
0!
0%
#636315000000
1!
1%
#636320000000
0!
0%
#636325000000
1!
1%
#636330000000
0!
0%
#636335000000
1!
1%
#636340000000
0!
0%
#636345000000
1!
1%
#636350000000
0!
0%
#636355000000
1!
1%
#636360000000
0!
0%
#636365000000
1!
1%
#636370000000
0!
0%
#636375000000
1!
1%
#636380000000
0!
0%
#636385000000
1!
1%
#636390000000
0!
0%
#636395000000
1!
1%
#636400000000
0!
0%
#636405000000
1!
1%
#636410000000
0!
0%
#636415000000
1!
1%
#636420000000
0!
0%
#636425000000
1!
1%
#636430000000
0!
0%
#636435000000
1!
1%
#636440000000
0!
0%
#636445000000
1!
1%
#636450000000
0!
0%
#636455000000
1!
1%
#636460000000
0!
0%
#636465000000
1!
1%
#636470000000
0!
0%
#636475000000
1!
1%
#636480000000
0!
0%
#636485000000
1!
1%
#636490000000
0!
0%
#636495000000
1!
1%
#636500000000
0!
0%
#636505000000
1!
1%
#636510000000
0!
0%
#636515000000
1!
1%
#636520000000
0!
0%
#636525000000
1!
1%
#636530000000
0!
0%
#636535000000
1!
1%
#636540000000
0!
0%
#636545000000
1!
1%
#636550000000
0!
0%
#636555000000
1!
1%
#636560000000
0!
0%
#636565000000
1!
1%
#636570000000
0!
0%
#636575000000
1!
1%
#636580000000
0!
0%
#636585000000
1!
1%
#636590000000
0!
0%
#636595000000
1!
1%
#636600000000
0!
0%
#636605000000
1!
1%
#636610000000
0!
0%
#636615000000
1!
1%
#636620000000
0!
0%
#636625000000
1!
1%
#636630000000
0!
0%
#636635000000
1!
1%
#636640000000
0!
0%
#636645000000
1!
1%
#636650000000
0!
0%
#636655000000
1!
1%
#636660000000
0!
0%
#636665000000
1!
1%
#636670000000
0!
0%
#636675000000
1!
1%
#636680000000
0!
0%
#636685000000
1!
1%
#636690000000
0!
0%
#636695000000
1!
1%
#636700000000
0!
0%
#636705000000
1!
1%
#636710000000
0!
0%
#636715000000
1!
1%
#636720000000
0!
0%
#636725000000
1!
1%
#636730000000
0!
0%
#636735000000
1!
1%
#636740000000
0!
0%
#636745000000
1!
1%
#636750000000
0!
0%
#636755000000
1!
1%
#636760000000
0!
0%
#636765000000
1!
1%
#636770000000
0!
0%
#636775000000
1!
1%
#636780000000
0!
0%
#636785000000
1!
1%
#636790000000
0!
0%
#636795000000
1!
1%
#636800000000
0!
0%
#636805000000
1!
1%
#636810000000
0!
0%
#636815000000
1!
1%
#636820000000
0!
0%
#636825000000
1!
1%
#636830000000
0!
0%
#636835000000
1!
1%
#636840000000
0!
0%
#636845000000
1!
1%
#636850000000
0!
0%
#636855000000
1!
1%
#636860000000
0!
0%
#636865000000
1!
1%
#636870000000
0!
0%
#636875000000
1!
1%
#636880000000
0!
0%
#636885000000
1!
1%
#636890000000
0!
0%
#636895000000
1!
1%
#636900000000
0!
0%
#636905000000
1!
1%
#636910000000
0!
0%
#636915000000
1!
1%
#636920000000
0!
0%
#636925000000
1!
1%
#636930000000
0!
0%
#636935000000
1!
1%
#636940000000
0!
0%
#636945000000
1!
1%
#636950000000
0!
0%
#636955000000
1!
1%
#636960000000
0!
0%
#636965000000
1!
1%
#636970000000
0!
0%
#636975000000
1!
1%
#636980000000
0!
0%
#636985000000
1!
1%
#636990000000
0!
0%
#636995000000
1!
1%
#637000000000
0!
0%
#637005000000
1!
1%
#637010000000
0!
0%
#637015000000
1!
1%
#637020000000
0!
0%
#637025000000
1!
1%
#637030000000
0!
0%
#637035000000
1!
1%
#637040000000
0!
0%
#637045000000
1!
1%
#637050000000
0!
0%
#637055000000
1!
1%
#637060000000
0!
0%
#637065000000
1!
1%
#637070000000
0!
0%
#637075000000
1!
1%
#637080000000
0!
0%
#637085000000
1!
1%
#637090000000
0!
0%
#637095000000
1!
1%
#637100000000
0!
0%
#637105000000
1!
1%
#637110000000
0!
0%
#637115000000
1!
1%
#637120000000
0!
0%
#637125000000
1!
1%
#637130000000
0!
0%
#637135000000
1!
1%
#637140000000
0!
0%
#637145000000
1!
1%
#637150000000
0!
0%
#637155000000
1!
1%
#637160000000
0!
0%
#637165000000
1!
1%
#637170000000
0!
0%
#637175000000
1!
1%
#637180000000
0!
0%
#637185000000
1!
1%
#637190000000
0!
0%
#637195000000
1!
1%
#637200000000
0!
0%
#637205000000
1!
1%
#637210000000
0!
0%
#637215000000
1!
1%
#637220000000
0!
0%
#637225000000
1!
1%
#637230000000
0!
0%
#637235000000
1!
1%
#637240000000
0!
0%
#637245000000
1!
1%
#637250000000
0!
0%
#637255000000
1!
1%
#637260000000
0!
0%
#637265000000
1!
1%
#637270000000
0!
0%
#637275000000
1!
1%
#637280000000
0!
0%
#637285000000
1!
1%
#637290000000
0!
0%
#637295000000
1!
1%
#637300000000
0!
0%
#637305000000
1!
1%
#637310000000
0!
0%
#637315000000
1!
1%
#637320000000
0!
0%
#637325000000
1!
1%
#637330000000
0!
0%
#637335000000
1!
1%
#637340000000
0!
0%
#637345000000
1!
1%
#637350000000
0!
0%
#637355000000
1!
1%
#637360000000
0!
0%
#637365000000
1!
1%
#637370000000
0!
0%
#637375000000
1!
1%
#637380000000
0!
0%
#637385000000
1!
1%
#637390000000
0!
0%
#637395000000
1!
1%
#637400000000
0!
0%
#637405000000
1!
1%
#637410000000
0!
0%
#637415000000
1!
1%
#637420000000
0!
0%
#637425000000
1!
1%
#637430000000
0!
0%
#637435000000
1!
1%
#637440000000
0!
0%
#637445000000
1!
1%
#637450000000
0!
0%
#637455000000
1!
1%
#637460000000
0!
0%
#637465000000
1!
1%
#637470000000
0!
0%
#637475000000
1!
1%
#637480000000
0!
0%
#637485000000
1!
1%
#637490000000
0!
0%
#637495000000
1!
1%
#637500000000
0!
0%
#637505000000
1!
1%
#637510000000
0!
0%
#637515000000
1!
1%
#637520000000
0!
0%
#637525000000
1!
1%
#637530000000
0!
0%
#637535000000
1!
1%
#637540000000
0!
0%
#637545000000
1!
1%
#637550000000
0!
0%
#637555000000
1!
1%
#637560000000
0!
0%
#637565000000
1!
1%
#637570000000
0!
0%
#637575000000
1!
1%
#637580000000
0!
0%
#637585000000
1!
1%
#637590000000
0!
0%
#637595000000
1!
1%
#637600000000
0!
0%
#637605000000
1!
1%
#637610000000
0!
0%
#637615000000
1!
1%
#637620000000
0!
0%
#637625000000
1!
1%
#637630000000
0!
0%
#637635000000
1!
1%
#637640000000
0!
0%
#637645000000
1!
1%
#637650000000
0!
0%
#637655000000
1!
1%
#637660000000
0!
0%
#637665000000
1!
1%
#637670000000
0!
0%
#637675000000
1!
1%
#637680000000
0!
0%
#637685000000
1!
1%
#637690000000
0!
0%
#637695000000
1!
1%
#637700000000
0!
0%
#637705000000
1!
1%
#637710000000
0!
0%
#637715000000
1!
1%
#637720000000
0!
0%
#637725000000
1!
1%
#637730000000
0!
0%
#637735000000
1!
1%
#637740000000
0!
0%
#637745000000
1!
1%
#637750000000
0!
0%
#637755000000
1!
1%
#637760000000
0!
0%
#637765000000
1!
1%
#637770000000
0!
0%
#637775000000
1!
1%
#637780000000
0!
0%
#637785000000
1!
1%
#637790000000
0!
0%
#637795000000
1!
1%
#637800000000
0!
0%
#637805000000
1!
1%
#637810000000
0!
0%
#637815000000
1!
1%
#637820000000
0!
0%
#637825000000
1!
1%
#637830000000
0!
0%
#637835000000
1!
1%
#637840000000
0!
0%
#637845000000
1!
1%
#637850000000
0!
0%
#637855000000
1!
1%
#637860000000
0!
0%
#637865000000
1!
1%
#637870000000
0!
0%
#637875000000
1!
1%
#637880000000
0!
0%
#637885000000
1!
1%
#637890000000
0!
0%
#637895000000
1!
1%
#637900000000
0!
0%
#637905000000
1!
1%
#637910000000
0!
0%
#637915000000
1!
1%
#637920000000
0!
0%
#637925000000
1!
1%
#637930000000
0!
0%
#637935000000
1!
1%
#637940000000
0!
0%
#637945000000
1!
1%
#637950000000
0!
0%
#637955000000
1!
1%
#637960000000
0!
0%
#637965000000
1!
1%
#637970000000
0!
0%
#637975000000
1!
1%
#637980000000
0!
0%
#637985000000
1!
1%
#637990000000
0!
0%
#637995000000
1!
1%
#638000000000
0!
0%
#638005000000
1!
1%
#638010000000
0!
0%
#638015000000
1!
1%
#638020000000
0!
0%
#638025000000
1!
1%
#638030000000
0!
0%
#638035000000
1!
1%
#638040000000
0!
0%
#638045000000
1!
1%
#638050000000
0!
0%
#638055000000
1!
1%
#638060000000
0!
0%
#638065000000
1!
1%
#638070000000
0!
0%
#638075000000
1!
1%
#638080000000
0!
0%
#638085000000
1!
1%
#638090000000
0!
0%
#638095000000
1!
1%
#638100000000
0!
0%
#638105000000
1!
1%
#638110000000
0!
0%
#638115000000
1!
1%
#638120000000
0!
0%
#638125000000
1!
1%
#638130000000
0!
0%
#638135000000
1!
1%
#638140000000
0!
0%
#638145000000
1!
1%
#638150000000
0!
0%
#638155000000
1!
1%
#638160000000
0!
0%
#638165000000
1!
1%
#638170000000
0!
0%
#638175000000
1!
1%
#638180000000
0!
0%
#638185000000
1!
1%
#638190000000
0!
0%
#638195000000
1!
1%
#638200000000
0!
0%
#638205000000
1!
1%
#638210000000
0!
0%
#638215000000
1!
1%
#638220000000
0!
0%
#638225000000
1!
1%
#638230000000
0!
0%
#638235000000
1!
1%
#638240000000
0!
0%
#638245000000
1!
1%
#638250000000
0!
0%
#638255000000
1!
1%
#638260000000
0!
0%
#638265000000
1!
1%
#638270000000
0!
0%
#638275000000
1!
1%
#638280000000
0!
0%
#638285000000
1!
1%
#638290000000
0!
0%
#638295000000
1!
1%
#638300000000
0!
0%
#638305000000
1!
1%
#638310000000
0!
0%
#638315000000
1!
1%
#638320000000
0!
0%
#638325000000
1!
1%
#638330000000
0!
0%
#638335000000
1!
1%
#638340000000
0!
0%
#638345000000
1!
1%
#638350000000
0!
0%
#638355000000
1!
1%
#638360000000
0!
0%
#638365000000
1!
1%
#638370000000
0!
0%
#638375000000
1!
1%
#638380000000
0!
0%
#638385000000
1!
1%
#638390000000
0!
0%
#638395000000
1!
1%
#638400000000
0!
0%
#638405000000
1!
1%
#638410000000
0!
0%
#638415000000
1!
1%
#638420000000
0!
0%
#638425000000
1!
1%
#638430000000
0!
0%
#638435000000
1!
1%
#638440000000
0!
0%
#638445000000
1!
1%
#638450000000
0!
0%
#638455000000
1!
1%
#638460000000
0!
0%
#638465000000
1!
1%
#638470000000
0!
0%
#638475000000
1!
1%
#638480000000
0!
0%
#638485000000
1!
1%
#638490000000
0!
0%
#638495000000
1!
1%
#638500000000
0!
0%
#638505000000
1!
1%
#638510000000
0!
0%
#638515000000
1!
1%
#638520000000
0!
0%
#638525000000
1!
1%
#638530000000
0!
0%
#638535000000
1!
1%
#638540000000
0!
0%
#638545000000
1!
1%
#638550000000
0!
0%
#638555000000
1!
1%
#638560000000
0!
0%
#638565000000
1!
1%
#638570000000
0!
0%
#638575000000
1!
1%
#638580000000
0!
0%
#638585000000
1!
1%
#638590000000
0!
0%
#638595000000
1!
1%
#638600000000
0!
0%
#638605000000
1!
1%
#638610000000
0!
0%
#638615000000
1!
1%
#638620000000
0!
0%
#638625000000
1!
1%
#638630000000
0!
0%
#638635000000
1!
1%
#638640000000
0!
0%
#638645000000
1!
1%
#638650000000
0!
0%
#638655000000
1!
1%
#638660000000
0!
0%
#638665000000
1!
1%
#638670000000
0!
0%
#638675000000
1!
1%
#638680000000
0!
0%
#638685000000
1!
1%
#638690000000
0!
0%
#638695000000
1!
1%
#638700000000
0!
0%
#638705000000
1!
1%
#638710000000
0!
0%
#638715000000
1!
1%
#638720000000
0!
0%
#638725000000
1!
1%
#638730000000
0!
0%
#638735000000
1!
1%
#638740000000
0!
0%
#638745000000
1!
1%
#638750000000
0!
0%
#638755000000
1!
1%
#638760000000
0!
0%
#638765000000
1!
1%
#638770000000
0!
0%
#638775000000
1!
1%
#638780000000
0!
0%
#638785000000
1!
1%
#638790000000
0!
0%
#638795000000
1!
1%
#638800000000
0!
0%
#638805000000
1!
1%
#638810000000
0!
0%
#638815000000
1!
1%
#638820000000
0!
0%
#638825000000
1!
1%
#638830000000
0!
0%
#638835000000
1!
1%
#638840000000
0!
0%
#638845000000
1!
1%
#638850000000
0!
0%
#638855000000
1!
1%
#638860000000
0!
0%
#638865000000
1!
1%
#638870000000
0!
0%
#638875000000
1!
1%
#638880000000
0!
0%
#638885000000
1!
1%
#638890000000
0!
0%
#638895000000
1!
1%
#638900000000
0!
0%
#638905000000
1!
1%
#638910000000
0!
0%
#638915000000
1!
1%
#638920000000
0!
0%
#638925000000
1!
1%
#638930000000
0!
0%
#638935000000
1!
1%
#638940000000
0!
0%
#638945000000
1!
1%
#638950000000
0!
0%
#638955000000
1!
1%
#638960000000
0!
0%
#638965000000
1!
1%
#638970000000
0!
0%
#638975000000
1!
1%
#638980000000
0!
0%
#638985000000
1!
1%
#638990000000
0!
0%
#638995000000
1!
1%
#639000000000
0!
0%
#639005000000
1!
1%
#639010000000
0!
0%
#639015000000
1!
1%
#639020000000
0!
0%
#639025000000
1!
1%
#639030000000
0!
0%
#639035000000
1!
1%
#639040000000
0!
0%
#639045000000
1!
1%
#639050000000
0!
0%
#639055000000
1!
1%
#639060000000
0!
0%
#639065000000
1!
1%
#639070000000
0!
0%
#639075000000
1!
1%
#639080000000
0!
0%
#639085000000
1!
1%
#639090000000
0!
0%
#639095000000
1!
1%
#639100000000
0!
0%
#639105000000
1!
1%
#639110000000
0!
0%
#639115000000
1!
1%
#639120000000
0!
0%
#639125000000
1!
1%
#639130000000
0!
0%
#639135000000
1!
1%
#639140000000
0!
0%
#639145000000
1!
1%
#639150000000
0!
0%
#639155000000
1!
1%
#639160000000
0!
0%
#639165000000
1!
1%
#639170000000
0!
0%
#639175000000
1!
1%
#639180000000
0!
0%
#639185000000
1!
1%
#639190000000
0!
0%
#639195000000
1!
1%
#639200000000
0!
0%
#639205000000
1!
1%
#639210000000
0!
0%
#639215000000
1!
1%
#639220000000
0!
0%
#639225000000
1!
1%
#639230000000
0!
0%
#639235000000
1!
1%
#639240000000
0!
0%
#639245000000
1!
1%
#639250000000
0!
0%
#639255000000
1!
1%
#639260000000
0!
0%
#639265000000
1!
1%
#639270000000
0!
0%
#639275000000
1!
1%
#639280000000
0!
0%
#639285000000
1!
1%
#639290000000
0!
0%
#639295000000
1!
1%
#639300000000
0!
0%
#639305000000
1!
1%
#639310000000
0!
0%
#639315000000
1!
1%
#639320000000
0!
0%
#639325000000
1!
1%
#639330000000
0!
0%
#639335000000
1!
1%
#639340000000
0!
0%
#639345000000
1!
1%
#639350000000
0!
0%
#639355000000
1!
1%
#639360000000
0!
0%
#639365000000
1!
1%
#639370000000
0!
0%
#639375000000
1!
1%
#639380000000
0!
0%
#639385000000
1!
1%
#639390000000
0!
0%
#639395000000
1!
1%
#639400000000
0!
0%
#639405000000
1!
1%
#639410000000
0!
0%
#639415000000
1!
1%
#639420000000
0!
0%
#639425000000
1!
1%
#639430000000
0!
0%
#639435000000
1!
1%
#639440000000
0!
0%
#639445000000
1!
1%
#639450000000
0!
0%
#639455000000
1!
1%
#639460000000
0!
0%
#639465000000
1!
1%
#639470000000
0!
0%
#639475000000
1!
1%
#639480000000
0!
0%
#639485000000
1!
1%
#639490000000
0!
0%
#639495000000
1!
1%
#639500000000
0!
0%
#639505000000
1!
1%
#639510000000
0!
0%
#639515000000
1!
1%
#639520000000
0!
0%
#639525000000
1!
1%
#639530000000
0!
0%
#639535000000
1!
1%
#639540000000
0!
0%
#639545000000
1!
1%
#639550000000
0!
0%
#639555000000
1!
1%
#639560000000
0!
0%
#639565000000
1!
1%
#639570000000
0!
0%
#639575000000
1!
1%
#639580000000
0!
0%
#639585000000
1!
1%
#639590000000
0!
0%
#639595000000
1!
1%
#639600000000
0!
0%
#639605000000
1!
1%
#639610000000
0!
0%
#639615000000
1!
1%
#639620000000
0!
0%
#639625000000
1!
1%
#639630000000
0!
0%
#639635000000
1!
1%
#639640000000
0!
0%
#639645000000
1!
1%
#639650000000
0!
0%
#639655000000
1!
1%
#639660000000
0!
0%
#639665000000
1!
1%
#639670000000
0!
0%
#639675000000
1!
1%
#639680000000
0!
0%
#639685000000
1!
1%
#639690000000
0!
0%
#639695000000
1!
1%
#639700000000
0!
0%
#639705000000
1!
1%
#639710000000
0!
0%
#639715000000
1!
1%
#639720000000
0!
0%
#639725000000
1!
1%
#639730000000
0!
0%
#639735000000
1!
1%
#639740000000
0!
0%
#639745000000
1!
1%
#639750000000
0!
0%
#639755000000
1!
1%
#639760000000
0!
0%
#639765000000
1!
1%
#639770000000
0!
0%
#639775000000
1!
1%
#639780000000
0!
0%
#639785000000
1!
1%
#639790000000
0!
0%
#639795000000
1!
1%
#639800000000
0!
0%
#639805000000
1!
1%
#639810000000
0!
0%
#639815000000
1!
1%
#639820000000
0!
0%
#639825000000
1!
1%
#639830000000
0!
0%
#639835000000
1!
1%
#639840000000
0!
0%
#639845000000
1!
1%
#639850000000
0!
0%
#639855000000
1!
1%
#639860000000
0!
0%
#639865000000
1!
1%
#639870000000
0!
0%
#639875000000
1!
1%
#639880000000
0!
0%
#639885000000
1!
1%
#639890000000
0!
0%
#639895000000
1!
1%
#639900000000
0!
0%
#639905000000
1!
1%
#639910000000
0!
0%
#639915000000
1!
1%
#639920000000
0!
0%
#639925000000
1!
1%
#639930000000
0!
0%
#639935000000
1!
1%
#639940000000
0!
0%
#639945000000
1!
1%
#639950000000
0!
0%
#639955000000
1!
1%
#639960000000
0!
0%
#639965000000
1!
1%
#639970000000
0!
0%
#639975000000
1!
1%
#639980000000
0!
0%
#639985000000
1!
1%
#639990000000
0!
0%
#639995000000
1!
1%
#640000000000
0!
0%
#640005000000
1!
1%
#640010000000
0!
0%
#640015000000
1!
1%
#640020000000
0!
0%
#640025000000
1!
1%
#640030000000
0!
0%
#640035000000
1!
1%
#640040000000
0!
0%
#640045000000
1!
1%
#640050000000
0!
0%
#640055000000
1!
1%
#640060000000
0!
0%
#640065000000
1!
1%
#640070000000
0!
0%
#640075000000
1!
1%
#640080000000
0!
0%
#640085000000
1!
1%
#640090000000
0!
0%
#640095000000
1!
1%
#640100000000
0!
0%
#640105000000
1!
1%
#640110000000
0!
0%
#640115000000
1!
1%
#640120000000
0!
0%
#640125000000
1!
1%
#640130000000
0!
0%
#640135000000
1!
1%
#640140000000
0!
0%
#640145000000
1!
1%
#640150000000
0!
0%
#640155000000
1!
1%
#640160000000
0!
0%
#640165000000
1!
1%
#640170000000
0!
0%
#640175000000
1!
1%
#640180000000
0!
0%
#640185000000
1!
1%
#640190000000
0!
0%
#640195000000
1!
1%
#640200000000
0!
0%
#640205000000
1!
1%
#640210000000
0!
0%
#640215000000
1!
1%
#640220000000
0!
0%
#640225000000
1!
1%
#640230000000
0!
0%
#640235000000
1!
1%
#640240000000
0!
0%
#640245000000
1!
1%
#640250000000
0!
0%
#640255000000
1!
1%
#640260000000
0!
0%
#640265000000
1!
1%
#640270000000
0!
0%
#640275000000
1!
1%
#640280000000
0!
0%
#640285000000
1!
1%
#640290000000
0!
0%
#640295000000
1!
1%
#640300000000
0!
0%
#640305000000
1!
1%
#640310000000
0!
0%
#640315000000
1!
1%
#640320000000
0!
0%
#640325000000
1!
1%
#640330000000
0!
0%
#640335000000
1!
1%
#640340000000
0!
0%
#640345000000
1!
1%
#640350000000
0!
0%
#640355000000
1!
1%
#640360000000
0!
0%
#640365000000
1!
1%
#640370000000
0!
0%
#640375000000
1!
1%
#640380000000
0!
0%
#640385000000
1!
1%
#640390000000
0!
0%
#640395000000
1!
1%
#640400000000
0!
0%
#640405000000
1!
1%
#640410000000
0!
0%
#640415000000
1!
1%
#640420000000
0!
0%
#640425000000
1!
1%
#640430000000
0!
0%
#640435000000
1!
1%
#640440000000
0!
0%
#640445000000
1!
1%
#640450000000
0!
0%
#640455000000
1!
1%
#640460000000
0!
0%
#640465000000
1!
1%
#640470000000
0!
0%
#640475000000
1!
1%
#640480000000
0!
0%
#640485000000
1!
1%
#640490000000
0!
0%
#640495000000
1!
1%
#640500000000
0!
0%
#640505000000
1!
1%
#640510000000
0!
0%
#640515000000
1!
1%
#640520000000
0!
0%
#640525000000
1!
1%
#640530000000
0!
0%
#640535000000
1!
1%
#640540000000
0!
0%
#640545000000
1!
1%
#640550000000
0!
0%
#640555000000
1!
1%
#640560000000
0!
0%
#640565000000
1!
1%
#640570000000
0!
0%
#640575000000
1!
1%
#640580000000
0!
0%
#640585000000
1!
1%
#640590000000
0!
0%
#640595000000
1!
1%
#640600000000
0!
0%
#640605000000
1!
1%
#640610000000
0!
0%
#640615000000
1!
1%
#640620000000
0!
0%
#640625000000
1!
1%
#640630000000
0!
0%
#640635000000
1!
1%
#640640000000
0!
0%
#640645000000
1!
1%
#640650000000
0!
0%
#640655000000
1!
1%
#640660000000
0!
0%
#640665000000
1!
1%
#640670000000
0!
0%
#640675000000
1!
1%
#640680000000
0!
0%
#640685000000
1!
1%
#640690000000
0!
0%
#640695000000
1!
1%
#640700000000
0!
0%
#640705000000
1!
1%
#640710000000
0!
0%
#640715000000
1!
1%
#640720000000
0!
0%
#640725000000
1!
1%
#640730000000
0!
0%
#640735000000
1!
1%
#640740000000
0!
0%
#640745000000
1!
1%
#640750000000
0!
0%
#640755000000
1!
1%
#640760000000
0!
0%
#640765000000
1!
1%
#640770000000
0!
0%
#640775000000
1!
1%
#640780000000
0!
0%
#640785000000
1!
1%
#640790000000
0!
0%
#640795000000
1!
1%
#640800000000
0!
0%
#640805000000
1!
1%
#640810000000
0!
0%
#640815000000
1!
1%
#640820000000
0!
0%
#640825000000
1!
1%
#640830000000
0!
0%
#640835000000
1!
1%
#640840000000
0!
0%
#640845000000
1!
1%
#640850000000
0!
0%
#640855000000
1!
1%
#640860000000
0!
0%
#640865000000
1!
1%
#640870000000
0!
0%
#640875000000
1!
1%
#640880000000
0!
0%
#640885000000
1!
1%
#640890000000
0!
0%
#640895000000
1!
1%
#640900000000
0!
0%
#640905000000
1!
1%
#640910000000
0!
0%
#640915000000
1!
1%
#640920000000
0!
0%
#640925000000
1!
1%
#640930000000
0!
0%
#640935000000
1!
1%
#640940000000
0!
0%
#640945000000
1!
1%
#640950000000
0!
0%
#640955000000
1!
1%
#640960000000
0!
0%
#640965000000
1!
1%
#640970000000
0!
0%
#640975000000
1!
1%
#640980000000
0!
0%
#640985000000
1!
1%
#640990000000
0!
0%
#640995000000
1!
1%
#641000000000
0!
0%
#641005000000
1!
1%
#641010000000
0!
0%
#641015000000
1!
1%
#641020000000
0!
0%
#641025000000
1!
1%
#641030000000
0!
0%
#641035000000
1!
1%
#641040000000
0!
0%
#641045000000
1!
1%
#641050000000
0!
0%
#641055000000
1!
1%
#641060000000
0!
0%
#641065000000
1!
1%
#641070000000
0!
0%
#641075000000
1!
1%
#641080000000
0!
0%
#641085000000
1!
1%
#641090000000
0!
0%
#641095000000
1!
1%
#641100000000
0!
0%
#641105000000
1!
1%
#641110000000
0!
0%
#641115000000
1!
1%
#641120000000
0!
0%
#641125000000
1!
1%
#641130000000
0!
0%
#641135000000
1!
1%
#641140000000
0!
0%
#641145000000
1!
1%
#641150000000
0!
0%
#641155000000
1!
1%
#641160000000
0!
0%
#641165000000
1!
1%
#641170000000
0!
0%
#641175000000
1!
1%
#641180000000
0!
0%
#641185000000
1!
1%
#641190000000
0!
0%
#641195000000
1!
1%
#641200000000
0!
0%
#641205000000
1!
1%
#641210000000
0!
0%
#641215000000
1!
1%
#641220000000
0!
0%
#641225000000
1!
1%
#641230000000
0!
0%
#641235000000
1!
1%
#641240000000
0!
0%
#641245000000
1!
1%
#641250000000
0!
0%
#641255000000
1!
1%
#641260000000
0!
0%
#641265000000
1!
1%
#641270000000
0!
0%
#641275000000
1!
1%
#641280000000
0!
0%
#641285000000
1!
1%
#641290000000
0!
0%
#641295000000
1!
1%
#641300000000
0!
0%
#641305000000
1!
1%
#641310000000
0!
0%
#641315000000
1!
1%
#641320000000
0!
0%
#641325000000
1!
1%
#641330000000
0!
0%
#641335000000
1!
1%
#641340000000
0!
0%
#641345000000
1!
1%
#641350000000
0!
0%
#641355000000
1!
1%
#641360000000
0!
0%
#641365000000
1!
1%
#641370000000
0!
0%
#641375000000
1!
1%
#641380000000
0!
0%
#641385000000
1!
1%
#641390000000
0!
0%
#641395000000
1!
1%
#641400000000
0!
0%
#641405000000
1!
1%
#641410000000
0!
0%
#641415000000
1!
1%
#641420000000
0!
0%
#641425000000
1!
1%
#641430000000
0!
0%
#641435000000
1!
1%
#641440000000
0!
0%
#641445000000
1!
1%
#641450000000
0!
0%
#641455000000
1!
1%
#641460000000
0!
0%
#641465000000
1!
1%
#641470000000
0!
0%
#641475000000
1!
1%
#641480000000
0!
0%
#641485000000
1!
1%
#641490000000
0!
0%
#641495000000
1!
1%
#641500000000
0!
0%
#641505000000
1!
1%
#641510000000
0!
0%
#641515000000
1!
1%
#641520000000
0!
0%
#641525000000
1!
1%
#641530000000
0!
0%
#641535000000
1!
1%
#641540000000
0!
0%
#641545000000
1!
1%
#641550000000
0!
0%
#641555000000
1!
1%
#641560000000
0!
0%
#641565000000
1!
1%
#641570000000
0!
0%
#641575000000
1!
1%
#641580000000
0!
0%
#641585000000
1!
1%
#641590000000
0!
0%
#641595000000
1!
1%
#641600000000
0!
0%
#641605000000
1!
1%
#641610000000
0!
0%
#641615000000
1!
1%
#641620000000
0!
0%
#641625000000
1!
1%
#641630000000
0!
0%
#641635000000
1!
1%
#641640000000
0!
0%
#641645000000
1!
1%
#641650000000
0!
0%
#641655000000
1!
1%
#641660000000
0!
0%
#641665000000
1!
1%
#641670000000
0!
0%
#641675000000
1!
1%
#641680000000
0!
0%
#641685000000
1!
1%
#641690000000
0!
0%
#641695000000
1!
1%
#641700000000
0!
0%
#641705000000
1!
1%
#641710000000
0!
0%
#641715000000
1!
1%
#641720000000
0!
0%
#641725000000
1!
1%
#641730000000
0!
0%
#641735000000
1!
1%
#641740000000
0!
0%
#641745000000
1!
1%
#641750000000
0!
0%
#641755000000
1!
1%
#641760000000
0!
0%
#641765000000
1!
1%
#641770000000
0!
0%
#641775000000
1!
1%
#641780000000
0!
0%
#641785000000
1!
1%
#641790000000
0!
0%
#641795000000
1!
1%
#641800000000
0!
0%
#641805000000
1!
1%
#641810000000
0!
0%
#641815000000
1!
1%
#641820000000
0!
0%
#641825000000
1!
1%
#641830000000
0!
0%
#641835000000
1!
1%
#641840000000
0!
0%
#641845000000
1!
1%
#641850000000
0!
0%
#641855000000
1!
1%
#641860000000
0!
0%
#641865000000
1!
1%
#641870000000
0!
0%
#641875000000
1!
1%
#641880000000
0!
0%
#641885000000
1!
1%
#641890000000
0!
0%
#641895000000
1!
1%
#641900000000
0!
0%
#641905000000
1!
1%
#641910000000
0!
0%
#641915000000
1!
1%
#641920000000
0!
0%
#641925000000
1!
1%
#641930000000
0!
0%
#641935000000
1!
1%
#641940000000
0!
0%
#641945000000
1!
1%
#641950000000
0!
0%
#641955000000
1!
1%
#641960000000
0!
0%
#641965000000
1!
1%
#641970000000
0!
0%
#641975000000
1!
1%
#641980000000
0!
0%
#641985000000
1!
1%
#641990000000
0!
0%
#641995000000
1!
1%
#642000000000
0!
0%
#642005000000
1!
1%
#642010000000
0!
0%
#642015000000
1!
1%
#642020000000
0!
0%
#642025000000
1!
1%
#642030000000
0!
0%
#642035000000
1!
1%
#642040000000
0!
0%
#642045000000
1!
1%
#642050000000
0!
0%
#642055000000
1!
1%
#642060000000
0!
0%
#642065000000
1!
1%
#642070000000
0!
0%
#642075000000
1!
1%
#642080000000
0!
0%
#642085000000
1!
1%
#642090000000
0!
0%
#642095000000
1!
1%
#642100000000
0!
0%
#642105000000
1!
1%
#642110000000
0!
0%
#642115000000
1!
1%
#642120000000
0!
0%
#642125000000
1!
1%
#642130000000
0!
0%
#642135000000
1!
1%
#642140000000
0!
0%
#642145000000
1!
1%
#642150000000
0!
0%
#642155000000
1!
1%
#642160000000
0!
0%
#642165000000
1!
1%
#642170000000
0!
0%
#642175000000
1!
1%
#642180000000
0!
0%
#642185000000
1!
1%
#642190000000
0!
0%
#642195000000
1!
1%
#642200000000
0!
0%
#642205000000
1!
1%
#642210000000
0!
0%
#642215000000
1!
1%
#642220000000
0!
0%
#642225000000
1!
1%
#642230000000
0!
0%
#642235000000
1!
1%
#642240000000
0!
0%
#642245000000
1!
1%
#642250000000
0!
0%
#642255000000
1!
1%
#642260000000
0!
0%
#642265000000
1!
1%
#642270000000
0!
0%
#642275000000
1!
1%
#642280000000
0!
0%
#642285000000
1!
1%
#642290000000
0!
0%
#642295000000
1!
1%
#642300000000
0!
0%
#642305000000
1!
1%
#642310000000
0!
0%
#642315000000
1!
1%
#642320000000
0!
0%
#642325000000
1!
1%
#642330000000
0!
0%
#642335000000
1!
1%
#642340000000
0!
0%
#642345000000
1!
1%
#642350000000
0!
0%
#642355000000
1!
1%
#642360000000
0!
0%
#642365000000
1!
1%
#642370000000
0!
0%
#642375000000
1!
1%
#642380000000
0!
0%
#642385000000
1!
1%
#642390000000
0!
0%
#642395000000
1!
1%
#642400000000
0!
0%
#642405000000
1!
1%
#642410000000
0!
0%
#642415000000
1!
1%
#642420000000
0!
0%
#642425000000
1!
1%
#642430000000
0!
0%
#642435000000
1!
1%
#642440000000
0!
0%
#642445000000
1!
1%
#642450000000
0!
0%
#642455000000
1!
1%
#642460000000
0!
0%
#642465000000
1!
1%
#642470000000
0!
0%
#642475000000
1!
1%
#642480000000
0!
0%
#642485000000
1!
1%
#642490000000
0!
0%
#642495000000
1!
1%
#642500000000
0!
0%
#642505000000
1!
1%
#642510000000
0!
0%
#642515000000
1!
1%
#642520000000
0!
0%
#642525000000
1!
1%
#642530000000
0!
0%
#642535000000
1!
1%
#642540000000
0!
0%
#642545000000
1!
1%
#642550000000
0!
0%
#642555000000
1!
1%
#642560000000
0!
0%
#642565000000
1!
1%
#642570000000
0!
0%
#642575000000
1!
1%
#642580000000
0!
0%
#642585000000
1!
1%
#642590000000
0!
0%
#642595000000
1!
1%
#642600000000
0!
0%
#642605000000
1!
1%
#642610000000
0!
0%
#642615000000
1!
1%
#642620000000
0!
0%
#642625000000
1!
1%
#642630000000
0!
0%
#642635000000
1!
1%
#642640000000
0!
0%
#642645000000
1!
1%
#642650000000
0!
0%
#642655000000
1!
1%
#642660000000
0!
0%
#642665000000
1!
1%
#642670000000
0!
0%
#642675000000
1!
1%
#642680000000
0!
0%
#642685000000
1!
1%
#642690000000
0!
0%
#642695000000
1!
1%
#642700000000
0!
0%
#642705000000
1!
1%
#642710000000
0!
0%
#642715000000
1!
1%
#642720000000
0!
0%
#642725000000
1!
1%
#642730000000
0!
0%
#642735000000
1!
1%
#642740000000
0!
0%
#642745000000
1!
1%
#642750000000
0!
0%
#642755000000
1!
1%
#642760000000
0!
0%
#642765000000
1!
1%
#642770000000
0!
0%
#642775000000
1!
1%
#642780000000
0!
0%
#642785000000
1!
1%
#642790000000
0!
0%
#642795000000
1!
1%
#642800000000
0!
0%
#642805000000
1!
1%
#642810000000
0!
0%
#642815000000
1!
1%
#642820000000
0!
0%
#642825000000
1!
1%
#642830000000
0!
0%
#642835000000
1!
1%
#642840000000
0!
0%
#642845000000
1!
1%
#642850000000
0!
0%
#642855000000
1!
1%
#642860000000
0!
0%
#642865000000
1!
1%
#642870000000
0!
0%
#642875000000
1!
1%
#642880000000
0!
0%
#642885000000
1!
1%
#642890000000
0!
0%
#642895000000
1!
1%
#642900000000
0!
0%
#642905000000
1!
1%
#642910000000
0!
0%
#642915000000
1!
1%
#642920000000
0!
0%
#642925000000
1!
1%
#642930000000
0!
0%
#642935000000
1!
1%
#642940000000
0!
0%
#642945000000
1!
1%
#642950000000
0!
0%
#642955000000
1!
1%
#642960000000
0!
0%
#642965000000
1!
1%
#642970000000
0!
0%
#642975000000
1!
1%
#642980000000
0!
0%
#642985000000
1!
1%
#642990000000
0!
0%
#642995000000
1!
1%
#643000000000
0!
0%
#643005000000
1!
1%
#643010000000
0!
0%
#643015000000
1!
1%
#643020000000
0!
0%
#643025000000
1!
1%
#643030000000
0!
0%
#643035000000
1!
1%
#643040000000
0!
0%
#643045000000
1!
1%
#643050000000
0!
0%
#643055000000
1!
1%
#643060000000
0!
0%
#643065000000
1!
1%
#643070000000
0!
0%
#643075000000
1!
1%
#643080000000
0!
0%
#643085000000
1!
1%
#643090000000
0!
0%
#643095000000
1!
1%
#643100000000
0!
0%
#643105000000
1!
1%
#643110000000
0!
0%
#643115000000
1!
1%
#643120000000
0!
0%
#643125000000
1!
1%
#643130000000
0!
0%
#643135000000
1!
1%
#643140000000
0!
0%
#643145000000
1!
1%
#643150000000
0!
0%
#643155000000
1!
1%
#643160000000
0!
0%
#643165000000
1!
1%
#643170000000
0!
0%
#643175000000
1!
1%
#643180000000
0!
0%
#643185000000
1!
1%
#643190000000
0!
0%
#643195000000
1!
1%
#643200000000
0!
0%
#643205000000
1!
1%
#643210000000
0!
0%
#643215000000
1!
1%
#643220000000
0!
0%
#643225000000
1!
1%
#643230000000
0!
0%
#643235000000
1!
1%
#643240000000
0!
0%
#643245000000
1!
1%
#643250000000
0!
0%
#643255000000
1!
1%
#643260000000
0!
0%
#643265000000
1!
1%
#643270000000
0!
0%
#643275000000
1!
1%
#643280000000
0!
0%
#643285000000
1!
1%
#643290000000
0!
0%
#643295000000
1!
1%
#643300000000
0!
0%
#643305000000
1!
1%
#643310000000
0!
0%
#643315000000
1!
1%
#643320000000
0!
0%
#643325000000
1!
1%
#643330000000
0!
0%
#643335000000
1!
1%
#643340000000
0!
0%
#643345000000
1!
1%
#643350000000
0!
0%
#643355000000
1!
1%
#643360000000
0!
0%
#643365000000
1!
1%
#643370000000
0!
0%
#643375000000
1!
1%
#643380000000
0!
0%
#643385000000
1!
1%
#643390000000
0!
0%
#643395000000
1!
1%
#643400000000
0!
0%
#643405000000
1!
1%
#643410000000
0!
0%
#643415000000
1!
1%
#643420000000
0!
0%
#643425000000
1!
1%
#643430000000
0!
0%
#643435000000
1!
1%
#643440000000
0!
0%
#643445000000
1!
1%
#643450000000
0!
0%
#643455000000
1!
1%
#643460000000
0!
0%
#643465000000
1!
1%
#643470000000
0!
0%
#643475000000
1!
1%
#643480000000
0!
0%
#643485000000
1!
1%
#643490000000
0!
0%
#643495000000
1!
1%
#643500000000
0!
0%
#643505000000
1!
1%
#643510000000
0!
0%
#643515000000
1!
1%
#643520000000
0!
0%
#643525000000
1!
1%
#643530000000
0!
0%
#643535000000
1!
1%
#643540000000
0!
0%
#643545000000
1!
1%
#643550000000
0!
0%
#643555000000
1!
1%
#643560000000
0!
0%
#643565000000
1!
1%
#643570000000
0!
0%
#643575000000
1!
1%
#643580000000
0!
0%
#643585000000
1!
1%
#643590000000
0!
0%
#643595000000
1!
1%
#643600000000
0!
0%
#643605000000
1!
1%
#643610000000
0!
0%
#643615000000
1!
1%
#643620000000
0!
0%
#643625000000
1!
1%
#643630000000
0!
0%
#643635000000
1!
1%
#643640000000
0!
0%
#643645000000
1!
1%
#643650000000
0!
0%
#643655000000
1!
1%
#643660000000
0!
0%
#643665000000
1!
1%
#643670000000
0!
0%
#643675000000
1!
1%
#643680000000
0!
0%
#643685000000
1!
1%
#643690000000
0!
0%
#643695000000
1!
1%
#643700000000
0!
0%
#643705000000
1!
1%
#643710000000
0!
0%
#643715000000
1!
1%
#643720000000
0!
0%
#643725000000
1!
1%
#643730000000
0!
0%
#643735000000
1!
1%
#643740000000
0!
0%
#643745000000
1!
1%
#643750000000
0!
0%
#643755000000
1!
1%
#643760000000
0!
0%
#643765000000
1!
1%
#643770000000
0!
0%
#643775000000
1!
1%
#643780000000
0!
0%
#643785000000
1!
1%
#643790000000
0!
0%
#643795000000
1!
1%
#643800000000
0!
0%
#643805000000
1!
1%
#643810000000
0!
0%
#643815000000
1!
1%
#643820000000
0!
0%
#643825000000
1!
1%
#643830000000
0!
0%
#643835000000
1!
1%
#643840000000
0!
0%
#643845000000
1!
1%
#643850000000
0!
0%
#643855000000
1!
1%
#643860000000
0!
0%
#643865000000
1!
1%
#643870000000
0!
0%
#643875000000
1!
1%
#643880000000
0!
0%
#643885000000
1!
1%
#643890000000
0!
0%
#643895000000
1!
1%
#643900000000
0!
0%
#643905000000
1!
1%
#643910000000
0!
0%
#643915000000
1!
1%
#643920000000
0!
0%
#643925000000
1!
1%
#643930000000
0!
0%
#643935000000
1!
1%
#643940000000
0!
0%
#643945000000
1!
1%
#643950000000
0!
0%
#643955000000
1!
1%
#643960000000
0!
0%
#643965000000
1!
1%
#643970000000
0!
0%
#643975000000
1!
1%
#643980000000
0!
0%
#643985000000
1!
1%
#643990000000
0!
0%
#643995000000
1!
1%
#644000000000
0!
0%
#644005000000
1!
1%
#644010000000
0!
0%
#644015000000
1!
1%
#644020000000
0!
0%
#644025000000
1!
1%
#644030000000
0!
0%
#644035000000
1!
1%
#644040000000
0!
0%
#644045000000
1!
1%
#644050000000
0!
0%
#644055000000
1!
1%
#644060000000
0!
0%
#644065000000
1!
1%
#644070000000
0!
0%
#644075000000
1!
1%
#644080000000
0!
0%
#644085000000
1!
1%
#644090000000
0!
0%
#644095000000
1!
1%
#644100000000
0!
0%
#644105000000
1!
1%
#644110000000
0!
0%
#644115000000
1!
1%
#644120000000
0!
0%
#644125000000
1!
1%
#644130000000
0!
0%
#644135000000
1!
1%
#644140000000
0!
0%
#644145000000
1!
1%
#644150000000
0!
0%
#644155000000
1!
1%
#644160000000
0!
0%
#644165000000
1!
1%
#644170000000
0!
0%
#644175000000
1!
1%
#644180000000
0!
0%
#644185000000
1!
1%
#644190000000
0!
0%
#644195000000
1!
1%
#644200000000
0!
0%
#644205000000
1!
1%
#644210000000
0!
0%
#644215000000
1!
1%
#644220000000
0!
0%
#644225000000
1!
1%
#644230000000
0!
0%
#644235000000
1!
1%
#644240000000
0!
0%
#644245000000
1!
1%
#644250000000
0!
0%
#644255000000
1!
1%
#644260000000
0!
0%
#644265000000
1!
1%
#644270000000
0!
0%
#644275000000
1!
1%
#644280000000
0!
0%
#644285000000
1!
1%
#644290000000
0!
0%
#644295000000
1!
1%
#644300000000
0!
0%
#644305000000
1!
1%
#644310000000
0!
0%
#644315000000
1!
1%
#644320000000
0!
0%
#644325000000
1!
1%
#644330000000
0!
0%
#644335000000
1!
1%
#644340000000
0!
0%
#644345000000
1!
1%
#644350000000
0!
0%
#644355000000
1!
1%
#644360000000
0!
0%
#644365000000
1!
1%
#644370000000
0!
0%
#644375000000
1!
1%
#644380000000
0!
0%
#644385000000
1!
1%
#644390000000
0!
0%
#644395000000
1!
1%
#644400000000
0!
0%
#644405000000
1!
1%
#644410000000
0!
0%
#644415000000
1!
1%
#644420000000
0!
0%
#644425000000
1!
1%
#644430000000
0!
0%
#644435000000
1!
1%
#644440000000
0!
0%
#644445000000
1!
1%
#644450000000
0!
0%
#644455000000
1!
1%
#644460000000
0!
0%
#644465000000
1!
1%
#644470000000
0!
0%
#644475000000
1!
1%
#644480000000
0!
0%
#644485000000
1!
1%
#644490000000
0!
0%
#644495000000
1!
1%
#644500000000
0!
0%
#644505000000
1!
1%
#644510000000
0!
0%
#644515000000
1!
1%
#644520000000
0!
0%
#644525000000
1!
1%
#644530000000
0!
0%
#644535000000
1!
1%
#644540000000
0!
0%
#644545000000
1!
1%
#644550000000
0!
0%
#644555000000
1!
1%
#644560000000
0!
0%
#644565000000
1!
1%
#644570000000
0!
0%
#644575000000
1!
1%
#644580000000
0!
0%
#644585000000
1!
1%
#644590000000
0!
0%
#644595000000
1!
1%
#644600000000
0!
0%
#644605000000
1!
1%
#644610000000
0!
0%
#644615000000
1!
1%
#644620000000
0!
0%
#644625000000
1!
1%
#644630000000
0!
0%
#644635000000
1!
1%
#644640000000
0!
0%
#644645000000
1!
1%
#644650000000
0!
0%
#644655000000
1!
1%
#644660000000
0!
0%
#644665000000
1!
1%
#644670000000
0!
0%
#644675000000
1!
1%
#644680000000
0!
0%
#644685000000
1!
1%
#644690000000
0!
0%
#644695000000
1!
1%
#644700000000
0!
0%
#644705000000
1!
1%
#644710000000
0!
0%
#644715000000
1!
1%
#644720000000
0!
0%
#644725000000
1!
1%
#644730000000
0!
0%
#644735000000
1!
1%
#644740000000
0!
0%
#644745000000
1!
1%
#644750000000
0!
0%
#644755000000
1!
1%
#644760000000
0!
0%
#644765000000
1!
1%
#644770000000
0!
0%
#644775000000
1!
1%
#644780000000
0!
0%
#644785000000
1!
1%
#644790000000
0!
0%
#644795000000
1!
1%
#644800000000
0!
0%
#644805000000
1!
1%
#644810000000
0!
0%
#644815000000
1!
1%
#644820000000
0!
0%
#644825000000
1!
1%
#644830000000
0!
0%
#644835000000
1!
1%
#644840000000
0!
0%
#644845000000
1!
1%
#644850000000
0!
0%
#644855000000
1!
1%
#644860000000
0!
0%
#644865000000
1!
1%
#644870000000
0!
0%
#644875000000
1!
1%
#644880000000
0!
0%
#644885000000
1!
1%
#644890000000
0!
0%
#644895000000
1!
1%
#644900000000
0!
0%
#644905000000
1!
1%
#644910000000
0!
0%
#644915000000
1!
1%
#644920000000
0!
0%
#644925000000
1!
1%
#644930000000
0!
0%
#644935000000
1!
1%
#644940000000
0!
0%
#644945000000
1!
1%
#644950000000
0!
0%
#644955000000
1!
1%
#644960000000
0!
0%
#644965000000
1!
1%
#644970000000
0!
0%
#644975000000
1!
1%
#644980000000
0!
0%
#644985000000
1!
1%
#644990000000
0!
0%
#644995000000
1!
1%
#645000000000
0!
0%
#645005000000
1!
1%
#645010000000
0!
0%
#645015000000
1!
1%
#645020000000
0!
0%
#645025000000
1!
1%
#645030000000
0!
0%
#645035000000
1!
1%
#645040000000
0!
0%
#645045000000
1!
1%
#645050000000
0!
0%
#645055000000
1!
1%
#645060000000
0!
0%
#645065000000
1!
1%
#645070000000
0!
0%
#645075000000
1!
1%
#645080000000
0!
0%
#645085000000
1!
1%
#645090000000
0!
0%
#645095000000
1!
1%
#645100000000
0!
0%
#645105000000
1!
1%
#645110000000
0!
0%
#645115000000
1!
1%
#645120000000
0!
0%
#645125000000
1!
1%
#645130000000
0!
0%
#645135000000
1!
1%
#645140000000
0!
0%
#645145000000
1!
1%
#645150000000
0!
0%
#645155000000
1!
1%
#645160000000
0!
0%
#645165000000
1!
1%
#645170000000
0!
0%
#645175000000
1!
1%
#645180000000
0!
0%
#645185000000
1!
1%
#645190000000
0!
0%
#645195000000
1!
1%
#645200000000
0!
0%
#645205000000
1!
1%
#645210000000
0!
0%
#645215000000
1!
1%
#645220000000
0!
0%
#645225000000
1!
1%
#645230000000
0!
0%
#645235000000
1!
1%
#645240000000
0!
0%
#645245000000
1!
1%
#645250000000
0!
0%
#645255000000
1!
1%
#645260000000
0!
0%
#645265000000
1!
1%
#645270000000
0!
0%
#645275000000
1!
1%
#645280000000
0!
0%
#645285000000
1!
1%
#645290000000
0!
0%
#645295000000
1!
1%
#645300000000
0!
0%
#645305000000
1!
1%
#645310000000
0!
0%
#645315000000
1!
1%
#645320000000
0!
0%
#645325000000
1!
1%
#645330000000
0!
0%
#645335000000
1!
1%
#645340000000
0!
0%
#645345000000
1!
1%
#645350000000
0!
0%
#645355000000
1!
1%
#645360000000
0!
0%
#645365000000
1!
1%
#645370000000
0!
0%
#645375000000
1!
1%
#645380000000
0!
0%
#645385000000
1!
1%
#645390000000
0!
0%
#645395000000
1!
1%
#645400000000
0!
0%
#645405000000
1!
1%
#645410000000
0!
0%
#645415000000
1!
1%
#645420000000
0!
0%
#645425000000
1!
1%
#645430000000
0!
0%
#645435000000
1!
1%
#645440000000
0!
0%
#645445000000
1!
1%
#645450000000
0!
0%
#645455000000
1!
1%
#645460000000
0!
0%
#645465000000
1!
1%
#645470000000
0!
0%
#645475000000
1!
1%
#645480000000
0!
0%
#645485000000
1!
1%
#645490000000
0!
0%
#645495000000
1!
1%
#645500000000
0!
0%
#645505000000
1!
1%
#645510000000
0!
0%
#645515000000
1!
1%
#645520000000
0!
0%
#645525000000
1!
1%
#645530000000
0!
0%
#645535000000
1!
1%
#645540000000
0!
0%
#645545000000
1!
1%
#645550000000
0!
0%
#645555000000
1!
1%
#645560000000
0!
0%
#645565000000
1!
1%
#645570000000
0!
0%
#645575000000
1!
1%
#645580000000
0!
0%
#645585000000
1!
1%
#645590000000
0!
0%
#645595000000
1!
1%
#645600000000
0!
0%
#645605000000
1!
1%
#645610000000
0!
0%
#645615000000
1!
1%
#645620000000
0!
0%
#645625000000
1!
1%
#645630000000
0!
0%
#645635000000
1!
1%
#645640000000
0!
0%
#645645000000
1!
1%
#645650000000
0!
0%
#645655000000
1!
1%
#645660000000
0!
0%
#645665000000
1!
1%
#645670000000
0!
0%
#645675000000
1!
1%
#645680000000
0!
0%
#645685000000
1!
1%
#645690000000
0!
0%
#645695000000
1!
1%
#645700000000
0!
0%
#645705000000
1!
1%
#645710000000
0!
0%
#645715000000
1!
1%
#645720000000
0!
0%
#645725000000
1!
1%
#645730000000
0!
0%
#645735000000
1!
1%
#645740000000
0!
0%
#645745000000
1!
1%
#645750000000
0!
0%
#645755000000
1!
1%
#645760000000
0!
0%
#645765000000
1!
1%
#645770000000
0!
0%
#645775000000
1!
1%
#645780000000
0!
0%
#645785000000
1!
1%
#645790000000
0!
0%
#645795000000
1!
1%
#645800000000
0!
0%
#645805000000
1!
1%
#645810000000
0!
0%
#645815000000
1!
1%
#645820000000
0!
0%
#645825000000
1!
1%
#645830000000
0!
0%
#645835000000
1!
1%
#645840000000
0!
0%
#645845000000
1!
1%
#645850000000
0!
0%
#645855000000
1!
1%
#645860000000
0!
0%
#645865000000
1!
1%
#645870000000
0!
0%
#645875000000
1!
1%
#645880000000
0!
0%
#645885000000
1!
1%
#645890000000
0!
0%
#645895000000
1!
1%
#645900000000
0!
0%
#645905000000
1!
1%
#645910000000
0!
0%
#645915000000
1!
1%
#645920000000
0!
0%
#645925000000
1!
1%
#645930000000
0!
0%
#645935000000
1!
1%
#645940000000
0!
0%
#645945000000
1!
1%
#645950000000
0!
0%
#645955000000
1!
1%
#645960000000
0!
0%
#645965000000
1!
1%
#645970000000
0!
0%
#645975000000
1!
1%
#645980000000
0!
0%
#645985000000
1!
1%
#645990000000
0!
0%
#645995000000
1!
1%
#646000000000
0!
0%
#646005000000
1!
1%
#646010000000
0!
0%
#646015000000
1!
1%
#646020000000
0!
0%
#646025000000
1!
1%
#646030000000
0!
0%
#646035000000
1!
1%
#646040000000
0!
0%
#646045000000
1!
1%
#646050000000
0!
0%
#646055000000
1!
1%
#646060000000
0!
0%
#646065000000
1!
1%
#646070000000
0!
0%
#646075000000
1!
1%
#646080000000
0!
0%
#646085000000
1!
1%
#646090000000
0!
0%
#646095000000
1!
1%
#646100000000
0!
0%
#646105000000
1!
1%
#646110000000
0!
0%
#646115000000
1!
1%
#646120000000
0!
0%
#646125000000
1!
1%
#646130000000
0!
0%
#646135000000
1!
1%
#646140000000
0!
0%
#646145000000
1!
1%
#646150000000
0!
0%
#646155000000
1!
1%
#646160000000
0!
0%
#646165000000
1!
1%
#646170000000
0!
0%
#646175000000
1!
1%
#646180000000
0!
0%
#646185000000
1!
1%
#646190000000
0!
0%
#646195000000
1!
1%
#646200000000
0!
0%
#646205000000
1!
1%
#646210000000
0!
0%
#646215000000
1!
1%
#646220000000
0!
0%
#646225000000
1!
1%
#646230000000
0!
0%
#646235000000
1!
1%
#646240000000
0!
0%
#646245000000
1!
1%
#646250000000
0!
0%
#646255000000
1!
1%
#646260000000
0!
0%
#646265000000
1!
1%
#646270000000
0!
0%
#646275000000
1!
1%
#646280000000
0!
0%
#646285000000
1!
1%
#646290000000
0!
0%
#646295000000
1!
1%
#646300000000
0!
0%
#646305000000
1!
1%
#646310000000
0!
0%
#646315000000
1!
1%
#646320000000
0!
0%
#646325000000
1!
1%
#646330000000
0!
0%
#646335000000
1!
1%
#646340000000
0!
0%
#646345000000
1!
1%
#646350000000
0!
0%
#646355000000
1!
1%
#646360000000
0!
0%
#646365000000
1!
1%
#646370000000
0!
0%
#646375000000
1!
1%
#646380000000
0!
0%
#646385000000
1!
1%
#646390000000
0!
0%
#646395000000
1!
1%
#646400000000
0!
0%
#646405000000
1!
1%
#646410000000
0!
0%
#646415000000
1!
1%
#646420000000
0!
0%
#646425000000
1!
1%
#646430000000
0!
0%
#646435000000
1!
1%
#646440000000
0!
0%
#646445000000
1!
1%
#646450000000
0!
0%
#646455000000
1!
1%
#646460000000
0!
0%
#646465000000
1!
1%
#646470000000
0!
0%
#646475000000
1!
1%
#646480000000
0!
0%
#646485000000
1!
1%
#646490000000
0!
0%
#646495000000
1!
1%
#646500000000
0!
0%
#646505000000
1!
1%
#646510000000
0!
0%
#646515000000
1!
1%
#646520000000
0!
0%
#646525000000
1!
1%
#646530000000
0!
0%
#646535000000
1!
1%
#646540000000
0!
0%
#646545000000
1!
1%
#646550000000
0!
0%
#646555000000
1!
1%
#646560000000
0!
0%
#646565000000
1!
1%
#646570000000
0!
0%
#646575000000
1!
1%
#646580000000
0!
0%
#646585000000
1!
1%
#646590000000
0!
0%
#646595000000
1!
1%
#646600000000
0!
0%
#646605000000
1!
1%
#646610000000
0!
0%
#646615000000
1!
1%
#646620000000
0!
0%
#646625000000
1!
1%
#646630000000
0!
0%
#646635000000
1!
1%
#646640000000
0!
0%
#646645000000
1!
1%
#646650000000
0!
0%
#646655000000
1!
1%
#646660000000
0!
0%
#646665000000
1!
1%
#646670000000
0!
0%
#646675000000
1!
1%
#646680000000
0!
0%
#646685000000
1!
1%
#646690000000
0!
0%
#646695000000
1!
1%
#646700000000
0!
0%
#646705000000
1!
1%
#646710000000
0!
0%
#646715000000
1!
1%
#646720000000
0!
0%
#646725000000
1!
1%
#646730000000
0!
0%
#646735000000
1!
1%
#646740000000
0!
0%
#646745000000
1!
1%
#646750000000
0!
0%
#646755000000
1!
1%
#646760000000
0!
0%
#646765000000
1!
1%
#646770000000
0!
0%
#646775000000
1!
1%
#646780000000
0!
0%
#646785000000
1!
1%
#646790000000
0!
0%
#646795000000
1!
1%
#646800000000
0!
0%
#646805000000
1!
1%
#646810000000
0!
0%
#646815000000
1!
1%
#646820000000
0!
0%
#646825000000
1!
1%
#646830000000
0!
0%
#646835000000
1!
1%
#646840000000
0!
0%
#646845000000
1!
1%
#646850000000
0!
0%
#646855000000
1!
1%
#646860000000
0!
0%
#646865000000
1!
1%
#646870000000
0!
0%
#646875000000
1!
1%
#646880000000
0!
0%
#646885000000
1!
1%
#646890000000
0!
0%
#646895000000
1!
1%
#646900000000
0!
0%
#646905000000
1!
1%
#646910000000
0!
0%
#646915000000
1!
1%
#646920000000
0!
0%
#646925000000
1!
1%
#646930000000
0!
0%
#646935000000
1!
1%
#646940000000
0!
0%
#646945000000
1!
1%
#646950000000
0!
0%
#646955000000
1!
1%
#646960000000
0!
0%
#646965000000
1!
1%
#646970000000
0!
0%
#646975000000
1!
1%
#646980000000
0!
0%
#646985000000
1!
1%
#646990000000
0!
0%
#646995000000
1!
1%
#647000000000
0!
0%
#647005000000
1!
1%
#647010000000
0!
0%
#647015000000
1!
1%
#647020000000
0!
0%
#647025000000
1!
1%
#647030000000
0!
0%
#647035000000
1!
1%
#647040000000
0!
0%
#647045000000
1!
1%
#647050000000
0!
0%
#647055000000
1!
1%
#647060000000
0!
0%
#647065000000
1!
1%
#647070000000
0!
0%
#647075000000
1!
1%
#647080000000
0!
0%
#647085000000
1!
1%
#647090000000
0!
0%
#647095000000
1!
1%
#647100000000
0!
0%
#647105000000
1!
1%
#647110000000
0!
0%
#647115000000
1!
1%
#647120000000
0!
0%
#647125000000
1!
1%
#647130000000
0!
0%
#647135000000
1!
1%
#647140000000
0!
0%
#647145000000
1!
1%
#647150000000
0!
0%
#647155000000
1!
1%
#647160000000
0!
0%
#647165000000
1!
1%
#647170000000
0!
0%
#647175000000
1!
1%
#647180000000
0!
0%
#647185000000
1!
1%
#647190000000
0!
0%
#647195000000
1!
1%
#647200000000
0!
0%
#647205000000
1!
1%
#647210000000
0!
0%
#647215000000
1!
1%
#647220000000
0!
0%
#647225000000
1!
1%
#647230000000
0!
0%
#647235000000
1!
1%
#647240000000
0!
0%
#647245000000
1!
1%
#647250000000
0!
0%
#647255000000
1!
1%
#647260000000
0!
0%
#647265000000
1!
1%
#647270000000
0!
0%
#647275000000
1!
1%
#647280000000
0!
0%
#647285000000
1!
1%
#647290000000
0!
0%
#647295000000
1!
1%
#647300000000
0!
0%
#647305000000
1!
1%
#647310000000
0!
0%
#647315000000
1!
1%
#647320000000
0!
0%
#647325000000
1!
1%
#647330000000
0!
0%
#647335000000
1!
1%
#647340000000
0!
0%
#647345000000
1!
1%
#647350000000
0!
0%
#647355000000
1!
1%
#647360000000
0!
0%
#647365000000
1!
1%
#647370000000
0!
0%
#647375000000
1!
1%
#647380000000
0!
0%
#647385000000
1!
1%
#647390000000
0!
0%
#647395000000
1!
1%
#647400000000
0!
0%
#647405000000
1!
1%
#647410000000
0!
0%
#647415000000
1!
1%
#647420000000
0!
0%
#647425000000
1!
1%
#647430000000
0!
0%
#647435000000
1!
1%
#647440000000
0!
0%
#647445000000
1!
1%
#647450000000
0!
0%
#647455000000
1!
1%
#647460000000
0!
0%
#647465000000
1!
1%
#647470000000
0!
0%
#647475000000
1!
1%
#647480000000
0!
0%
#647485000000
1!
1%
#647490000000
0!
0%
#647495000000
1!
1%
#647500000000
0!
0%
#647505000000
1!
1%
#647510000000
0!
0%
#647515000000
1!
1%
#647520000000
0!
0%
#647525000000
1!
1%
#647530000000
0!
0%
#647535000000
1!
1%
#647540000000
0!
0%
#647545000000
1!
1%
#647550000000
0!
0%
#647555000000
1!
1%
#647560000000
0!
0%
#647565000000
1!
1%
#647570000000
0!
0%
#647575000000
1!
1%
#647580000000
0!
0%
#647585000000
1!
1%
#647590000000
0!
0%
#647595000000
1!
1%
#647600000000
0!
0%
#647605000000
1!
1%
#647610000000
0!
0%
#647615000000
1!
1%
#647620000000
0!
0%
#647625000000
1!
1%
#647630000000
0!
0%
#647635000000
1!
1%
#647640000000
0!
0%
#647645000000
1!
1%
#647650000000
0!
0%
#647655000000
1!
1%
#647660000000
0!
0%
#647665000000
1!
1%
#647670000000
0!
0%
#647675000000
1!
1%
#647680000000
0!
0%
#647685000000
1!
1%
#647690000000
0!
0%
#647695000000
1!
1%
#647700000000
0!
0%
#647705000000
1!
1%
#647710000000
0!
0%
#647715000000
1!
1%
#647720000000
0!
0%
#647725000000
1!
1%
#647730000000
0!
0%
#647735000000
1!
1%
#647740000000
0!
0%
#647745000000
1!
1%
#647750000000
0!
0%
#647755000000
1!
1%
#647760000000
0!
0%
#647765000000
1!
1%
#647770000000
0!
0%
#647775000000
1!
1%
#647780000000
0!
0%
#647785000000
1!
1%
#647790000000
0!
0%
#647795000000
1!
1%
#647800000000
0!
0%
#647805000000
1!
1%
#647810000000
0!
0%
#647815000000
1!
1%
#647820000000
0!
0%
#647825000000
1!
1%
#647830000000
0!
0%
#647835000000
1!
1%
#647840000000
0!
0%
#647845000000
1!
1%
#647850000000
0!
0%
#647855000000
1!
1%
#647860000000
0!
0%
#647865000000
1!
1%
#647870000000
0!
0%
#647875000000
1!
1%
#647880000000
0!
0%
#647885000000
1!
1%
#647890000000
0!
0%
#647895000000
1!
1%
#647900000000
0!
0%
#647905000000
1!
1%
#647910000000
0!
0%
#647915000000
1!
1%
#647920000000
0!
0%
#647925000000
1!
1%
#647930000000
0!
0%
#647935000000
1!
1%
#647940000000
0!
0%
#647945000000
1!
1%
#647950000000
0!
0%
#647955000000
1!
1%
#647960000000
0!
0%
#647965000000
1!
1%
#647970000000
0!
0%
#647975000000
1!
1%
#647980000000
0!
0%
#647985000000
1!
1%
#647990000000
0!
0%
#647995000000
1!
1%
#648000000000
0!
0%
#648005000000
1!
1%
#648010000000
0!
0%
#648015000000
1!
1%
#648020000000
0!
0%
#648025000000
1!
1%
#648030000000
0!
0%
#648035000000
1!
1%
#648040000000
0!
0%
#648045000000
1!
1%
#648050000000
0!
0%
#648055000000
1!
1%
#648060000000
0!
0%
#648065000000
1!
1%
#648070000000
0!
0%
#648075000000
1!
1%
#648080000000
0!
0%
#648085000000
1!
1%
#648090000000
0!
0%
#648095000000
1!
1%
#648100000000
0!
0%
#648105000000
1!
1%
#648110000000
0!
0%
#648115000000
1!
1%
#648120000000
0!
0%
#648125000000
1!
1%
#648130000000
0!
0%
#648135000000
1!
1%
#648140000000
0!
0%
#648145000000
1!
1%
#648150000000
0!
0%
#648155000000
1!
1%
#648160000000
0!
0%
#648165000000
1!
1%
#648170000000
0!
0%
#648175000000
1!
1%
#648180000000
0!
0%
#648185000000
1!
1%
#648190000000
0!
0%
#648195000000
1!
1%
#648200000000
0!
0%
#648205000000
1!
1%
#648210000000
0!
0%
#648215000000
1!
1%
#648220000000
0!
0%
#648225000000
1!
1%
#648230000000
0!
0%
#648235000000
1!
1%
#648240000000
0!
0%
#648245000000
1!
1%
#648250000000
0!
0%
#648255000000
1!
1%
#648260000000
0!
0%
#648265000000
1!
1%
#648270000000
0!
0%
#648275000000
1!
1%
#648280000000
0!
0%
#648285000000
1!
1%
#648290000000
0!
0%
#648295000000
1!
1%
#648300000000
0!
0%
#648305000000
1!
1%
#648310000000
0!
0%
#648315000000
1!
1%
#648320000000
0!
0%
#648325000000
1!
1%
#648330000000
0!
0%
#648335000000
1!
1%
#648340000000
0!
0%
#648345000000
1!
1%
#648350000000
0!
0%
#648355000000
1!
1%
#648360000000
0!
0%
#648365000000
1!
1%
#648370000000
0!
0%
#648375000000
1!
1%
#648380000000
0!
0%
#648385000000
1!
1%
#648390000000
0!
0%
#648395000000
1!
1%
#648400000000
0!
0%
#648405000000
1!
1%
#648410000000
0!
0%
#648415000000
1!
1%
#648420000000
0!
0%
#648425000000
1!
1%
#648430000000
0!
0%
#648435000000
1!
1%
#648440000000
0!
0%
#648445000000
1!
1%
#648450000000
0!
0%
#648455000000
1!
1%
#648460000000
0!
0%
#648465000000
1!
1%
#648470000000
0!
0%
#648475000000
1!
1%
#648480000000
0!
0%
#648485000000
1!
1%
#648490000000
0!
0%
#648495000000
1!
1%
#648500000000
0!
0%
#648505000000
1!
1%
#648510000000
0!
0%
#648515000000
1!
1%
#648520000000
0!
0%
#648525000000
1!
1%
#648530000000
0!
0%
#648535000000
1!
1%
#648540000000
0!
0%
#648545000000
1!
1%
#648550000000
0!
0%
#648555000000
1!
1%
#648560000000
0!
0%
#648565000000
1!
1%
#648570000000
0!
0%
#648575000000
1!
1%
#648580000000
0!
0%
#648585000000
1!
1%
#648590000000
0!
0%
#648595000000
1!
1%
#648600000000
0!
0%
#648605000000
1!
1%
#648610000000
0!
0%
#648615000000
1!
1%
#648620000000
0!
0%
#648625000000
1!
1%
#648630000000
0!
0%
#648635000000
1!
1%
#648640000000
0!
0%
#648645000000
1!
1%
#648650000000
0!
0%
#648655000000
1!
1%
#648660000000
0!
0%
#648665000000
1!
1%
#648670000000
0!
0%
#648675000000
1!
1%
#648680000000
0!
0%
#648685000000
1!
1%
#648690000000
0!
0%
#648695000000
1!
1%
#648700000000
0!
0%
#648705000000
1!
1%
#648710000000
0!
0%
#648715000000
1!
1%
#648720000000
0!
0%
#648725000000
1!
1%
#648730000000
0!
0%
#648735000000
1!
1%
#648740000000
0!
0%
#648745000000
1!
1%
#648750000000
0!
0%
#648755000000
1!
1%
#648760000000
0!
0%
#648765000000
1!
1%
#648770000000
0!
0%
#648775000000
1!
1%
#648780000000
0!
0%
#648785000000
1!
1%
#648790000000
0!
0%
#648795000000
1!
1%
#648800000000
0!
0%
#648805000000
1!
1%
#648810000000
0!
0%
#648815000000
1!
1%
#648820000000
0!
0%
#648825000000
1!
1%
#648830000000
0!
0%
#648835000000
1!
1%
#648840000000
0!
0%
#648845000000
1!
1%
#648850000000
0!
0%
#648855000000
1!
1%
#648860000000
0!
0%
#648865000000
1!
1%
#648870000000
0!
0%
#648875000000
1!
1%
#648880000000
0!
0%
#648885000000
1!
1%
#648890000000
0!
0%
#648895000000
1!
1%
#648900000000
0!
0%
#648905000000
1!
1%
#648910000000
0!
0%
#648915000000
1!
1%
#648920000000
0!
0%
#648925000000
1!
1%
#648930000000
0!
0%
#648935000000
1!
1%
#648940000000
0!
0%
#648945000000
1!
1%
#648950000000
0!
0%
#648955000000
1!
1%
#648960000000
0!
0%
#648965000000
1!
1%
#648970000000
0!
0%
#648975000000
1!
1%
#648980000000
0!
0%
#648985000000
1!
1%
#648990000000
0!
0%
#648995000000
1!
1%
#649000000000
0!
0%
#649005000000
1!
1%
#649010000000
0!
0%
#649015000000
1!
1%
#649020000000
0!
0%
#649025000000
1!
1%
#649030000000
0!
0%
#649035000000
1!
1%
#649040000000
0!
0%
#649045000000
1!
1%
#649050000000
0!
0%
#649055000000
1!
1%
#649060000000
0!
0%
#649065000000
1!
1%
#649070000000
0!
0%
#649075000000
1!
1%
#649080000000
0!
0%
#649085000000
1!
1%
#649090000000
0!
0%
#649095000000
1!
1%
#649100000000
0!
0%
#649105000000
1!
1%
#649110000000
0!
0%
#649115000000
1!
1%
#649120000000
0!
0%
#649125000000
1!
1%
#649130000000
0!
0%
#649135000000
1!
1%
#649140000000
0!
0%
#649145000000
1!
1%
#649150000000
0!
0%
#649155000000
1!
1%
#649160000000
0!
0%
#649165000000
1!
1%
#649170000000
0!
0%
#649175000000
1!
1%
#649180000000
0!
0%
#649185000000
1!
1%
#649190000000
0!
0%
#649195000000
1!
1%
#649200000000
0!
0%
#649205000000
1!
1%
#649210000000
0!
0%
#649215000000
1!
1%
#649220000000
0!
0%
#649225000000
1!
1%
#649230000000
0!
0%
#649235000000
1!
1%
#649240000000
0!
0%
#649245000000
1!
1%
#649250000000
0!
0%
#649255000000
1!
1%
#649260000000
0!
0%
#649265000000
1!
1%
#649270000000
0!
0%
#649275000000
1!
1%
#649280000000
0!
0%
#649285000000
1!
1%
#649290000000
0!
0%
#649295000000
1!
1%
#649300000000
0!
0%
#649305000000
1!
1%
#649310000000
0!
0%
#649315000000
1!
1%
#649320000000
0!
0%
#649325000000
1!
1%
#649330000000
0!
0%
#649335000000
1!
1%
#649340000000
0!
0%
#649345000000
1!
1%
#649350000000
0!
0%
#649355000000
1!
1%
#649360000000
0!
0%
#649365000000
1!
1%
#649370000000
0!
0%
#649375000000
1!
1%
#649380000000
0!
0%
#649385000000
1!
1%
#649390000000
0!
0%
#649395000000
1!
1%
#649400000000
0!
0%
#649405000000
1!
1%
#649410000000
0!
0%
#649415000000
1!
1%
#649420000000
0!
0%
#649425000000
1!
1%
#649430000000
0!
0%
#649435000000
1!
1%
#649440000000
0!
0%
#649445000000
1!
1%
#649450000000
0!
0%
#649455000000
1!
1%
#649460000000
0!
0%
#649465000000
1!
1%
#649470000000
0!
0%
#649475000000
1!
1%
#649480000000
0!
0%
#649485000000
1!
1%
#649490000000
0!
0%
#649495000000
1!
1%
#649500000000
0!
0%
#649505000000
1!
1%
#649510000000
0!
0%
#649515000000
1!
1%
#649520000000
0!
0%
#649525000000
1!
1%
#649530000000
0!
0%
#649535000000
1!
1%
#649540000000
0!
0%
#649545000000
1!
1%
#649550000000
0!
0%
#649555000000
1!
1%
#649560000000
0!
0%
#649565000000
1!
1%
#649570000000
0!
0%
#649575000000
1!
1%
#649580000000
0!
0%
#649585000000
1!
1%
#649590000000
0!
0%
#649595000000
1!
1%
#649600000000
0!
0%
#649605000000
1!
1%
#649610000000
0!
0%
#649615000000
1!
1%
#649620000000
0!
0%
#649625000000
1!
1%
#649630000000
0!
0%
#649635000000
1!
1%
#649640000000
0!
0%
#649645000000
1!
1%
#649650000000
0!
0%
#649655000000
1!
1%
#649660000000
0!
0%
#649665000000
1!
1%
#649670000000
0!
0%
#649675000000
1!
1%
#649680000000
0!
0%
#649685000000
1!
1%
#649690000000
0!
0%
#649695000000
1!
1%
#649700000000
0!
0%
#649705000000
1!
1%
#649710000000
0!
0%
#649715000000
1!
1%
#649720000000
0!
0%
#649725000000
1!
1%
#649730000000
0!
0%
#649735000000
1!
1%
#649740000000
0!
0%
#649745000000
1!
1%
#649750000000
0!
0%
#649755000000
1!
1%
#649760000000
0!
0%
#649765000000
1!
1%
#649770000000
0!
0%
#649775000000
1!
1%
#649780000000
0!
0%
#649785000000
1!
1%
#649790000000
0!
0%
#649795000000
1!
1%
#649800000000
0!
0%
#649805000000
1!
1%
#649810000000
0!
0%
#649815000000
1!
1%
#649820000000
0!
0%
#649825000000
1!
1%
#649830000000
0!
0%
#649835000000
1!
1%
#649840000000
0!
0%
#649845000000
1!
1%
#649850000000
0!
0%
#649855000000
1!
1%
#649860000000
0!
0%
#649865000000
1!
1%
#649870000000
0!
0%
#649875000000
1!
1%
#649880000000
0!
0%
#649885000000
1!
1%
#649890000000
0!
0%
#649895000000
1!
1%
#649900000000
0!
0%
#649905000000
1!
1%
#649910000000
0!
0%
#649915000000
1!
1%
#649920000000
0!
0%
#649925000000
1!
1%
#649930000000
0!
0%
#649935000000
1!
1%
#649940000000
0!
0%
#649945000000
1!
1%
#649950000000
0!
0%
#649955000000
1!
1%
#649960000000
0!
0%
#649965000000
1!
1%
#649970000000
0!
0%
#649975000000
1!
1%
#649980000000
0!
0%
#649985000000
1!
1%
#649990000000
0!
0%
#649995000000
1!
1%
#650000000000
0!
0%
#650005000000
1!
1%
#650010000000
0!
0%
#650015000000
1!
1%
#650020000000
0!
0%
#650025000000
1!
1%
#650030000000
0!
0%
#650035000000
1!
1%
#650040000000
0!
0%
#650045000000
1!
1%
#650050000000
0!
0%
#650055000000
1!
1%
#650060000000
0!
0%
#650065000000
1!
1%
#650070000000
0!
0%
#650075000000
1!
1%
#650080000000
0!
0%
#650085000000
1!
1%
#650090000000
0!
0%
#650095000000
1!
1%
#650100000000
0!
0%
#650105000000
1!
1%
#650110000000
0!
0%
#650115000000
1!
1%
#650120000000
0!
0%
#650125000000
1!
1%
#650130000000
0!
0%
#650135000000
1!
1%
#650140000000
0!
0%
#650145000000
1!
1%
#650150000000
0!
0%
#650155000000
1!
1%
#650160000000
0!
0%
#650165000000
1!
1%
#650170000000
0!
0%
#650175000000
1!
1%
#650180000000
0!
0%
#650185000000
1!
1%
#650190000000
0!
0%
#650195000000
1!
1%
#650200000000
0!
0%
#650205000000
1!
1%
#650210000000
0!
0%
#650215000000
1!
1%
#650220000000
0!
0%
#650225000000
1!
1%
#650230000000
0!
0%
#650235000000
1!
1%
#650240000000
0!
0%
#650245000000
1!
1%
#650250000000
0!
0%
#650255000000
1!
1%
#650260000000
0!
0%
#650265000000
1!
1%
#650270000000
0!
0%
#650275000000
1!
1%
#650280000000
0!
0%
#650285000000
1!
1%
#650290000000
0!
0%
#650295000000
1!
1%
#650300000000
0!
0%
#650305000000
1!
1%
#650310000000
0!
0%
#650315000000
1!
1%
#650320000000
0!
0%
#650325000000
1!
1%
#650330000000
0!
0%
#650335000000
1!
1%
#650340000000
0!
0%
#650345000000
1!
1%
#650350000000
0!
0%
#650355000000
1!
1%
#650360000000
0!
0%
#650365000000
1!
1%
#650370000000
0!
0%
#650375000000
1!
1%
#650380000000
0!
0%
#650385000000
1!
1%
#650390000000
0!
0%
#650395000000
1!
1%
#650400000000
0!
0%
#650405000000
1!
1%
#650410000000
0!
0%
#650415000000
1!
1%
#650420000000
0!
0%
#650425000000
1!
1%
#650430000000
0!
0%
#650435000000
1!
1%
#650440000000
0!
0%
#650445000000
1!
1%
#650450000000
0!
0%
#650455000000
1!
1%
#650460000000
0!
0%
#650465000000
1!
1%
#650470000000
0!
0%
#650475000000
1!
1%
#650480000000
0!
0%
#650485000000
1!
1%
#650490000000
0!
0%
#650495000000
1!
1%
#650500000000
0!
0%
#650505000000
1!
1%
#650510000000
0!
0%
#650515000000
1!
1%
#650520000000
0!
0%
#650525000000
1!
1%
#650530000000
0!
0%
#650535000000
1!
1%
#650540000000
0!
0%
#650545000000
1!
1%
#650550000000
0!
0%
#650555000000
1!
1%
#650560000000
0!
0%
#650565000000
1!
1%
#650570000000
0!
0%
#650575000000
1!
1%
#650580000000
0!
0%
#650585000000
1!
1%
#650590000000
0!
0%
#650595000000
1!
1%
#650600000000
0!
0%
#650605000000
1!
1%
#650610000000
0!
0%
#650615000000
1!
1%
#650620000000
0!
0%
#650625000000
1!
1%
#650630000000
0!
0%
#650635000000
1!
1%
#650640000000
0!
0%
#650645000000
1!
1%
#650650000000
0!
0%
#650655000000
1!
1%
#650660000000
0!
0%
#650665000000
1!
1%
#650670000000
0!
0%
#650675000000
1!
1%
#650680000000
0!
0%
#650685000000
1!
1%
#650690000000
0!
0%
#650695000000
1!
1%
#650700000000
0!
0%
#650705000000
1!
1%
#650710000000
0!
0%
#650715000000
1!
1%
#650720000000
0!
0%
#650725000000
1!
1%
#650730000000
0!
0%
#650735000000
1!
1%
#650740000000
0!
0%
#650745000000
1!
1%
#650750000000
0!
0%
#650755000000
1!
1%
#650760000000
0!
0%
#650765000000
1!
1%
#650770000000
0!
0%
#650775000000
1!
1%
#650780000000
0!
0%
#650785000000
1!
1%
#650790000000
0!
0%
#650795000000
1!
1%
#650800000000
0!
0%
#650805000000
1!
1%
#650810000000
0!
0%
#650815000000
1!
1%
#650820000000
0!
0%
#650825000000
1!
1%
#650830000000
0!
0%
#650835000000
1!
1%
#650840000000
0!
0%
#650845000000
1!
1%
#650850000000
0!
0%
#650855000000
1!
1%
#650860000000
0!
0%
#650865000000
1!
1%
#650870000000
0!
0%
#650875000000
1!
1%
#650880000000
0!
0%
#650885000000
1!
1%
#650890000000
0!
0%
#650895000000
1!
1%
#650900000000
0!
0%
#650905000000
1!
1%
#650910000000
0!
0%
#650915000000
1!
1%
#650920000000
0!
0%
#650925000000
1!
1%
#650930000000
0!
0%
#650935000000
1!
1%
#650940000000
0!
0%
#650945000000
1!
1%
#650950000000
0!
0%
#650955000000
1!
1%
#650960000000
0!
0%
#650965000000
1!
1%
#650970000000
0!
0%
#650975000000
1!
1%
#650980000000
0!
0%
#650985000000
1!
1%
#650990000000
0!
0%
#650995000000
1!
1%
#651000000000
0!
0%
#651005000000
1!
1%
#651010000000
0!
0%
#651015000000
1!
1%
#651020000000
0!
0%
#651025000000
1!
1%
#651030000000
0!
0%
#651035000000
1!
1%
#651040000000
0!
0%
#651045000000
1!
1%
#651050000000
0!
0%
#651055000000
1!
1%
#651060000000
0!
0%
#651065000000
1!
1%
#651070000000
0!
0%
#651075000000
1!
1%
#651080000000
0!
0%
#651085000000
1!
1%
#651090000000
0!
0%
#651095000000
1!
1%
#651100000000
0!
0%
#651105000000
1!
1%
#651110000000
0!
0%
#651115000000
1!
1%
#651120000000
0!
0%
#651125000000
1!
1%
#651130000000
0!
0%
#651135000000
1!
1%
#651140000000
0!
0%
#651145000000
1!
1%
#651150000000
0!
0%
#651155000000
1!
1%
#651160000000
0!
0%
#651165000000
1!
1%
#651170000000
0!
0%
#651175000000
1!
1%
#651180000000
0!
0%
#651185000000
1!
1%
#651190000000
0!
0%
#651195000000
1!
1%
#651200000000
0!
0%
#651205000000
1!
1%
#651210000000
0!
0%
#651215000000
1!
1%
#651220000000
0!
0%
#651225000000
1!
1%
#651230000000
0!
0%
#651235000000
1!
1%
#651240000000
0!
0%
#651245000000
1!
1%
#651250000000
0!
0%
#651255000000
1!
1%
#651260000000
0!
0%
#651265000000
1!
1%
#651270000000
0!
0%
#651275000000
1!
1%
#651280000000
0!
0%
#651285000000
1!
1%
#651290000000
0!
0%
#651295000000
1!
1%
#651300000000
0!
0%
#651305000000
1!
1%
#651310000000
0!
0%
#651315000000
1!
1%
#651320000000
0!
0%
#651325000000
1!
1%
#651330000000
0!
0%
#651335000000
1!
1%
#651340000000
0!
0%
#651345000000
1!
1%
#651350000000
0!
0%
#651355000000
1!
1%
#651360000000
0!
0%
#651365000000
1!
1%
#651370000000
0!
0%
#651375000000
1!
1%
#651380000000
0!
0%
#651385000000
1!
1%
#651390000000
0!
0%
#651395000000
1!
1%
#651400000000
0!
0%
#651405000000
1!
1%
#651410000000
0!
0%
#651415000000
1!
1%
#651420000000
0!
0%
#651425000000
1!
1%
#651430000000
0!
0%
#651435000000
1!
1%
#651440000000
0!
0%
#651445000000
1!
1%
#651450000000
0!
0%
#651455000000
1!
1%
#651460000000
0!
0%
#651465000000
1!
1%
#651470000000
0!
0%
#651475000000
1!
1%
#651480000000
0!
0%
#651485000000
1!
1%
#651490000000
0!
0%
#651495000000
1!
1%
#651500000000
0!
0%
#651505000000
1!
1%
#651510000000
0!
0%
#651515000000
1!
1%
#651520000000
0!
0%
#651525000000
1!
1%
#651530000000
0!
0%
#651535000000
1!
1%
#651540000000
0!
0%
#651545000000
1!
1%
#651550000000
0!
0%
#651555000000
1!
1%
#651560000000
0!
0%
#651565000000
1!
1%
#651570000000
0!
0%
#651575000000
1!
1%
#651580000000
0!
0%
#651585000000
1!
1%
#651590000000
0!
0%
#651595000000
1!
1%
#651600000000
0!
0%
#651605000000
1!
1%
#651610000000
0!
0%
#651615000000
1!
1%
#651620000000
0!
0%
#651625000000
1!
1%
#651630000000
0!
0%
#651635000000
1!
1%
#651640000000
0!
0%
#651645000000
1!
1%
#651650000000
0!
0%
#651655000000
1!
1%
#651660000000
0!
0%
#651665000000
1!
1%
#651670000000
0!
0%
#651675000000
1!
1%
#651680000000
0!
0%
#651685000000
1!
1%
#651690000000
0!
0%
#651695000000
1!
1%
#651700000000
0!
0%
#651705000000
1!
1%
#651710000000
0!
0%
#651715000000
1!
1%
#651720000000
0!
0%
#651725000000
1!
1%
#651730000000
0!
0%
#651735000000
1!
1%
#651740000000
0!
0%
#651745000000
1!
1%
#651750000000
0!
0%
#651755000000
1!
1%
#651760000000
0!
0%
#651765000000
1!
1%
#651770000000
0!
0%
#651775000000
1!
1%
#651780000000
0!
0%
#651785000000
1!
1%
#651790000000
0!
0%
#651795000000
1!
1%
#651800000000
0!
0%
#651805000000
1!
1%
#651810000000
0!
0%
#651815000000
1!
1%
#651820000000
0!
0%
#651825000000
1!
1%
#651830000000
0!
0%
#651835000000
1!
1%
#651840000000
0!
0%
#651845000000
1!
1%
#651850000000
0!
0%
#651855000000
1!
1%
#651860000000
0!
0%
#651865000000
1!
1%
#651870000000
0!
0%
#651875000000
1!
1%
#651880000000
0!
0%
#651885000000
1!
1%
#651890000000
0!
0%
#651895000000
1!
1%
#651900000000
0!
0%
#651905000000
1!
1%
#651910000000
0!
0%
#651915000000
1!
1%
#651920000000
0!
0%
#651925000000
1!
1%
#651930000000
0!
0%
#651935000000
1!
1%
#651940000000
0!
0%
#651945000000
1!
1%
#651950000000
0!
0%
#651955000000
1!
1%
#651960000000
0!
0%
#651965000000
1!
1%
#651970000000
0!
0%
#651975000000
1!
1%
#651980000000
0!
0%
#651985000000
1!
1%
#651990000000
0!
0%
#651995000000
1!
1%
#652000000000
0!
0%
#652005000000
1!
1%
#652010000000
0!
0%
#652015000000
1!
1%
#652020000000
0!
0%
#652025000000
1!
1%
#652030000000
0!
0%
#652035000000
1!
1%
#652040000000
0!
0%
#652045000000
1!
1%
#652050000000
0!
0%
#652055000000
1!
1%
#652060000000
0!
0%
#652065000000
1!
1%
#652070000000
0!
0%
#652075000000
1!
1%
#652080000000
0!
0%
#652085000000
1!
1%
#652090000000
0!
0%
#652095000000
1!
1%
#652100000000
0!
0%
#652105000000
1!
1%
#652110000000
0!
0%
#652115000000
1!
1%
#652120000000
0!
0%
#652125000000
1!
1%
#652130000000
0!
0%
#652135000000
1!
1%
#652140000000
0!
0%
#652145000000
1!
1%
#652150000000
0!
0%
#652155000000
1!
1%
#652160000000
0!
0%
#652165000000
1!
1%
#652170000000
0!
0%
#652175000000
1!
1%
#652180000000
0!
0%
#652185000000
1!
1%
#652190000000
0!
0%
#652195000000
1!
1%
#652200000000
0!
0%
#652205000000
1!
1%
#652210000000
0!
0%
#652215000000
1!
1%
#652220000000
0!
0%
#652225000000
1!
1%
#652230000000
0!
0%
#652235000000
1!
1%
#652240000000
0!
0%
#652245000000
1!
1%
#652250000000
0!
0%
#652255000000
1!
1%
#652260000000
0!
0%
#652265000000
1!
1%
#652270000000
0!
0%
#652275000000
1!
1%
#652280000000
0!
0%
#652285000000
1!
1%
#652290000000
0!
0%
#652295000000
1!
1%
#652300000000
0!
0%
#652305000000
1!
1%
#652310000000
0!
0%
#652315000000
1!
1%
#652320000000
0!
0%
#652325000000
1!
1%
#652330000000
0!
0%
#652335000000
1!
1%
#652340000000
0!
0%
#652345000000
1!
1%
#652350000000
0!
0%
#652355000000
1!
1%
#652360000000
0!
0%
#652365000000
1!
1%
#652370000000
0!
0%
#652375000000
1!
1%
#652380000000
0!
0%
#652385000000
1!
1%
#652390000000
0!
0%
#652395000000
1!
1%
#652400000000
0!
0%
#652405000000
1!
1%
#652410000000
0!
0%
#652415000000
1!
1%
#652420000000
0!
0%
#652425000000
1!
1%
#652430000000
0!
0%
#652435000000
1!
1%
#652440000000
0!
0%
#652445000000
1!
1%
#652450000000
0!
0%
#652455000000
1!
1%
#652460000000
0!
0%
#652465000000
1!
1%
#652470000000
0!
0%
#652475000000
1!
1%
#652480000000
0!
0%
#652485000000
1!
1%
#652490000000
0!
0%
#652495000000
1!
1%
#652500000000
0!
0%
#652505000000
1!
1%
#652510000000
0!
0%
#652515000000
1!
1%
#652520000000
0!
0%
#652525000000
1!
1%
#652530000000
0!
0%
#652535000000
1!
1%
#652540000000
0!
0%
#652545000000
1!
1%
#652550000000
0!
0%
#652555000000
1!
1%
#652560000000
0!
0%
#652565000000
1!
1%
#652570000000
0!
0%
#652575000000
1!
1%
#652580000000
0!
0%
#652585000000
1!
1%
#652590000000
0!
0%
#652595000000
1!
1%
#652600000000
0!
0%
#652605000000
1!
1%
#652610000000
0!
0%
#652615000000
1!
1%
#652620000000
0!
0%
#652625000000
1!
1%
#652630000000
0!
0%
#652635000000
1!
1%
#652640000000
0!
0%
#652645000000
1!
1%
#652650000000
0!
0%
#652655000000
1!
1%
#652660000000
0!
0%
#652665000000
1!
1%
#652670000000
0!
0%
#652675000000
1!
1%
#652680000000
0!
0%
#652685000000
1!
1%
#652690000000
0!
0%
#652695000000
1!
1%
#652700000000
0!
0%
#652705000000
1!
1%
#652710000000
0!
0%
#652715000000
1!
1%
#652720000000
0!
0%
#652725000000
1!
1%
#652730000000
0!
0%
#652735000000
1!
1%
#652740000000
0!
0%
#652745000000
1!
1%
#652750000000
0!
0%
#652755000000
1!
1%
#652760000000
0!
0%
#652765000000
1!
1%
#652770000000
0!
0%
#652775000000
1!
1%
#652780000000
0!
0%
#652785000000
1!
1%
#652790000000
0!
0%
#652795000000
1!
1%
#652800000000
0!
0%
#652805000000
1!
1%
#652810000000
0!
0%
#652815000000
1!
1%
#652820000000
0!
0%
#652825000000
1!
1%
#652830000000
0!
0%
#652835000000
1!
1%
#652840000000
0!
0%
#652845000000
1!
1%
#652850000000
0!
0%
#652855000000
1!
1%
#652860000000
0!
0%
#652865000000
1!
1%
#652870000000
0!
0%
#652875000000
1!
1%
#652880000000
0!
0%
#652885000000
1!
1%
#652890000000
0!
0%
#652895000000
1!
1%
#652900000000
0!
0%
#652905000000
1!
1%
#652910000000
0!
0%
#652915000000
1!
1%
#652920000000
0!
0%
#652925000000
1!
1%
#652930000000
0!
0%
#652935000000
1!
1%
#652940000000
0!
0%
#652945000000
1!
1%
#652950000000
0!
0%
#652955000000
1!
1%
#652960000000
0!
0%
#652965000000
1!
1%
#652970000000
0!
0%
#652975000000
1!
1%
#652980000000
0!
0%
#652985000000
1!
1%
#652990000000
0!
0%
#652995000000
1!
1%
#653000000000
0!
0%
#653005000000
1!
1%
#653010000000
0!
0%
#653015000000
1!
1%
#653020000000
0!
0%
#653025000000
1!
1%
#653030000000
0!
0%
#653035000000
1!
1%
#653040000000
0!
0%
#653045000000
1!
1%
#653050000000
0!
0%
#653055000000
1!
1%
#653060000000
0!
0%
#653065000000
1!
1%
#653070000000
0!
0%
#653075000000
1!
1%
#653080000000
0!
0%
#653085000000
1!
1%
#653090000000
0!
0%
#653095000000
1!
1%
#653100000000
0!
0%
#653105000000
1!
1%
#653110000000
0!
0%
#653115000000
1!
1%
#653120000000
0!
0%
#653125000000
1!
1%
#653130000000
0!
0%
#653135000000
1!
1%
#653140000000
0!
0%
#653145000000
1!
1%
#653150000000
0!
0%
#653155000000
1!
1%
#653160000000
0!
0%
#653165000000
1!
1%
#653170000000
0!
0%
#653175000000
1!
1%
#653180000000
0!
0%
#653185000000
1!
1%
#653190000000
0!
0%
#653195000000
1!
1%
#653200000000
0!
0%
#653205000000
1!
1%
#653210000000
0!
0%
#653215000000
1!
1%
#653220000000
0!
0%
#653225000000
1!
1%
#653230000000
0!
0%
#653235000000
1!
1%
#653240000000
0!
0%
#653245000000
1!
1%
#653250000000
0!
0%
#653255000000
1!
1%
#653260000000
0!
0%
#653265000000
1!
1%
#653270000000
0!
0%
#653275000000
1!
1%
#653280000000
0!
0%
#653285000000
1!
1%
#653290000000
0!
0%
#653295000000
1!
1%
#653300000000
0!
0%
#653305000000
1!
1%
#653310000000
0!
0%
#653315000000
1!
1%
#653320000000
0!
0%
#653325000000
1!
1%
#653330000000
0!
0%
#653335000000
1!
1%
#653340000000
0!
0%
#653345000000
1!
1%
#653350000000
0!
0%
#653355000000
1!
1%
#653360000000
0!
0%
#653365000000
1!
1%
#653370000000
0!
0%
#653375000000
1!
1%
#653380000000
0!
0%
#653385000000
1!
1%
#653390000000
0!
0%
#653395000000
1!
1%
#653400000000
0!
0%
#653405000000
1!
1%
#653410000000
0!
0%
#653415000000
1!
1%
#653420000000
0!
0%
#653425000000
1!
1%
#653430000000
0!
0%
#653435000000
1!
1%
#653440000000
0!
0%
#653445000000
1!
1%
#653450000000
0!
0%
#653455000000
1!
1%
#653460000000
0!
0%
#653465000000
1!
1%
#653470000000
0!
0%
#653475000000
1!
1%
#653480000000
0!
0%
#653485000000
1!
1%
#653490000000
0!
0%
#653495000000
1!
1%
#653500000000
0!
0%
#653505000000
1!
1%
#653510000000
0!
0%
#653515000000
1!
1%
#653520000000
0!
0%
#653525000000
1!
1%
#653530000000
0!
0%
#653535000000
1!
1%
#653540000000
0!
0%
#653545000000
1!
1%
#653550000000
0!
0%
#653555000000
1!
1%
#653560000000
0!
0%
#653565000000
1!
1%
#653570000000
0!
0%
#653575000000
1!
1%
#653580000000
0!
0%
#653585000000
1!
1%
#653590000000
0!
0%
#653595000000
1!
1%
#653600000000
0!
0%
#653605000000
1!
1%
#653610000000
0!
0%
#653615000000
1!
1%
#653620000000
0!
0%
#653625000000
1!
1%
#653630000000
0!
0%
#653635000000
1!
1%
#653640000000
0!
0%
#653645000000
1!
1%
#653650000000
0!
0%
#653655000000
1!
1%
#653660000000
0!
0%
#653665000000
1!
1%
#653670000000
0!
0%
#653675000000
1!
1%
#653680000000
0!
0%
#653685000000
1!
1%
#653690000000
0!
0%
#653695000000
1!
1%
#653700000000
0!
0%
#653705000000
1!
1%
#653710000000
0!
0%
#653715000000
1!
1%
#653720000000
0!
0%
#653725000000
1!
1%
#653730000000
0!
0%
#653735000000
1!
1%
#653740000000
0!
0%
#653745000000
1!
1%
#653750000000
0!
0%
#653755000000
1!
1%
#653760000000
0!
0%
#653765000000
1!
1%
#653770000000
0!
0%
#653775000000
1!
1%
#653780000000
0!
0%
#653785000000
1!
1%
#653790000000
0!
0%
#653795000000
1!
1%
#653800000000
0!
0%
#653805000000
1!
1%
#653810000000
0!
0%
#653815000000
1!
1%
#653820000000
0!
0%
#653825000000
1!
1%
#653830000000
0!
0%
#653835000000
1!
1%
#653840000000
0!
0%
#653845000000
1!
1%
#653850000000
0!
0%
#653855000000
1!
1%
#653860000000
0!
0%
#653865000000
1!
1%
#653870000000
0!
0%
#653875000000
1!
1%
#653880000000
0!
0%
#653885000000
1!
1%
#653890000000
0!
0%
#653895000000
1!
1%
#653900000000
0!
0%
#653905000000
1!
1%
#653910000000
0!
0%
#653915000000
1!
1%
#653920000000
0!
0%
#653925000000
1!
1%
#653930000000
0!
0%
#653935000000
1!
1%
#653940000000
0!
0%
#653945000000
1!
1%
#653950000000
0!
0%
#653955000000
1!
1%
#653960000000
0!
0%
#653965000000
1!
1%
#653970000000
0!
0%
#653975000000
1!
1%
#653980000000
0!
0%
#653985000000
1!
1%
#653990000000
0!
0%
#653995000000
1!
1%
#654000000000
0!
0%
#654005000000
1!
1%
#654010000000
0!
0%
#654015000000
1!
1%
#654020000000
0!
0%
#654025000000
1!
1%
#654030000000
0!
0%
#654035000000
1!
1%
#654040000000
0!
0%
#654045000000
1!
1%
#654050000000
0!
0%
#654055000000
1!
1%
#654060000000
0!
0%
#654065000000
1!
1%
#654070000000
0!
0%
#654075000000
1!
1%
#654080000000
0!
0%
#654085000000
1!
1%
#654090000000
0!
0%
#654095000000
1!
1%
#654100000000
0!
0%
#654105000000
1!
1%
#654110000000
0!
0%
#654115000000
1!
1%
#654120000000
0!
0%
#654125000000
1!
1%
#654130000000
0!
0%
#654135000000
1!
1%
#654140000000
0!
0%
#654145000000
1!
1%
#654150000000
0!
0%
#654155000000
1!
1%
#654160000000
0!
0%
#654165000000
1!
1%
#654170000000
0!
0%
#654175000000
1!
1%
#654180000000
0!
0%
#654185000000
1!
1%
#654190000000
0!
0%
#654195000000
1!
1%
#654200000000
0!
0%
#654205000000
1!
1%
#654210000000
0!
0%
#654215000000
1!
1%
#654220000000
0!
0%
#654225000000
1!
1%
#654230000000
0!
0%
#654235000000
1!
1%
#654240000000
0!
0%
#654245000000
1!
1%
#654250000000
0!
0%
#654255000000
1!
1%
#654260000000
0!
0%
#654265000000
1!
1%
#654270000000
0!
0%
#654275000000
1!
1%
#654280000000
0!
0%
#654285000000
1!
1%
#654290000000
0!
0%
#654295000000
1!
1%
#654300000000
0!
0%
#654305000000
1!
1%
#654310000000
0!
0%
#654315000000
1!
1%
#654320000000
0!
0%
#654325000000
1!
1%
#654330000000
0!
0%
#654335000000
1!
1%
#654340000000
0!
0%
#654345000000
1!
1%
#654350000000
0!
0%
#654355000000
1!
1%
#654360000000
0!
0%
#654365000000
1!
1%
#654370000000
0!
0%
#654375000000
1!
1%
#654380000000
0!
0%
#654385000000
1!
1%
#654390000000
0!
0%
#654395000000
1!
1%
#654400000000
0!
0%
#654405000000
1!
1%
#654410000000
0!
0%
#654415000000
1!
1%
#654420000000
0!
0%
#654425000000
1!
1%
#654430000000
0!
0%
#654435000000
1!
1%
#654440000000
0!
0%
#654445000000
1!
1%
#654450000000
0!
0%
#654455000000
1!
1%
#654460000000
0!
0%
#654465000000
1!
1%
#654470000000
0!
0%
#654475000000
1!
1%
#654480000000
0!
0%
#654485000000
1!
1%
#654490000000
0!
0%
#654495000000
1!
1%
#654500000000
0!
0%
#654505000000
1!
1%
#654510000000
0!
0%
#654515000000
1!
1%
#654520000000
0!
0%
#654525000000
1!
1%
#654530000000
0!
0%
#654535000000
1!
1%
#654540000000
0!
0%
#654545000000
1!
1%
#654550000000
0!
0%
#654555000000
1!
1%
#654560000000
0!
0%
#654565000000
1!
1%
#654570000000
0!
0%
#654575000000
1!
1%
#654580000000
0!
0%
#654585000000
1!
1%
#654590000000
0!
0%
#654595000000
1!
1%
#654600000000
0!
0%
#654605000000
1!
1%
#654610000000
0!
0%
#654615000000
1!
1%
#654620000000
0!
0%
#654625000000
1!
1%
#654630000000
0!
0%
#654635000000
1!
1%
#654640000000
0!
0%
#654645000000
1!
1%
#654650000000
0!
0%
#654655000000
1!
1%
#654660000000
0!
0%
#654665000000
1!
1%
#654670000000
0!
0%
#654675000000
1!
1%
#654680000000
0!
0%
#654685000000
1!
1%
#654690000000
0!
0%
#654695000000
1!
1%
#654700000000
0!
0%
#654705000000
1!
1%
#654710000000
0!
0%
#654715000000
1!
1%
#654720000000
0!
0%
#654725000000
1!
1%
#654730000000
0!
0%
#654735000000
1!
1%
#654740000000
0!
0%
#654745000000
1!
1%
#654750000000
0!
0%
#654755000000
1!
1%
#654760000000
0!
0%
#654765000000
1!
1%
#654770000000
0!
0%
#654775000000
1!
1%
#654780000000
0!
0%
#654785000000
1!
1%
#654790000000
0!
0%
#654795000000
1!
1%
#654800000000
0!
0%
#654805000000
1!
1%
#654810000000
0!
0%
#654815000000
1!
1%
#654820000000
0!
0%
#654825000000
1!
1%
#654830000000
0!
0%
#654835000000
1!
1%
#654840000000
0!
0%
#654845000000
1!
1%
#654850000000
0!
0%
#654855000000
1!
1%
#654860000000
0!
0%
#654865000000
1!
1%
#654870000000
0!
0%
#654875000000
1!
1%
#654880000000
0!
0%
#654885000000
1!
1%
#654890000000
0!
0%
#654895000000
1!
1%
#654900000000
0!
0%
#654905000000
1!
1%
#654910000000
0!
0%
#654915000000
1!
1%
#654920000000
0!
0%
#654925000000
1!
1%
#654930000000
0!
0%
#654935000000
1!
1%
#654940000000
0!
0%
#654945000000
1!
1%
#654950000000
0!
0%
#654955000000
1!
1%
#654960000000
0!
0%
#654965000000
1!
1%
#654970000000
0!
0%
#654975000000
1!
1%
#654980000000
0!
0%
#654985000000
1!
1%
#654990000000
0!
0%
#654995000000
1!
1%
#655000000000
0!
0%
#655005000000
1!
1%
#655010000000
0!
0%
#655015000000
1!
1%
#655020000000
0!
0%
#655025000000
1!
1%
#655030000000
0!
0%
#655035000000
1!
1%
#655040000000
0!
0%
#655045000000
1!
1%
#655050000000
0!
0%
#655055000000
1!
1%
#655060000000
0!
0%
#655065000000
1!
1%
#655070000000
0!
0%
#655075000000
1!
1%
#655080000000
0!
0%
#655085000000
1!
1%
#655090000000
0!
0%
#655095000000
1!
1%
#655100000000
0!
0%
#655105000000
1!
1%
#655110000000
0!
0%
#655115000000
1!
1%
#655120000000
0!
0%
#655125000000
1!
1%
#655130000000
0!
0%
#655135000000
1!
1%
#655140000000
0!
0%
#655145000000
1!
1%
#655150000000
0!
0%
#655155000000
1!
1%
#655160000000
0!
0%
#655165000000
1!
1%
#655170000000
0!
0%
#655175000000
1!
1%
#655180000000
0!
0%
#655185000000
1!
1%
#655190000000
0!
0%
#655195000000
1!
1%
#655200000000
0!
0%
#655205000000
1!
1%
#655210000000
0!
0%
#655215000000
1!
1%
#655220000000
0!
0%
#655225000000
1!
1%
#655230000000
0!
0%
#655235000000
1!
1%
#655240000000
0!
0%
#655245000000
1!
1%
#655250000000
0!
0%
#655255000000
1!
1%
#655260000000
0!
0%
#655265000000
1!
1%
#655270000000
0!
0%
#655275000000
1!
1%
#655280000000
0!
0%
#655285000000
1!
1%
#655290000000
0!
0%
#655295000000
1!
1%
#655300000000
0!
0%
#655305000000
1!
1%
#655310000000
0!
0%
#655315000000
1!
1%
#655320000000
0!
0%
#655325000000
1!
1%
#655330000000
0!
0%
#655335000000
1!
1%
#655340000000
0!
0%
#655345000000
1!
1%
#655350000000
0!
0%
#655355000000
1!
1%
#655360000000
0!
0%
#655365000000
1!
1%
#655370000000
0!
0%
#655375000000
1!
1%
#655380000000
0!
0%
#655385000000
1!
1%
#655390000000
0!
0%
#655395000000
1!
1%
#655400000000
0!
0%
#655405000000
1!
1%
#655410000000
0!
0%
#655415000000
1!
1%
#655420000000
0!
0%
#655425000000
1!
1%
#655430000000
0!
0%
#655435000000
1!
1%
#655440000000
0!
0%
#655445000000
1!
1%
#655450000000
0!
0%
#655455000000
1!
1%
#655460000000
0!
0%
#655465000000
1!
1%
#655470000000
0!
0%
#655475000000
1!
1%
#655480000000
0!
0%
#655485000000
1!
1%
#655490000000
0!
0%
#655495000000
1!
1%
#655500000000
0!
0%
#655505000000
1!
1%
#655510000000
0!
0%
#655515000000
1!
1%
#655520000000
0!
0%
#655525000000
1!
1%
#655530000000
0!
0%
#655535000000
1!
1%
#655540000000
0!
0%
#655545000000
1!
1%
#655550000000
0!
0%
#655555000000
1!
1%
#655560000000
0!
0%
#655565000000
1!
1%
#655570000000
0!
0%
#655575000000
1!
1%
#655580000000
0!
0%
#655585000000
1!
1%
#655590000000
0!
0%
#655595000000
1!
1%
#655600000000
0!
0%
#655605000000
1!
1%
#655610000000
0!
0%
#655615000000
1!
1%
#655620000000
0!
0%
#655625000000
1!
1%
#655630000000
0!
0%
#655635000000
1!
1%
#655640000000
0!
0%
#655645000000
1!
1%
#655650000000
0!
0%
#655655000000
1!
1%
#655660000000
0!
0%
#655665000000
1!
1%
#655670000000
0!
0%
#655675000000
1!
1%
#655680000000
0!
0%
#655685000000
1!
1%
#655690000000
0!
0%
#655695000000
1!
1%
#655700000000
0!
0%
#655705000000
1!
1%
#655710000000
0!
0%
#655715000000
1!
1%
#655720000000
0!
0%
#655725000000
1!
1%
#655730000000
0!
0%
#655735000000
1!
1%
#655740000000
0!
0%
#655745000000
1!
1%
#655750000000
0!
0%
#655755000000
1!
1%
#655760000000
0!
0%
#655765000000
1!
1%
#655770000000
0!
0%
#655775000000
1!
1%
#655780000000
0!
0%
#655785000000
1!
1%
#655790000000
0!
0%
#655795000000
1!
1%
#655800000000
0!
0%
#655805000000
1!
1%
#655810000000
0!
0%
#655815000000
1!
1%
#655820000000
0!
0%
#655825000000
1!
1%
#655830000000
0!
0%
#655835000000
1!
1%
#655840000000
0!
0%
#655845000000
1!
1%
#655850000000
0!
0%
#655855000000
1!
1%
#655860000000
0!
0%
#655865000000
1!
1%
#655870000000
0!
0%
#655875000000
1!
1%
#655880000000
0!
0%
#655885000000
1!
1%
#655890000000
0!
0%
#655895000000
1!
1%
#655900000000
0!
0%
#655905000000
1!
1%
#655910000000
0!
0%
#655915000000
1!
1%
#655920000000
0!
0%
#655925000000
1!
1%
#655930000000
0!
0%
#655935000000
1!
1%
#655940000000
0!
0%
#655945000000
1!
1%
#655950000000
0!
0%
#655955000000
1!
1%
#655960000000
0!
0%
#655965000000
1!
1%
#655970000000
0!
0%
#655975000000
1!
1%
#655980000000
0!
0%
#655985000000
1!
1%
#655990000000
0!
0%
#655995000000
1!
1%
#656000000000
0!
0%
#656005000000
1!
1%
#656010000000
0!
0%
#656015000000
1!
1%
#656020000000
0!
0%
#656025000000
1!
1%
#656030000000
0!
0%
#656035000000
1!
1%
#656040000000
0!
0%
#656045000000
1!
1%
#656050000000
0!
0%
#656055000000
1!
1%
#656060000000
0!
0%
#656065000000
1!
1%
#656070000000
0!
0%
#656075000000
1!
1%
#656080000000
0!
0%
#656085000000
1!
1%
#656090000000
0!
0%
#656095000000
1!
1%
#656100000000
0!
0%
#656105000000
1!
1%
#656110000000
0!
0%
#656115000000
1!
1%
#656120000000
0!
0%
#656125000000
1!
1%
#656130000000
0!
0%
#656135000000
1!
1%
#656140000000
0!
0%
#656145000000
1!
1%
#656150000000
0!
0%
#656155000000
1!
1%
#656160000000
0!
0%
#656165000000
1!
1%
#656170000000
0!
0%
#656175000000
1!
1%
#656180000000
0!
0%
#656185000000
1!
1%
#656190000000
0!
0%
#656195000000
1!
1%
#656200000000
0!
0%
#656205000000
1!
1%
#656210000000
0!
0%
#656215000000
1!
1%
#656220000000
0!
0%
#656225000000
1!
1%
#656230000000
0!
0%
#656235000000
1!
1%
#656240000000
0!
0%
#656245000000
1!
1%
#656250000000
0!
0%
#656255000000
1!
1%
#656260000000
0!
0%
#656265000000
1!
1%
#656270000000
0!
0%
#656275000000
1!
1%
#656280000000
0!
0%
#656285000000
1!
1%
#656290000000
0!
0%
#656295000000
1!
1%
#656300000000
0!
0%
#656305000000
1!
1%
#656310000000
0!
0%
#656315000000
1!
1%
#656320000000
0!
0%
#656325000000
1!
1%
#656330000000
0!
0%
#656335000000
1!
1%
#656340000000
0!
0%
#656345000000
1!
1%
#656350000000
0!
0%
#656355000000
1!
1%
#656360000000
0!
0%
#656365000000
1!
1%
#656370000000
0!
0%
#656375000000
1!
1%
#656380000000
0!
0%
#656385000000
1!
1%
#656390000000
0!
0%
#656395000000
1!
1%
#656400000000
0!
0%
#656405000000
1!
1%
#656410000000
0!
0%
#656415000000
1!
1%
#656420000000
0!
0%
#656425000000
1!
1%
#656430000000
0!
0%
#656435000000
1!
1%
#656440000000
0!
0%
#656445000000
1!
1%
#656450000000
0!
0%
#656455000000
1!
1%
#656460000000
0!
0%
#656465000000
1!
1%
#656470000000
0!
0%
#656475000000
1!
1%
#656480000000
0!
0%
#656485000000
1!
1%
#656490000000
0!
0%
#656495000000
1!
1%
#656500000000
0!
0%
#656505000000
1!
1%
#656510000000
0!
0%
#656515000000
1!
1%
#656520000000
0!
0%
#656525000000
1!
1%
#656530000000
0!
0%
#656535000000
1!
1%
#656540000000
0!
0%
#656545000000
1!
1%
#656550000000
0!
0%
#656555000000
1!
1%
#656560000000
0!
0%
#656565000000
1!
1%
#656570000000
0!
0%
#656575000000
1!
1%
#656580000000
0!
0%
#656585000000
1!
1%
#656590000000
0!
0%
#656595000000
1!
1%
#656600000000
0!
0%
#656605000000
1!
1%
#656610000000
0!
0%
#656615000000
1!
1%
#656620000000
0!
0%
#656625000000
1!
1%
#656630000000
0!
0%
#656635000000
1!
1%
#656640000000
0!
0%
#656645000000
1!
1%
#656650000000
0!
0%
#656655000000
1!
1%
#656660000000
0!
0%
#656665000000
1!
1%
#656670000000
0!
0%
#656675000000
1!
1%
#656680000000
0!
0%
#656685000000
1!
1%
#656690000000
0!
0%
#656695000000
1!
1%
#656700000000
0!
0%
#656705000000
1!
1%
#656710000000
0!
0%
#656715000000
1!
1%
#656720000000
0!
0%
#656725000000
1!
1%
#656730000000
0!
0%
#656735000000
1!
1%
#656740000000
0!
0%
#656745000000
1!
1%
#656750000000
0!
0%
#656755000000
1!
1%
#656760000000
0!
0%
#656765000000
1!
1%
#656770000000
0!
0%
#656775000000
1!
1%
#656780000000
0!
0%
#656785000000
1!
1%
#656790000000
0!
0%
#656795000000
1!
1%
#656800000000
0!
0%
#656805000000
1!
1%
#656810000000
0!
0%
#656815000000
1!
1%
#656820000000
0!
0%
#656825000000
1!
1%
#656830000000
0!
0%
#656835000000
1!
1%
#656840000000
0!
0%
#656845000000
1!
1%
#656850000000
0!
0%
#656855000000
1!
1%
#656860000000
0!
0%
#656865000000
1!
1%
#656870000000
0!
0%
#656875000000
1!
1%
#656880000000
0!
0%
#656885000000
1!
1%
#656890000000
0!
0%
#656895000000
1!
1%
#656900000000
0!
0%
#656905000000
1!
1%
#656910000000
0!
0%
#656915000000
1!
1%
#656920000000
0!
0%
#656925000000
1!
1%
#656930000000
0!
0%
#656935000000
1!
1%
#656940000000
0!
0%
#656945000000
1!
1%
#656950000000
0!
0%
#656955000000
1!
1%
#656960000000
0!
0%
#656965000000
1!
1%
#656970000000
0!
0%
#656975000000
1!
1%
#656980000000
0!
0%
#656985000000
1!
1%
#656990000000
0!
0%
#656995000000
1!
1%
#657000000000
0!
0%
#657005000000
1!
1%
#657010000000
0!
0%
#657015000000
1!
1%
#657020000000
0!
0%
#657025000000
1!
1%
#657030000000
0!
0%
#657035000000
1!
1%
#657040000000
0!
0%
#657045000000
1!
1%
#657050000000
0!
0%
#657055000000
1!
1%
#657060000000
0!
0%
#657065000000
1!
1%
#657070000000
0!
0%
#657075000000
1!
1%
#657080000000
0!
0%
#657085000000
1!
1%
#657090000000
0!
0%
#657095000000
1!
1%
#657100000000
0!
0%
#657105000000
1!
1%
#657110000000
0!
0%
#657115000000
1!
1%
#657120000000
0!
0%
#657125000000
1!
1%
#657130000000
0!
0%
#657135000000
1!
1%
#657140000000
0!
0%
#657145000000
1!
1%
#657150000000
0!
0%
#657155000000
1!
1%
#657160000000
0!
0%
#657165000000
1!
1%
#657170000000
0!
0%
#657175000000
1!
1%
#657180000000
0!
0%
#657185000000
1!
1%
#657190000000
0!
0%
#657195000000
1!
1%
#657200000000
0!
0%
#657205000000
1!
1%
#657210000000
0!
0%
#657215000000
1!
1%
#657220000000
0!
0%
#657225000000
1!
1%
#657230000000
0!
0%
#657235000000
1!
1%
#657240000000
0!
0%
#657245000000
1!
1%
#657250000000
0!
0%
#657255000000
1!
1%
#657260000000
0!
0%
#657265000000
1!
1%
#657270000000
0!
0%
#657275000000
1!
1%
#657280000000
0!
0%
#657285000000
1!
1%
#657290000000
0!
0%
#657295000000
1!
1%
#657300000000
0!
0%
#657305000000
1!
1%
#657310000000
0!
0%
#657315000000
1!
1%
#657320000000
0!
0%
#657325000000
1!
1%
#657330000000
0!
0%
#657335000000
1!
1%
#657340000000
0!
0%
#657345000000
1!
1%
#657350000000
0!
0%
#657355000000
1!
1%
#657360000000
0!
0%
#657365000000
1!
1%
#657370000000
0!
0%
#657375000000
1!
1%
#657380000000
0!
0%
#657385000000
1!
1%
#657390000000
0!
0%
#657395000000
1!
1%
#657400000000
0!
0%
#657405000000
1!
1%
#657410000000
0!
0%
#657415000000
1!
1%
#657420000000
0!
0%
#657425000000
1!
1%
#657430000000
0!
0%
#657435000000
1!
1%
#657440000000
0!
0%
#657445000000
1!
1%
#657450000000
0!
0%
#657455000000
1!
1%
#657460000000
0!
0%
#657465000000
1!
1%
#657470000000
0!
0%
#657475000000
1!
1%
#657480000000
0!
0%
#657485000000
1!
1%
#657490000000
0!
0%
#657495000000
1!
1%
#657500000000
0!
0%
#657505000000
1!
1%
#657510000000
0!
0%
#657515000000
1!
1%
#657520000000
0!
0%
#657525000000
1!
1%
#657530000000
0!
0%
#657535000000
1!
1%
#657540000000
0!
0%
#657545000000
1!
1%
#657550000000
0!
0%
#657555000000
1!
1%
#657560000000
0!
0%
#657565000000
1!
1%
#657570000000
0!
0%
#657575000000
1!
1%
#657580000000
0!
0%
#657585000000
1!
1%
#657590000000
0!
0%
#657595000000
1!
1%
#657600000000
0!
0%
#657605000000
1!
1%
#657610000000
0!
0%
#657615000000
1!
1%
#657620000000
0!
0%
#657625000000
1!
1%
#657630000000
0!
0%
#657635000000
1!
1%
#657640000000
0!
0%
#657645000000
1!
1%
#657650000000
0!
0%
#657655000000
1!
1%
#657660000000
0!
0%
#657665000000
1!
1%
#657670000000
0!
0%
#657675000000
1!
1%
#657680000000
0!
0%
#657685000000
1!
1%
#657690000000
0!
0%
#657695000000
1!
1%
#657700000000
0!
0%
#657705000000
1!
1%
#657710000000
0!
0%
#657715000000
1!
1%
#657720000000
0!
0%
#657725000000
1!
1%
#657730000000
0!
0%
#657735000000
1!
1%
#657740000000
0!
0%
#657745000000
1!
1%
#657750000000
0!
0%
#657755000000
1!
1%
#657760000000
0!
0%
#657765000000
1!
1%
#657770000000
0!
0%
#657775000000
1!
1%
#657780000000
0!
0%
#657785000000
1!
1%
#657790000000
0!
0%
#657795000000
1!
1%
#657800000000
0!
0%
#657805000000
1!
1%
#657810000000
0!
0%
#657815000000
1!
1%
#657820000000
0!
0%
#657825000000
1!
1%
#657830000000
0!
0%
#657835000000
1!
1%
#657840000000
0!
0%
#657845000000
1!
1%
#657850000000
0!
0%
#657855000000
1!
1%
#657860000000
0!
0%
#657865000000
1!
1%
#657870000000
0!
0%
#657875000000
1!
1%
#657880000000
0!
0%
#657885000000
1!
1%
#657890000000
0!
0%
#657895000000
1!
1%
#657900000000
0!
0%
#657905000000
1!
1%
#657910000000
0!
0%
#657915000000
1!
1%
#657920000000
0!
0%
#657925000000
1!
1%
#657930000000
0!
0%
#657935000000
1!
1%
#657940000000
0!
0%
#657945000000
1!
1%
#657950000000
0!
0%
#657955000000
1!
1%
#657960000000
0!
0%
#657965000000
1!
1%
#657970000000
0!
0%
#657975000000
1!
1%
#657980000000
0!
0%
#657985000000
1!
1%
#657990000000
0!
0%
#657995000000
1!
1%
#658000000000
0!
0%
#658005000000
1!
1%
#658010000000
0!
0%
#658015000000
1!
1%
#658020000000
0!
0%
#658025000000
1!
1%
#658030000000
0!
0%
#658035000000
1!
1%
#658040000000
0!
0%
#658045000000
1!
1%
#658050000000
0!
0%
#658055000000
1!
1%
#658060000000
0!
0%
#658065000000
1!
1%
#658070000000
0!
0%
#658075000000
1!
1%
#658080000000
0!
0%
#658085000000
1!
1%
#658090000000
0!
0%
#658095000000
1!
1%
#658100000000
0!
0%
#658105000000
1!
1%
#658110000000
0!
0%
#658115000000
1!
1%
#658120000000
0!
0%
#658125000000
1!
1%
#658130000000
0!
0%
#658135000000
1!
1%
#658140000000
0!
0%
#658145000000
1!
1%
#658150000000
0!
0%
#658155000000
1!
1%
#658160000000
0!
0%
#658165000000
1!
1%
#658170000000
0!
0%
#658175000000
1!
1%
#658180000000
0!
0%
#658185000000
1!
1%
#658190000000
0!
0%
#658195000000
1!
1%
#658200000000
0!
0%
#658205000000
1!
1%
#658210000000
0!
0%
#658215000000
1!
1%
#658220000000
0!
0%
#658225000000
1!
1%
#658230000000
0!
0%
#658235000000
1!
1%
#658240000000
0!
0%
#658245000000
1!
1%
#658250000000
0!
0%
#658255000000
1!
1%
#658260000000
0!
0%
#658265000000
1!
1%
#658270000000
0!
0%
#658275000000
1!
1%
#658280000000
0!
0%
#658285000000
1!
1%
#658290000000
0!
0%
#658295000000
1!
1%
#658300000000
0!
0%
#658305000000
1!
1%
#658310000000
0!
0%
#658315000000
1!
1%
#658320000000
0!
0%
#658325000000
1!
1%
#658330000000
0!
0%
#658335000000
1!
1%
#658340000000
0!
0%
#658345000000
1!
1%
#658350000000
0!
0%
#658355000000
1!
1%
#658360000000
0!
0%
#658365000000
1!
1%
#658370000000
0!
0%
#658375000000
1!
1%
#658380000000
0!
0%
#658385000000
1!
1%
#658390000000
0!
0%
#658395000000
1!
1%
#658400000000
0!
0%
#658405000000
1!
1%
#658410000000
0!
0%
#658415000000
1!
1%
#658420000000
0!
0%
#658425000000
1!
1%
#658430000000
0!
0%
#658435000000
1!
1%
#658440000000
0!
0%
#658445000000
1!
1%
#658450000000
0!
0%
#658455000000
1!
1%
#658460000000
0!
0%
#658465000000
1!
1%
#658470000000
0!
0%
#658475000000
1!
1%
#658480000000
0!
0%
#658485000000
1!
1%
#658490000000
0!
0%
#658495000000
1!
1%
#658500000000
0!
0%
#658505000000
1!
1%
#658510000000
0!
0%
#658515000000
1!
1%
#658520000000
0!
0%
#658525000000
1!
1%
#658530000000
0!
0%
#658535000000
1!
1%
#658540000000
0!
0%
#658545000000
1!
1%
#658550000000
0!
0%
#658555000000
1!
1%
#658560000000
0!
0%
#658565000000
1!
1%
#658570000000
0!
0%
#658575000000
1!
1%
#658580000000
0!
0%
#658585000000
1!
1%
#658590000000
0!
0%
#658595000000
1!
1%
#658600000000
0!
0%
#658605000000
1!
1%
#658610000000
0!
0%
#658615000000
1!
1%
#658620000000
0!
0%
#658625000000
1!
1%
#658630000000
0!
0%
#658635000000
1!
1%
#658640000000
0!
0%
#658645000000
1!
1%
#658650000000
0!
0%
#658655000000
1!
1%
#658660000000
0!
0%
#658665000000
1!
1%
#658670000000
0!
0%
#658675000000
1!
1%
#658680000000
0!
0%
#658685000000
1!
1%
#658690000000
0!
0%
#658695000000
1!
1%
#658700000000
0!
0%
#658705000000
1!
1%
#658710000000
0!
0%
#658715000000
1!
1%
#658720000000
0!
0%
#658725000000
1!
1%
#658730000000
0!
0%
#658735000000
1!
1%
#658740000000
0!
0%
#658745000000
1!
1%
#658750000000
0!
0%
#658755000000
1!
1%
#658760000000
0!
0%
#658765000000
1!
1%
#658770000000
0!
0%
#658775000000
1!
1%
#658780000000
0!
0%
#658785000000
1!
1%
#658790000000
0!
0%
#658795000000
1!
1%
#658800000000
0!
0%
#658805000000
1!
1%
#658810000000
0!
0%
#658815000000
1!
1%
#658820000000
0!
0%
#658825000000
1!
1%
#658830000000
0!
0%
#658835000000
1!
1%
#658840000000
0!
0%
#658845000000
1!
1%
#658850000000
0!
0%
#658855000000
1!
1%
#658860000000
0!
0%
#658865000000
1!
1%
#658870000000
0!
0%
#658875000000
1!
1%
#658880000000
0!
0%
#658885000000
1!
1%
#658890000000
0!
0%
#658895000000
1!
1%
#658900000000
0!
0%
#658905000000
1!
1%
#658910000000
0!
0%
#658915000000
1!
1%
#658920000000
0!
0%
#658925000000
1!
1%
#658930000000
0!
0%
#658935000000
1!
1%
#658940000000
0!
0%
#658945000000
1!
1%
#658950000000
0!
0%
#658955000000
1!
1%
#658960000000
0!
0%
#658965000000
1!
1%
#658970000000
0!
0%
#658975000000
1!
1%
#658980000000
0!
0%
#658985000000
1!
1%
#658990000000
0!
0%
#658995000000
1!
1%
#659000000000
0!
0%
#659005000000
1!
1%
#659010000000
0!
0%
#659015000000
1!
1%
#659020000000
0!
0%
#659025000000
1!
1%
#659030000000
0!
0%
#659035000000
1!
1%
#659040000000
0!
0%
#659045000000
1!
1%
#659050000000
0!
0%
#659055000000
1!
1%
#659060000000
0!
0%
#659065000000
1!
1%
#659070000000
0!
0%
#659075000000
1!
1%
#659080000000
0!
0%
#659085000000
1!
1%
#659090000000
0!
0%
#659095000000
1!
1%
#659100000000
0!
0%
#659105000000
1!
1%
#659110000000
0!
0%
#659115000000
1!
1%
#659120000000
0!
0%
#659125000000
1!
1%
#659130000000
0!
0%
#659135000000
1!
1%
#659140000000
0!
0%
#659145000000
1!
1%
#659150000000
0!
0%
#659155000000
1!
1%
#659160000000
0!
0%
#659165000000
1!
1%
#659170000000
0!
0%
#659175000000
1!
1%
#659180000000
0!
0%
#659185000000
1!
1%
#659190000000
0!
0%
#659195000000
1!
1%
#659200000000
0!
0%
#659205000000
1!
1%
#659210000000
0!
0%
#659215000000
1!
1%
#659220000000
0!
0%
#659225000000
1!
1%
#659230000000
0!
0%
#659235000000
1!
1%
#659240000000
0!
0%
#659245000000
1!
1%
#659250000000
0!
0%
#659255000000
1!
1%
#659260000000
0!
0%
#659265000000
1!
1%
#659270000000
0!
0%
#659275000000
1!
1%
#659280000000
0!
0%
#659285000000
1!
1%
#659290000000
0!
0%
#659295000000
1!
1%
#659300000000
0!
0%
#659305000000
1!
1%
#659310000000
0!
0%
#659315000000
1!
1%
#659320000000
0!
0%
#659325000000
1!
1%
#659330000000
0!
0%
#659335000000
1!
1%
#659340000000
0!
0%
#659345000000
1!
1%
#659350000000
0!
0%
#659355000000
1!
1%
#659360000000
0!
0%
#659365000000
1!
1%
#659370000000
0!
0%
#659375000000
1!
1%
#659380000000
0!
0%
#659385000000
1!
1%
#659390000000
0!
0%
#659395000000
1!
1%
#659400000000
0!
0%
#659405000000
1!
1%
#659410000000
0!
0%
#659415000000
1!
1%
#659420000000
0!
0%
#659425000000
1!
1%
#659430000000
0!
0%
#659435000000
1!
1%
#659440000000
0!
0%
#659445000000
1!
1%
#659450000000
0!
0%
#659455000000
1!
1%
#659460000000
0!
0%
#659465000000
1!
1%
#659470000000
0!
0%
#659475000000
1!
1%
#659480000000
0!
0%
#659485000000
1!
1%
#659490000000
0!
0%
#659495000000
1!
1%
#659500000000
0!
0%
#659505000000
1!
1%
#659510000000
0!
0%
#659515000000
1!
1%
#659520000000
0!
0%
#659525000000
1!
1%
#659530000000
0!
0%
#659535000000
1!
1%
#659540000000
0!
0%
#659545000000
1!
1%
#659550000000
0!
0%
#659555000000
1!
1%
#659560000000
0!
0%
#659565000000
1!
1%
#659570000000
0!
0%
#659575000000
1!
1%
#659580000000
0!
0%
#659585000000
1!
1%
#659590000000
0!
0%
#659595000000
1!
1%
#659600000000
0!
0%
#659605000000
1!
1%
#659610000000
0!
0%
#659615000000
1!
1%
#659620000000
0!
0%
#659625000000
1!
1%
#659630000000
0!
0%
#659635000000
1!
1%
#659640000000
0!
0%
#659645000000
1!
1%
#659650000000
0!
0%
#659655000000
1!
1%
#659660000000
0!
0%
#659665000000
1!
1%
#659670000000
0!
0%
#659675000000
1!
1%
#659680000000
0!
0%
#659685000000
1!
1%
#659690000000
0!
0%
#659695000000
1!
1%
#659700000000
0!
0%
#659705000000
1!
1%
#659710000000
0!
0%
#659715000000
1!
1%
#659720000000
0!
0%
#659725000000
1!
1%
#659730000000
0!
0%
#659735000000
1!
1%
#659740000000
0!
0%
#659745000000
1!
1%
#659750000000
0!
0%
#659755000000
1!
1%
#659760000000
0!
0%
#659765000000
1!
1%
#659770000000
0!
0%
#659775000000
1!
1%
#659780000000
0!
0%
#659785000000
1!
1%
#659790000000
0!
0%
#659795000000
1!
1%
#659800000000
0!
0%
#659805000000
1!
1%
#659810000000
0!
0%
#659815000000
1!
1%
#659820000000
0!
0%
#659825000000
1!
1%
#659830000000
0!
0%
#659835000000
1!
1%
#659840000000
0!
0%
#659845000000
1!
1%
#659850000000
0!
0%
#659855000000
1!
1%
#659860000000
0!
0%
#659865000000
1!
1%
#659870000000
0!
0%
#659875000000
1!
1%
#659880000000
0!
0%
#659885000000
1!
1%
#659890000000
0!
0%
#659895000000
1!
1%
#659900000000
0!
0%
#659905000000
1!
1%
#659910000000
0!
0%
#659915000000
1!
1%
#659920000000
0!
0%
#659925000000
1!
1%
#659930000000
0!
0%
#659935000000
1!
1%
#659940000000
0!
0%
#659945000000
1!
1%
#659950000000
0!
0%
#659955000000
1!
1%
#659960000000
0!
0%
#659965000000
1!
1%
#659970000000
0!
0%
#659975000000
1!
1%
#659980000000
0!
0%
#659985000000
1!
1%
#659990000000
0!
0%
#659995000000
1!
1%
#660000000000
0!
0%
#660005000000
1!
1%
#660010000000
0!
0%
#660015000000
1!
1%
#660020000000
0!
0%
#660025000000
1!
1%
#660030000000
0!
0%
#660035000000
1!
1%
#660040000000
0!
0%
#660045000000
1!
1%
#660050000000
0!
0%
#660055000000
1!
1%
#660060000000
0!
0%
#660065000000
1!
1%
#660070000000
0!
0%
#660075000000
1!
1%
#660080000000
0!
0%
#660085000000
1!
1%
#660090000000
0!
0%
#660095000000
1!
1%
#660100000000
0!
0%
#660105000000
1!
1%
#660110000000
0!
0%
#660115000000
1!
1%
#660120000000
0!
0%
#660125000000
1!
1%
#660130000000
0!
0%
#660135000000
1!
1%
#660140000000
0!
0%
#660145000000
1!
1%
#660150000000
0!
0%
#660155000000
1!
1%
#660160000000
0!
0%
#660165000000
1!
1%
#660170000000
0!
0%
#660175000000
1!
1%
#660180000000
0!
0%
#660185000000
1!
1%
#660190000000
0!
0%
#660195000000
1!
1%
#660200000000
0!
0%
#660205000000
1!
1%
#660210000000
0!
0%
#660215000000
1!
1%
#660220000000
0!
0%
#660225000000
1!
1%
#660230000000
0!
0%
#660235000000
1!
1%
#660240000000
0!
0%
#660245000000
1!
1%
#660250000000
0!
0%
#660255000000
1!
1%
#660260000000
0!
0%
#660265000000
1!
1%
#660270000000
0!
0%
#660275000000
1!
1%
#660280000000
0!
0%
#660285000000
1!
1%
#660290000000
0!
0%
#660295000000
1!
1%
#660300000000
0!
0%
#660305000000
1!
1%
#660310000000
0!
0%
#660315000000
1!
1%
#660320000000
0!
0%
#660325000000
1!
1%
#660330000000
0!
0%
#660335000000
1!
1%
#660340000000
0!
0%
#660345000000
1!
1%
#660350000000
0!
0%
#660355000000
1!
1%
#660360000000
0!
0%
#660365000000
1!
1%
#660370000000
0!
0%
#660375000000
1!
1%
#660380000000
0!
0%
#660385000000
1!
1%
#660390000000
0!
0%
#660395000000
1!
1%
#660400000000
0!
0%
#660405000000
1!
1%
#660410000000
0!
0%
#660415000000
1!
1%
#660420000000
0!
0%
#660425000000
1!
1%
#660430000000
0!
0%
#660435000000
1!
1%
#660440000000
0!
0%
#660445000000
1!
1%
#660450000000
0!
0%
#660455000000
1!
1%
#660460000000
0!
0%
#660465000000
1!
1%
#660470000000
0!
0%
#660475000000
1!
1%
#660480000000
0!
0%
#660485000000
1!
1%
#660490000000
0!
0%
#660495000000
1!
1%
#660500000000
0!
0%
#660505000000
1!
1%
#660510000000
0!
0%
#660515000000
1!
1%
#660520000000
0!
0%
#660525000000
1!
1%
#660530000000
0!
0%
#660535000000
1!
1%
#660540000000
0!
0%
#660545000000
1!
1%
#660550000000
0!
0%
#660555000000
1!
1%
#660560000000
0!
0%
#660565000000
1!
1%
#660570000000
0!
0%
#660575000000
1!
1%
#660580000000
0!
0%
#660585000000
1!
1%
#660590000000
0!
0%
#660595000000
1!
1%
#660600000000
0!
0%
#660605000000
1!
1%
#660610000000
0!
0%
#660615000000
1!
1%
#660620000000
0!
0%
#660625000000
1!
1%
#660630000000
0!
0%
#660635000000
1!
1%
#660640000000
0!
0%
#660645000000
1!
1%
#660650000000
0!
0%
#660655000000
1!
1%
#660660000000
0!
0%
#660665000000
1!
1%
#660670000000
0!
0%
#660675000000
1!
1%
#660680000000
0!
0%
#660685000000
1!
1%
#660690000000
0!
0%
#660695000000
1!
1%
#660700000000
0!
0%
#660705000000
1!
1%
#660710000000
0!
0%
#660715000000
1!
1%
#660720000000
0!
0%
#660725000000
1!
1%
#660730000000
0!
0%
#660735000000
1!
1%
#660740000000
0!
0%
#660745000000
1!
1%
#660750000000
0!
0%
#660755000000
1!
1%
#660760000000
0!
0%
#660765000000
1!
1%
#660770000000
0!
0%
#660775000000
1!
1%
#660780000000
0!
0%
#660785000000
1!
1%
#660790000000
0!
0%
#660795000000
1!
1%
#660800000000
0!
0%
#660805000000
1!
1%
#660810000000
0!
0%
#660815000000
1!
1%
#660820000000
0!
0%
#660825000000
1!
1%
#660830000000
0!
0%
#660835000000
1!
1%
#660840000000
0!
0%
#660845000000
1!
1%
#660850000000
0!
0%
#660855000000
1!
1%
#660860000000
0!
0%
#660865000000
1!
1%
#660870000000
0!
0%
#660875000000
1!
1%
#660880000000
0!
0%
#660885000000
1!
1%
#660890000000
0!
0%
#660895000000
1!
1%
#660900000000
0!
0%
#660905000000
1!
1%
#660910000000
0!
0%
#660915000000
1!
1%
#660920000000
0!
0%
#660925000000
1!
1%
#660930000000
0!
0%
#660935000000
1!
1%
#660940000000
0!
0%
#660945000000
1!
1%
#660950000000
0!
0%
#660955000000
1!
1%
#660960000000
0!
0%
#660965000000
1!
1%
#660970000000
0!
0%
#660975000000
1!
1%
#660980000000
0!
0%
#660985000000
1!
1%
#660990000000
0!
0%
#660995000000
1!
1%
#661000000000
0!
0%
#661005000000
1!
1%
#661010000000
0!
0%
#661015000000
1!
1%
#661020000000
0!
0%
#661025000000
1!
1%
#661030000000
0!
0%
#661035000000
1!
1%
#661040000000
0!
0%
#661045000000
1!
1%
#661050000000
0!
0%
#661055000000
1!
1%
#661060000000
0!
0%
#661065000000
1!
1%
#661070000000
0!
0%
#661075000000
1!
1%
#661080000000
0!
0%
#661085000000
1!
1%
#661090000000
0!
0%
#661095000000
1!
1%
#661100000000
0!
0%
#661105000000
1!
1%
#661110000000
0!
0%
#661115000000
1!
1%
#661120000000
0!
0%
#661125000000
1!
1%
#661130000000
0!
0%
#661135000000
1!
1%
#661140000000
0!
0%
#661145000000
1!
1%
#661150000000
0!
0%
#661155000000
1!
1%
#661160000000
0!
0%
#661165000000
1!
1%
#661170000000
0!
0%
#661175000000
1!
1%
#661180000000
0!
0%
#661185000000
1!
1%
#661190000000
0!
0%
#661195000000
1!
1%
#661200000000
0!
0%
#661205000000
1!
1%
#661210000000
0!
0%
#661215000000
1!
1%
#661220000000
0!
0%
#661225000000
1!
1%
#661230000000
0!
0%
#661235000000
1!
1%
#661240000000
0!
0%
#661245000000
1!
1%
#661250000000
0!
0%
#661255000000
1!
1%
#661260000000
0!
0%
#661265000000
1!
1%
#661270000000
0!
0%
#661275000000
1!
1%
#661280000000
0!
0%
#661285000000
1!
1%
#661290000000
0!
0%
#661295000000
1!
1%
#661300000000
0!
0%
#661305000000
1!
1%
#661310000000
0!
0%
#661315000000
1!
1%
#661320000000
0!
0%
#661325000000
1!
1%
#661330000000
0!
0%
#661335000000
1!
1%
#661340000000
0!
0%
#661345000000
1!
1%
#661350000000
0!
0%
#661355000000
1!
1%
#661360000000
0!
0%
#661365000000
1!
1%
#661370000000
0!
0%
#661375000000
1!
1%
#661380000000
0!
0%
#661385000000
1!
1%
#661390000000
0!
0%
#661395000000
1!
1%
#661400000000
0!
0%
#661405000000
1!
1%
#661410000000
0!
0%
#661415000000
1!
1%
#661420000000
0!
0%
#661425000000
1!
1%
#661430000000
0!
0%
#661435000000
1!
1%
#661440000000
0!
0%
#661445000000
1!
1%
#661450000000
0!
0%
#661455000000
1!
1%
#661460000000
0!
0%
#661465000000
1!
1%
#661470000000
0!
0%
#661475000000
1!
1%
#661480000000
0!
0%
#661485000000
1!
1%
#661490000000
0!
0%
#661495000000
1!
1%
#661500000000
0!
0%
#661505000000
1!
1%
#661510000000
0!
0%
#661515000000
1!
1%
#661520000000
0!
0%
#661525000000
1!
1%
#661530000000
0!
0%
#661535000000
1!
1%
#661540000000
0!
0%
#661545000000
1!
1%
#661550000000
0!
0%
#661555000000
1!
1%
#661560000000
0!
0%
#661565000000
1!
1%
#661570000000
0!
0%
#661575000000
1!
1%
#661580000000
0!
0%
#661585000000
1!
1%
#661590000000
0!
0%
#661595000000
1!
1%
#661600000000
0!
0%
#661605000000
1!
1%
#661610000000
0!
0%
#661615000000
1!
1%
#661620000000
0!
0%
#661625000000
1!
1%
#661630000000
0!
0%
#661635000000
1!
1%
#661640000000
0!
0%
#661645000000
1!
1%
#661650000000
0!
0%
#661655000000
1!
1%
#661660000000
0!
0%
#661665000000
1!
1%
#661670000000
0!
0%
#661675000000
1!
1%
#661680000000
0!
0%
#661685000000
1!
1%
#661690000000
0!
0%
#661695000000
1!
1%
#661700000000
0!
0%
#661705000000
1!
1%
#661710000000
0!
0%
#661715000000
1!
1%
#661720000000
0!
0%
#661725000000
1!
1%
#661730000000
0!
0%
#661735000000
1!
1%
#661740000000
0!
0%
#661745000000
1!
1%
#661750000000
0!
0%
#661755000000
1!
1%
#661760000000
0!
0%
#661765000000
1!
1%
#661770000000
0!
0%
#661775000000
1!
1%
#661780000000
0!
0%
#661785000000
1!
1%
#661790000000
0!
0%
#661795000000
1!
1%
#661800000000
0!
0%
#661805000000
1!
1%
#661810000000
0!
0%
#661815000000
1!
1%
#661820000000
0!
0%
#661825000000
1!
1%
#661830000000
0!
0%
#661835000000
1!
1%
#661840000000
0!
0%
#661845000000
1!
1%
#661850000000
0!
0%
#661855000000
1!
1%
#661860000000
0!
0%
#661865000000
1!
1%
#661870000000
0!
0%
#661875000000
1!
1%
#661880000000
0!
0%
#661885000000
1!
1%
#661890000000
0!
0%
#661895000000
1!
1%
#661900000000
0!
0%
#661905000000
1!
1%
#661910000000
0!
0%
#661915000000
1!
1%
#661920000000
0!
0%
#661925000000
1!
1%
#661930000000
0!
0%
#661935000000
1!
1%
#661940000000
0!
0%
#661945000000
1!
1%
#661950000000
0!
0%
#661955000000
1!
1%
#661960000000
0!
0%
#661965000000
1!
1%
#661970000000
0!
0%
#661975000000
1!
1%
#661980000000
0!
0%
#661985000000
1!
1%
#661990000000
0!
0%
#661995000000
1!
1%
#662000000000
0!
0%
#662005000000
1!
1%
#662010000000
0!
0%
#662015000000
1!
1%
#662020000000
0!
0%
#662025000000
1!
1%
#662030000000
0!
0%
#662035000000
1!
1%
#662040000000
0!
0%
#662045000000
1!
1%
#662050000000
0!
0%
#662055000000
1!
1%
#662060000000
0!
0%
#662065000000
1!
1%
#662070000000
0!
0%
#662075000000
1!
1%
#662080000000
0!
0%
#662085000000
1!
1%
#662090000000
0!
0%
#662095000000
1!
1%
#662100000000
0!
0%
#662105000000
1!
1%
#662110000000
0!
0%
#662115000000
1!
1%
#662120000000
0!
0%
#662125000000
1!
1%
#662130000000
0!
0%
#662135000000
1!
1%
#662140000000
0!
0%
#662145000000
1!
1%
#662150000000
0!
0%
#662155000000
1!
1%
#662160000000
0!
0%
#662165000000
1!
1%
#662170000000
0!
0%
#662175000000
1!
1%
#662180000000
0!
0%
#662185000000
1!
1%
#662190000000
0!
0%
#662195000000
1!
1%
#662200000000
0!
0%
#662205000000
1!
1%
#662210000000
0!
0%
#662215000000
1!
1%
#662220000000
0!
0%
#662225000000
1!
1%
#662230000000
0!
0%
#662235000000
1!
1%
#662240000000
0!
0%
#662245000000
1!
1%
#662250000000
0!
0%
#662255000000
1!
1%
#662260000000
0!
0%
#662265000000
1!
1%
#662270000000
0!
0%
#662275000000
1!
1%
#662280000000
0!
0%
#662285000000
1!
1%
#662290000000
0!
0%
#662295000000
1!
1%
#662300000000
0!
0%
#662305000000
1!
1%
#662310000000
0!
0%
#662315000000
1!
1%
#662320000000
0!
0%
#662325000000
1!
1%
#662330000000
0!
0%
#662335000000
1!
1%
#662340000000
0!
0%
#662345000000
1!
1%
#662350000000
0!
0%
#662355000000
1!
1%
#662360000000
0!
0%
#662365000000
1!
1%
#662370000000
0!
0%
#662375000000
1!
1%
#662380000000
0!
0%
#662385000000
1!
1%
#662390000000
0!
0%
#662395000000
1!
1%
#662400000000
0!
0%
#662405000000
1!
1%
#662410000000
0!
0%
#662415000000
1!
1%
#662420000000
0!
0%
#662425000000
1!
1%
#662430000000
0!
0%
#662435000000
1!
1%
#662440000000
0!
0%
#662445000000
1!
1%
#662450000000
0!
0%
#662455000000
1!
1%
#662460000000
0!
0%
#662465000000
1!
1%
#662470000000
0!
0%
#662475000000
1!
1%
#662480000000
0!
0%
#662485000000
1!
1%
#662490000000
0!
0%
#662495000000
1!
1%
#662500000000
0!
0%
#662505000000
1!
1%
#662510000000
0!
0%
#662515000000
1!
1%
#662520000000
0!
0%
#662525000000
1!
1%
#662530000000
0!
0%
#662535000000
1!
1%
#662540000000
0!
0%
#662545000000
1!
1%
#662550000000
0!
0%
#662555000000
1!
1%
#662560000000
0!
0%
#662565000000
1!
1%
#662570000000
0!
0%
#662575000000
1!
1%
#662580000000
0!
0%
#662585000000
1!
1%
#662590000000
0!
0%
#662595000000
1!
1%
#662600000000
0!
0%
#662605000000
1!
1%
#662610000000
0!
0%
#662615000000
1!
1%
#662620000000
0!
0%
#662625000000
1!
1%
#662630000000
0!
0%
#662635000000
1!
1%
#662640000000
0!
0%
#662645000000
1!
1%
#662650000000
0!
0%
#662655000000
1!
1%
#662660000000
0!
0%
#662665000000
1!
1%
#662670000000
0!
0%
#662675000000
1!
1%
#662680000000
0!
0%
#662685000000
1!
1%
#662690000000
0!
0%
#662695000000
1!
1%
#662700000000
0!
0%
#662705000000
1!
1%
#662710000000
0!
0%
#662715000000
1!
1%
#662720000000
0!
0%
#662725000000
1!
1%
#662730000000
0!
0%
#662735000000
1!
1%
#662740000000
0!
0%
#662745000000
1!
1%
#662750000000
0!
0%
#662755000000
1!
1%
#662760000000
0!
0%
#662765000000
1!
1%
#662770000000
0!
0%
#662775000000
1!
1%
#662780000000
0!
0%
#662785000000
1!
1%
#662790000000
0!
0%
#662795000000
1!
1%
#662800000000
0!
0%
#662805000000
1!
1%
#662810000000
0!
0%
#662815000000
1!
1%
#662820000000
0!
0%
#662825000000
1!
1%
#662830000000
0!
0%
#662835000000
1!
1%
#662840000000
0!
0%
#662845000000
1!
1%
#662850000000
0!
0%
#662855000000
1!
1%
#662860000000
0!
0%
#662865000000
1!
1%
#662870000000
0!
0%
#662875000000
1!
1%
#662880000000
0!
0%
#662885000000
1!
1%
#662890000000
0!
0%
#662895000000
1!
1%
#662900000000
0!
0%
#662905000000
1!
1%
#662910000000
0!
0%
#662915000000
1!
1%
#662920000000
0!
0%
#662925000000
1!
1%
#662930000000
0!
0%
#662935000000
1!
1%
#662940000000
0!
0%
#662945000000
1!
1%
#662950000000
0!
0%
#662955000000
1!
1%
#662960000000
0!
0%
#662965000000
1!
1%
#662970000000
0!
0%
#662975000000
1!
1%
#662980000000
0!
0%
#662985000000
1!
1%
#662990000000
0!
0%
#662995000000
1!
1%
#663000000000
0!
0%
#663005000000
1!
1%
#663010000000
0!
0%
#663015000000
1!
1%
#663020000000
0!
0%
#663025000000
1!
1%
#663030000000
0!
0%
#663035000000
1!
1%
#663040000000
0!
0%
#663045000000
1!
1%
#663050000000
0!
0%
#663055000000
1!
1%
#663060000000
0!
0%
#663065000000
1!
1%
#663070000000
0!
0%
#663075000000
1!
1%
#663080000000
0!
0%
#663085000000
1!
1%
#663090000000
0!
0%
#663095000000
1!
1%
#663100000000
0!
0%
#663105000000
1!
1%
#663110000000
0!
0%
#663115000000
1!
1%
#663120000000
0!
0%
#663125000000
1!
1%
#663130000000
0!
0%
#663135000000
1!
1%
#663140000000
0!
0%
#663145000000
1!
1%
#663150000000
0!
0%
#663155000000
1!
1%
#663160000000
0!
0%
#663165000000
1!
1%
#663170000000
0!
0%
#663175000000
1!
1%
#663180000000
0!
0%
#663185000000
1!
1%
#663190000000
0!
0%
#663195000000
1!
1%
#663200000000
0!
0%
#663205000000
1!
1%
#663210000000
0!
0%
#663215000000
1!
1%
#663220000000
0!
0%
#663225000000
1!
1%
#663230000000
0!
0%
#663235000000
1!
1%
#663240000000
0!
0%
#663245000000
1!
1%
#663250000000
0!
0%
#663255000000
1!
1%
#663260000000
0!
0%
#663265000000
1!
1%
#663270000000
0!
0%
#663275000000
1!
1%
#663280000000
0!
0%
#663285000000
1!
1%
#663290000000
0!
0%
#663295000000
1!
1%
#663300000000
0!
0%
#663305000000
1!
1%
#663310000000
0!
0%
#663315000000
1!
1%
#663320000000
0!
0%
#663325000000
1!
1%
#663330000000
0!
0%
#663335000000
1!
1%
#663340000000
0!
0%
#663345000000
1!
1%
#663350000000
0!
0%
#663355000000
1!
1%
#663360000000
0!
0%
#663365000000
1!
1%
#663370000000
0!
0%
#663375000000
1!
1%
#663380000000
0!
0%
#663385000000
1!
1%
#663390000000
0!
0%
#663395000000
1!
1%
#663400000000
0!
0%
#663405000000
1!
1%
#663410000000
0!
0%
#663415000000
1!
1%
#663420000000
0!
0%
#663425000000
1!
1%
#663430000000
0!
0%
#663435000000
1!
1%
#663440000000
0!
0%
#663445000000
1!
1%
#663450000000
0!
0%
#663455000000
1!
1%
#663460000000
0!
0%
#663465000000
1!
1%
#663470000000
0!
0%
#663475000000
1!
1%
#663480000000
0!
0%
#663485000000
1!
1%
#663490000000
0!
0%
#663495000000
1!
1%
#663500000000
0!
0%
#663505000000
1!
1%
#663510000000
0!
0%
#663515000000
1!
1%
#663520000000
0!
0%
#663525000000
1!
1%
#663530000000
0!
0%
#663535000000
1!
1%
#663540000000
0!
0%
#663545000000
1!
1%
#663550000000
0!
0%
#663555000000
1!
1%
#663560000000
0!
0%
#663565000000
1!
1%
#663570000000
0!
0%
#663575000000
1!
1%
#663580000000
0!
0%
#663585000000
1!
1%
#663590000000
0!
0%
#663595000000
1!
1%
#663600000000
0!
0%
#663605000000
1!
1%
#663610000000
0!
0%
#663615000000
1!
1%
#663620000000
0!
0%
#663625000000
1!
1%
#663630000000
0!
0%
#663635000000
1!
1%
#663640000000
0!
0%
#663645000000
1!
1%
#663650000000
0!
0%
#663655000000
1!
1%
#663660000000
0!
0%
#663665000000
1!
1%
#663670000000
0!
0%
#663675000000
1!
1%
#663680000000
0!
0%
#663685000000
1!
1%
#663690000000
0!
0%
#663695000000
1!
1%
#663700000000
0!
0%
#663705000000
1!
1%
#663710000000
0!
0%
#663715000000
1!
1%
#663720000000
0!
0%
#663725000000
1!
1%
#663730000000
0!
0%
#663735000000
1!
1%
#663740000000
0!
0%
#663745000000
1!
1%
#663750000000
0!
0%
#663755000000
1!
1%
#663760000000
0!
0%
#663765000000
1!
1%
#663770000000
0!
0%
#663775000000
1!
1%
#663780000000
0!
0%
#663785000000
1!
1%
#663790000000
0!
0%
#663795000000
1!
1%
#663800000000
0!
0%
#663805000000
1!
1%
#663810000000
0!
0%
#663815000000
1!
1%
#663820000000
0!
0%
#663825000000
1!
1%
#663830000000
0!
0%
#663835000000
1!
1%
#663840000000
0!
0%
#663845000000
1!
1%
#663850000000
0!
0%
#663855000000
1!
1%
#663860000000
0!
0%
#663865000000
1!
1%
#663870000000
0!
0%
#663875000000
1!
1%
#663880000000
0!
0%
#663885000000
1!
1%
#663890000000
0!
0%
#663895000000
1!
1%
#663900000000
0!
0%
#663905000000
1!
1%
#663910000000
0!
0%
#663915000000
1!
1%
#663920000000
0!
0%
#663925000000
1!
1%
#663930000000
0!
0%
#663935000000
1!
1%
#663940000000
0!
0%
#663945000000
1!
1%
#663950000000
0!
0%
#663955000000
1!
1%
#663960000000
0!
0%
#663965000000
1!
1%
#663970000000
0!
0%
#663975000000
1!
1%
#663980000000
0!
0%
#663985000000
1!
1%
#663990000000
0!
0%
#663995000000
1!
1%
#664000000000
0!
0%
#664005000000
1!
1%
#664010000000
0!
0%
#664015000000
1!
1%
#664020000000
0!
0%
#664025000000
1!
1%
#664030000000
0!
0%
#664035000000
1!
1%
#664040000000
0!
0%
#664045000000
1!
1%
#664050000000
0!
0%
#664055000000
1!
1%
#664060000000
0!
0%
#664065000000
1!
1%
#664070000000
0!
0%
#664075000000
1!
1%
#664080000000
0!
0%
#664085000000
1!
1%
#664090000000
0!
0%
#664095000000
1!
1%
#664100000000
0!
0%
#664105000000
1!
1%
#664110000000
0!
0%
#664115000000
1!
1%
#664120000000
0!
0%
#664125000000
1!
1%
#664130000000
0!
0%
#664135000000
1!
1%
#664140000000
0!
0%
#664145000000
1!
1%
#664150000000
0!
0%
#664155000000
1!
1%
#664160000000
0!
0%
#664165000000
1!
1%
#664170000000
0!
0%
#664175000000
1!
1%
#664180000000
0!
0%
#664185000000
1!
1%
#664190000000
0!
0%
#664195000000
1!
1%
#664200000000
0!
0%
#664205000000
1!
1%
#664210000000
0!
0%
#664215000000
1!
1%
#664220000000
0!
0%
#664225000000
1!
1%
#664230000000
0!
0%
#664235000000
1!
1%
#664240000000
0!
0%
#664245000000
1!
1%
#664250000000
0!
0%
#664255000000
1!
1%
#664260000000
0!
0%
#664265000000
1!
1%
#664270000000
0!
0%
#664275000000
1!
1%
#664280000000
0!
0%
#664285000000
1!
1%
#664290000000
0!
0%
#664295000000
1!
1%
#664300000000
0!
0%
#664305000000
1!
1%
#664310000000
0!
0%
#664315000000
1!
1%
#664320000000
0!
0%
#664325000000
1!
1%
#664330000000
0!
0%
#664335000000
1!
1%
#664340000000
0!
0%
#664345000000
1!
1%
#664350000000
0!
0%
#664355000000
1!
1%
#664360000000
0!
0%
#664365000000
1!
1%
#664370000000
0!
0%
#664375000000
1!
1%
#664380000000
0!
0%
#664385000000
1!
1%
#664390000000
0!
0%
#664395000000
1!
1%
#664400000000
0!
0%
#664405000000
1!
1%
#664410000000
0!
0%
#664415000000
1!
1%
#664420000000
0!
0%
#664425000000
1!
1%
#664430000000
0!
0%
#664435000000
1!
1%
#664440000000
0!
0%
#664445000000
1!
1%
#664450000000
0!
0%
#664455000000
1!
1%
#664460000000
0!
0%
#664465000000
1!
1%
#664470000000
0!
0%
#664475000000
1!
1%
#664480000000
0!
0%
#664485000000
1!
1%
#664490000000
0!
0%
#664495000000
1!
1%
#664500000000
0!
0%
#664505000000
1!
1%
#664510000000
0!
0%
#664515000000
1!
1%
#664520000000
0!
0%
#664525000000
1!
1%
#664530000000
0!
0%
#664535000000
1!
1%
#664540000000
0!
0%
#664545000000
1!
1%
#664550000000
0!
0%
#664555000000
1!
1%
#664560000000
0!
0%
#664565000000
1!
1%
#664570000000
0!
0%
#664575000000
1!
1%
#664580000000
0!
0%
#664585000000
1!
1%
#664590000000
0!
0%
#664595000000
1!
1%
#664600000000
0!
0%
#664605000000
1!
1%
#664610000000
0!
0%
#664615000000
1!
1%
#664620000000
0!
0%
#664625000000
1!
1%
#664630000000
0!
0%
#664635000000
1!
1%
#664640000000
0!
0%
#664645000000
1!
1%
#664650000000
0!
0%
#664655000000
1!
1%
#664660000000
0!
0%
#664665000000
1!
1%
#664670000000
0!
0%
#664675000000
1!
1%
#664680000000
0!
0%
#664685000000
1!
1%
#664690000000
0!
0%
#664695000000
1!
1%
#664700000000
0!
0%
#664705000000
1!
1%
#664710000000
0!
0%
#664715000000
1!
1%
#664720000000
0!
0%
#664725000000
1!
1%
#664730000000
0!
0%
#664735000000
1!
1%
#664740000000
0!
0%
#664745000000
1!
1%
#664750000000
0!
0%
#664755000000
1!
1%
#664760000000
0!
0%
#664765000000
1!
1%
#664770000000
0!
0%
#664775000000
1!
1%
#664780000000
0!
0%
#664785000000
1!
1%
#664790000000
0!
0%
#664795000000
1!
1%
#664800000000
0!
0%
#664805000000
1!
1%
#664810000000
0!
0%
#664815000000
1!
1%
#664820000000
0!
0%
#664825000000
1!
1%
#664830000000
0!
0%
#664835000000
1!
1%
#664840000000
0!
0%
#664845000000
1!
1%
#664850000000
0!
0%
#664855000000
1!
1%
#664860000000
0!
0%
#664865000000
1!
1%
#664870000000
0!
0%
#664875000000
1!
1%
#664880000000
0!
0%
#664885000000
1!
1%
#664890000000
0!
0%
#664895000000
1!
1%
#664900000000
0!
0%
#664905000000
1!
1%
#664910000000
0!
0%
#664915000000
1!
1%
#664920000000
0!
0%
#664925000000
1!
1%
#664930000000
0!
0%
#664935000000
1!
1%
#664940000000
0!
0%
#664945000000
1!
1%
#664950000000
0!
0%
#664955000000
1!
1%
#664960000000
0!
0%
#664965000000
1!
1%
#664970000000
0!
0%
#664975000000
1!
1%
#664980000000
0!
0%
#664985000000
1!
1%
#664990000000
0!
0%
#664995000000
1!
1%
#665000000000
0!
0%
#665005000000
1!
1%
#665010000000
0!
0%
#665015000000
1!
1%
#665020000000
0!
0%
#665025000000
1!
1%
#665030000000
0!
0%
#665035000000
1!
1%
#665040000000
0!
0%
#665045000000
1!
1%
#665050000000
0!
0%
#665055000000
1!
1%
#665060000000
0!
0%
#665065000000
1!
1%
#665070000000
0!
0%
#665075000000
1!
1%
#665080000000
0!
0%
#665085000000
1!
1%
#665090000000
0!
0%
#665095000000
1!
1%
#665100000000
0!
0%
#665105000000
1!
1%
#665110000000
0!
0%
#665115000000
1!
1%
#665120000000
0!
0%
#665125000000
1!
1%
#665130000000
0!
0%
#665135000000
1!
1%
#665140000000
0!
0%
#665145000000
1!
1%
#665150000000
0!
0%
#665155000000
1!
1%
#665160000000
0!
0%
#665165000000
1!
1%
#665170000000
0!
0%
#665175000000
1!
1%
#665180000000
0!
0%
#665185000000
1!
1%
#665190000000
0!
0%
#665195000000
1!
1%
#665200000000
0!
0%
#665205000000
1!
1%
#665210000000
0!
0%
#665215000000
1!
1%
#665220000000
0!
0%
#665225000000
1!
1%
#665230000000
0!
0%
#665235000000
1!
1%
#665240000000
0!
0%
#665245000000
1!
1%
#665250000000
0!
0%
#665255000000
1!
1%
#665260000000
0!
0%
#665265000000
1!
1%
#665270000000
0!
0%
#665275000000
1!
1%
#665280000000
0!
0%
#665285000000
1!
1%
#665290000000
0!
0%
#665295000000
1!
1%
#665300000000
0!
0%
#665305000000
1!
1%
#665310000000
0!
0%
#665315000000
1!
1%
#665320000000
0!
0%
#665325000000
1!
1%
#665330000000
0!
0%
#665335000000
1!
1%
#665340000000
0!
0%
#665345000000
1!
1%
#665350000000
0!
0%
#665355000000
1!
1%
#665360000000
0!
0%
#665365000000
1!
1%
#665370000000
0!
0%
#665375000000
1!
1%
#665380000000
0!
0%
#665385000000
1!
1%
#665390000000
0!
0%
#665395000000
1!
1%
#665400000000
0!
0%
#665405000000
1!
1%
#665410000000
0!
0%
#665415000000
1!
1%
#665420000000
0!
0%
#665425000000
1!
1%
#665430000000
0!
0%
#665435000000
1!
1%
#665440000000
0!
0%
#665445000000
1!
1%
#665450000000
0!
0%
#665455000000
1!
1%
#665460000000
0!
0%
#665465000000
1!
1%
#665470000000
0!
0%
#665475000000
1!
1%
#665480000000
0!
0%
#665485000000
1!
1%
#665490000000
0!
0%
#665495000000
1!
1%
#665500000000
0!
0%
#665505000000
1!
1%
#665510000000
0!
0%
#665515000000
1!
1%
#665520000000
0!
0%
#665525000000
1!
1%
#665530000000
0!
0%
#665535000000
1!
1%
#665540000000
0!
0%
#665545000000
1!
1%
#665550000000
0!
0%
#665555000000
1!
1%
#665560000000
0!
0%
#665565000000
1!
1%
#665570000000
0!
0%
#665575000000
1!
1%
#665580000000
0!
0%
#665585000000
1!
1%
#665590000000
0!
0%
#665595000000
1!
1%
#665600000000
0!
0%
#665605000000
1!
1%
#665610000000
0!
0%
#665615000000
1!
1%
#665620000000
0!
0%
#665625000000
1!
1%
#665630000000
0!
0%
#665635000000
1!
1%
#665640000000
0!
0%
#665645000000
1!
1%
#665650000000
0!
0%
#665655000000
1!
1%
#665660000000
0!
0%
#665665000000
1!
1%
#665670000000
0!
0%
#665675000000
1!
1%
#665680000000
0!
0%
#665685000000
1!
1%
#665690000000
0!
0%
#665695000000
1!
1%
#665700000000
0!
0%
#665705000000
1!
1%
#665710000000
0!
0%
#665715000000
1!
1%
#665720000000
0!
0%
#665725000000
1!
1%
#665730000000
0!
0%
#665735000000
1!
1%
#665740000000
0!
0%
#665745000000
1!
1%
#665750000000
0!
0%
#665755000000
1!
1%
#665760000000
0!
0%
#665765000000
1!
1%
#665770000000
0!
0%
#665775000000
1!
1%
#665780000000
0!
0%
#665785000000
1!
1%
#665790000000
0!
0%
#665795000000
1!
1%
#665800000000
0!
0%
#665805000000
1!
1%
#665810000000
0!
0%
#665815000000
1!
1%
#665820000000
0!
0%
#665825000000
1!
1%
#665830000000
0!
0%
#665835000000
1!
1%
#665840000000
0!
0%
#665845000000
1!
1%
#665850000000
0!
0%
#665855000000
1!
1%
#665860000000
0!
0%
#665865000000
1!
1%
#665870000000
0!
0%
#665875000000
1!
1%
#665880000000
0!
0%
#665885000000
1!
1%
#665890000000
0!
0%
#665895000000
1!
1%
#665900000000
0!
0%
#665905000000
1!
1%
#665910000000
0!
0%
#665915000000
1!
1%
#665920000000
0!
0%
#665925000000
1!
1%
#665930000000
0!
0%
#665935000000
1!
1%
#665940000000
0!
0%
#665945000000
1!
1%
#665950000000
0!
0%
#665955000000
1!
1%
#665960000000
0!
0%
#665965000000
1!
1%
#665970000000
0!
0%
#665975000000
1!
1%
#665980000000
0!
0%
#665985000000
1!
1%
#665990000000
0!
0%
#665995000000
1!
1%
#666000000000
0!
0%
#666005000000
1!
1%
#666010000000
0!
0%
#666015000000
1!
1%
#666020000000
0!
0%
#666025000000
1!
1%
#666030000000
0!
0%
#666035000000
1!
1%
#666040000000
0!
0%
#666045000000
1!
1%
#666050000000
0!
0%
#666055000000
1!
1%
#666060000000
0!
0%
#666065000000
1!
1%
#666070000000
0!
0%
#666075000000
1!
1%
#666080000000
0!
0%
#666085000000
1!
1%
#666090000000
0!
0%
#666095000000
1!
1%
#666100000000
0!
0%
#666105000000
1!
1%
#666110000000
0!
0%
#666115000000
1!
1%
#666120000000
0!
0%
#666125000000
1!
1%
#666130000000
0!
0%
#666135000000
1!
1%
#666140000000
0!
0%
#666145000000
1!
1%
#666150000000
0!
0%
#666155000000
1!
1%
#666160000000
0!
0%
#666165000000
1!
1%
#666170000000
0!
0%
#666175000000
1!
1%
#666180000000
0!
0%
#666185000000
1!
1%
#666190000000
0!
0%
#666195000000
1!
1%
#666200000000
0!
0%
#666205000000
1!
1%
#666210000000
0!
0%
#666215000000
1!
1%
#666220000000
0!
0%
#666225000000
1!
1%
#666230000000
0!
0%
#666235000000
1!
1%
#666240000000
0!
0%
#666245000000
1!
1%
#666250000000
0!
0%
#666255000000
1!
1%
#666260000000
0!
0%
#666265000000
1!
1%
#666270000000
0!
0%
#666275000000
1!
1%
#666280000000
0!
0%
#666285000000
1!
1%
#666290000000
0!
0%
#666295000000
1!
1%
#666300000000
0!
0%
#666305000000
1!
1%
#666310000000
0!
0%
#666315000000
1!
1%
#666320000000
0!
0%
#666325000000
1!
1%
#666330000000
0!
0%
#666335000000
1!
1%
#666340000000
0!
0%
#666345000000
1!
1%
#666350000000
0!
0%
#666355000000
1!
1%
#666360000000
0!
0%
#666365000000
1!
1%
#666370000000
0!
0%
#666375000000
1!
1%
#666380000000
0!
0%
#666385000000
1!
1%
#666390000000
0!
0%
#666395000000
1!
1%
#666400000000
0!
0%
#666405000000
1!
1%
#666410000000
0!
0%
#666415000000
1!
1%
#666420000000
0!
0%
#666425000000
1!
1%
#666430000000
0!
0%
#666435000000
1!
1%
#666440000000
0!
0%
#666445000000
1!
1%
#666450000000
0!
0%
#666455000000
1!
1%
#666460000000
0!
0%
#666465000000
1!
1%
#666470000000
0!
0%
#666475000000
1!
1%
#666480000000
0!
0%
#666485000000
1!
1%
#666490000000
0!
0%
#666495000000
1!
1%
#666500000000
0!
0%
#666505000000
1!
1%
#666510000000
0!
0%
#666515000000
1!
1%
#666520000000
0!
0%
#666525000000
1!
1%
#666530000000
0!
0%
#666535000000
1!
1%
#666540000000
0!
0%
#666545000000
1!
1%
#666550000000
0!
0%
#666555000000
1!
1%
#666560000000
0!
0%
#666565000000
1!
1%
#666570000000
0!
0%
#666575000000
1!
1%
#666580000000
0!
0%
#666585000000
1!
1%
#666590000000
0!
0%
#666595000000
1!
1%
#666600000000
0!
0%
#666605000000
1!
1%
#666610000000
0!
0%
#666615000000
1!
1%
#666620000000
0!
0%
#666625000000
1!
1%
#666630000000
0!
0%
#666635000000
1!
1%
#666640000000
0!
0%
#666645000000
1!
1%
#666650000000
0!
0%
#666655000000
1!
1%
#666660000000
0!
0%
#666665000000
1!
1%
#666670000000
0!
0%
#666675000000
1!
1%
#666680000000
0!
0%
#666685000000
1!
1%
#666690000000
0!
0%
#666695000000
1!
1%
#666700000000
0!
0%
#666705000000
1!
1%
#666710000000
0!
0%
#666715000000
1!
1%
#666720000000
0!
0%
#666725000000
1!
1%
#666730000000
0!
0%
#666735000000
1!
1%
#666740000000
0!
0%
#666745000000
1!
1%
#666750000000
0!
0%
#666755000000
1!
1%
#666760000000
0!
0%
#666765000000
1!
1%
#666770000000
0!
0%
#666775000000
1!
1%
#666780000000
0!
0%
#666785000000
1!
1%
#666790000000
0!
0%
#666795000000
1!
1%
#666800000000
0!
0%
#666805000000
1!
1%
#666810000000
0!
0%
#666815000000
1!
1%
#666820000000
0!
0%
#666825000000
1!
1%
#666830000000
0!
0%
#666835000000
1!
1%
#666840000000
0!
0%
#666845000000
1!
1%
#666850000000
0!
0%
#666855000000
1!
1%
#666860000000
0!
0%
#666865000000
1!
1%
#666870000000
0!
0%
#666875000000
1!
1%
#666880000000
0!
0%
#666885000000
1!
1%
#666890000000
0!
0%
#666895000000
1!
1%
#666900000000
0!
0%
#666905000000
1!
1%
#666910000000
0!
0%
#666915000000
1!
1%
#666920000000
0!
0%
#666925000000
1!
1%
#666930000000
0!
0%
#666935000000
1!
1%
#666940000000
0!
0%
#666945000000
1!
1%
#666950000000
0!
0%
#666955000000
1!
1%
#666960000000
0!
0%
#666965000000
1!
1%
#666970000000
0!
0%
#666975000000
1!
1%
#666980000000
0!
0%
#666985000000
1!
1%
#666990000000
0!
0%
#666995000000
1!
1%
#667000000000
0!
0%
#667005000000
1!
1%
#667010000000
0!
0%
#667015000000
1!
1%
#667020000000
0!
0%
#667025000000
1!
1%
#667030000000
0!
0%
#667035000000
1!
1%
#667040000000
0!
0%
#667045000000
1!
1%
#667050000000
0!
0%
#667055000000
1!
1%
#667060000000
0!
0%
#667065000000
1!
1%
#667070000000
0!
0%
#667075000000
1!
1%
#667080000000
0!
0%
#667085000000
1!
1%
#667090000000
0!
0%
#667095000000
1!
1%
#667100000000
0!
0%
#667105000000
1!
1%
#667110000000
0!
0%
#667115000000
1!
1%
#667120000000
0!
0%
#667125000000
1!
1%
#667130000000
0!
0%
#667135000000
1!
1%
#667140000000
0!
0%
#667145000000
1!
1%
#667150000000
0!
0%
#667155000000
1!
1%
#667160000000
0!
0%
#667165000000
1!
1%
#667170000000
0!
0%
#667175000000
1!
1%
#667180000000
0!
0%
#667185000000
1!
1%
#667190000000
0!
0%
#667195000000
1!
1%
#667200000000
0!
0%
#667205000000
1!
1%
#667210000000
0!
0%
#667215000000
1!
1%
#667220000000
0!
0%
#667225000000
1!
1%
#667230000000
0!
0%
#667235000000
1!
1%
#667240000000
0!
0%
#667245000000
1!
1%
#667250000000
0!
0%
#667255000000
1!
1%
#667260000000
0!
0%
#667265000000
1!
1%
#667270000000
0!
0%
#667275000000
1!
1%
#667280000000
0!
0%
#667285000000
1!
1%
#667290000000
0!
0%
#667295000000
1!
1%
#667300000000
0!
0%
#667305000000
1!
1%
#667310000000
0!
0%
#667315000000
1!
1%
#667320000000
0!
0%
#667325000000
1!
1%
#667330000000
0!
0%
#667335000000
1!
1%
#667340000000
0!
0%
#667345000000
1!
1%
#667350000000
0!
0%
#667355000000
1!
1%
#667360000000
0!
0%
#667365000000
1!
1%
#667370000000
0!
0%
#667375000000
1!
1%
#667380000000
0!
0%
#667385000000
1!
1%
#667390000000
0!
0%
#667395000000
1!
1%
#667400000000
0!
0%
#667405000000
1!
1%
#667410000000
0!
0%
#667415000000
1!
1%
#667420000000
0!
0%
#667425000000
1!
1%
#667430000000
0!
0%
#667435000000
1!
1%
#667440000000
0!
0%
#667445000000
1!
1%
#667450000000
0!
0%
#667455000000
1!
1%
#667460000000
0!
0%
#667465000000
1!
1%
#667470000000
0!
0%
#667475000000
1!
1%
#667480000000
0!
0%
#667485000000
1!
1%
#667490000000
0!
0%
#667495000000
1!
1%
#667500000000
0!
0%
#667505000000
1!
1%
#667510000000
0!
0%
#667515000000
1!
1%
#667520000000
0!
0%
#667525000000
1!
1%
#667530000000
0!
0%
#667535000000
1!
1%
#667540000000
0!
0%
#667545000000
1!
1%
#667550000000
0!
0%
#667555000000
1!
1%
#667560000000
0!
0%
#667565000000
1!
1%
#667570000000
0!
0%
#667575000000
1!
1%
#667580000000
0!
0%
#667585000000
1!
1%
#667590000000
0!
0%
#667595000000
1!
1%
#667600000000
0!
0%
#667605000000
1!
1%
#667610000000
0!
0%
#667615000000
1!
1%
#667620000000
0!
0%
#667625000000
1!
1%
#667630000000
0!
0%
#667635000000
1!
1%
#667640000000
0!
0%
#667645000000
1!
1%
#667650000000
0!
0%
#667655000000
1!
1%
#667660000000
0!
0%
#667665000000
1!
1%
#667670000000
0!
0%
#667675000000
1!
1%
#667680000000
0!
0%
#667685000000
1!
1%
#667690000000
0!
0%
#667695000000
1!
1%
#667700000000
0!
0%
#667705000000
1!
1%
#667710000000
0!
0%
#667715000000
1!
1%
#667720000000
0!
0%
#667725000000
1!
1%
#667730000000
0!
0%
#667735000000
1!
1%
#667740000000
0!
0%
#667745000000
1!
1%
#667750000000
0!
0%
#667755000000
1!
1%
#667760000000
0!
0%
#667765000000
1!
1%
#667770000000
0!
0%
#667775000000
1!
1%
#667780000000
0!
0%
#667785000000
1!
1%
#667790000000
0!
0%
#667795000000
1!
1%
#667800000000
0!
0%
#667805000000
1!
1%
#667810000000
0!
0%
#667815000000
1!
1%
#667820000000
0!
0%
#667825000000
1!
1%
#667830000000
0!
0%
#667835000000
1!
1%
#667840000000
0!
0%
#667845000000
1!
1%
#667850000000
0!
0%
#667855000000
1!
1%
#667860000000
0!
0%
#667865000000
1!
1%
#667870000000
0!
0%
#667875000000
1!
1%
#667880000000
0!
0%
#667885000000
1!
1%
#667890000000
0!
0%
#667895000000
1!
1%
#667900000000
0!
0%
#667905000000
1!
1%
#667910000000
0!
0%
#667915000000
1!
1%
#667920000000
0!
0%
#667925000000
1!
1%
#667930000000
0!
0%
#667935000000
1!
1%
#667940000000
0!
0%
#667945000000
1!
1%
#667950000000
0!
0%
#667955000000
1!
1%
#667960000000
0!
0%
#667965000000
1!
1%
#667970000000
0!
0%
#667975000000
1!
1%
#667980000000
0!
0%
#667985000000
1!
1%
#667990000000
0!
0%
#667995000000
1!
1%
#668000000000
0!
0%
#668005000000
1!
1%
#668010000000
0!
0%
#668015000000
1!
1%
#668020000000
0!
0%
#668025000000
1!
1%
#668030000000
0!
0%
#668035000000
1!
1%
#668040000000
0!
0%
#668045000000
1!
1%
#668050000000
0!
0%
#668055000000
1!
1%
#668060000000
0!
0%
#668065000000
1!
1%
#668070000000
0!
0%
#668075000000
1!
1%
#668080000000
0!
0%
#668085000000
1!
1%
#668090000000
0!
0%
#668095000000
1!
1%
#668100000000
0!
0%
#668105000000
1!
1%
#668110000000
0!
0%
#668115000000
1!
1%
#668120000000
0!
0%
#668125000000
1!
1%
#668130000000
0!
0%
#668135000000
1!
1%
#668140000000
0!
0%
#668145000000
1!
1%
#668150000000
0!
0%
#668155000000
1!
1%
#668160000000
0!
0%
#668165000000
1!
1%
#668170000000
0!
0%
#668175000000
1!
1%
#668180000000
0!
0%
#668185000000
1!
1%
#668190000000
0!
0%
#668195000000
1!
1%
#668200000000
0!
0%
#668205000000
1!
1%
#668210000000
0!
0%
#668215000000
1!
1%
#668220000000
0!
0%
#668225000000
1!
1%
#668230000000
0!
0%
#668235000000
1!
1%
#668240000000
0!
0%
#668245000000
1!
1%
#668250000000
0!
0%
#668255000000
1!
1%
#668260000000
0!
0%
#668265000000
1!
1%
#668270000000
0!
0%
#668275000000
1!
1%
#668280000000
0!
0%
#668285000000
1!
1%
#668290000000
0!
0%
#668295000000
1!
1%
#668300000000
0!
0%
#668305000000
1!
1%
#668310000000
0!
0%
#668315000000
1!
1%
#668320000000
0!
0%
#668325000000
1!
1%
#668330000000
0!
0%
#668335000000
1!
1%
#668340000000
0!
0%
#668345000000
1!
1%
#668350000000
0!
0%
#668355000000
1!
1%
#668360000000
0!
0%
#668365000000
1!
1%
#668370000000
0!
0%
#668375000000
1!
1%
#668380000000
0!
0%
#668385000000
1!
1%
#668390000000
0!
0%
#668395000000
1!
1%
#668400000000
0!
0%
#668405000000
1!
1%
#668410000000
0!
0%
#668415000000
1!
1%
#668420000000
0!
0%
#668425000000
1!
1%
#668430000000
0!
0%
#668435000000
1!
1%
#668440000000
0!
0%
#668445000000
1!
1%
#668450000000
0!
0%
#668455000000
1!
1%
#668460000000
0!
0%
#668465000000
1!
1%
#668470000000
0!
0%
#668475000000
1!
1%
#668480000000
0!
0%
#668485000000
1!
1%
#668490000000
0!
0%
#668495000000
1!
1%
#668500000000
0!
0%
#668505000000
1!
1%
#668510000000
0!
0%
#668515000000
1!
1%
#668520000000
0!
0%
#668525000000
1!
1%
#668530000000
0!
0%
#668535000000
1!
1%
#668540000000
0!
0%
#668545000000
1!
1%
#668550000000
0!
0%
#668555000000
1!
1%
#668560000000
0!
0%
#668565000000
1!
1%
#668570000000
0!
0%
#668575000000
1!
1%
#668580000000
0!
0%
#668585000000
1!
1%
#668590000000
0!
0%
#668595000000
1!
1%
#668600000000
0!
0%
#668605000000
1!
1%
#668610000000
0!
0%
#668615000000
1!
1%
#668620000000
0!
0%
#668625000000
1!
1%
#668630000000
0!
0%
#668635000000
1!
1%
#668640000000
0!
0%
#668645000000
1!
1%
#668650000000
0!
0%
#668655000000
1!
1%
#668660000000
0!
0%
#668665000000
1!
1%
#668670000000
0!
0%
#668675000000
1!
1%
#668680000000
0!
0%
#668685000000
1!
1%
#668690000000
0!
0%
#668695000000
1!
1%
#668700000000
0!
0%
#668705000000
1!
1%
#668710000000
0!
0%
#668715000000
1!
1%
#668720000000
0!
0%
#668725000000
1!
1%
#668730000000
0!
0%
#668735000000
1!
1%
#668740000000
0!
0%
#668745000000
1!
1%
#668750000000
0!
0%
#668755000000
1!
1%
#668760000000
0!
0%
#668765000000
1!
1%
#668770000000
0!
0%
#668775000000
1!
1%
#668780000000
0!
0%
#668785000000
1!
1%
#668790000000
0!
0%
#668795000000
1!
1%
#668800000000
0!
0%
#668805000000
1!
1%
#668810000000
0!
0%
#668815000000
1!
1%
#668820000000
0!
0%
#668825000000
1!
1%
#668830000000
0!
0%
#668835000000
1!
1%
#668840000000
0!
0%
#668845000000
1!
1%
#668850000000
0!
0%
#668855000000
1!
1%
#668860000000
0!
0%
#668865000000
1!
1%
#668870000000
0!
0%
#668875000000
1!
1%
#668880000000
0!
0%
#668885000000
1!
1%
#668890000000
0!
0%
#668895000000
1!
1%
#668900000000
0!
0%
#668905000000
1!
1%
#668910000000
0!
0%
#668915000000
1!
1%
#668920000000
0!
0%
#668925000000
1!
1%
#668930000000
0!
0%
#668935000000
1!
1%
#668940000000
0!
0%
#668945000000
1!
1%
#668950000000
0!
0%
#668955000000
1!
1%
#668960000000
0!
0%
#668965000000
1!
1%
#668970000000
0!
0%
#668975000000
1!
1%
#668980000000
0!
0%
#668985000000
1!
1%
#668990000000
0!
0%
#668995000000
1!
1%
#669000000000
0!
0%
#669005000000
1!
1%
#669010000000
0!
0%
#669015000000
1!
1%
#669020000000
0!
0%
#669025000000
1!
1%
#669030000000
0!
0%
#669035000000
1!
1%
#669040000000
0!
0%
#669045000000
1!
1%
#669050000000
0!
0%
#669055000000
1!
1%
#669060000000
0!
0%
#669065000000
1!
1%
#669070000000
0!
0%
#669075000000
1!
1%
#669080000000
0!
0%
#669085000000
1!
1%
#669090000000
0!
0%
#669095000000
1!
1%
#669100000000
0!
0%
#669105000000
1!
1%
#669110000000
0!
0%
#669115000000
1!
1%
#669120000000
0!
0%
#669125000000
1!
1%
#669130000000
0!
0%
#669135000000
1!
1%
#669140000000
0!
0%
#669145000000
1!
1%
#669150000000
0!
0%
#669155000000
1!
1%
#669160000000
0!
0%
#669165000000
1!
1%
#669170000000
0!
0%
#669175000000
1!
1%
#669180000000
0!
0%
#669185000000
1!
1%
#669190000000
0!
0%
#669195000000
1!
1%
#669200000000
0!
0%
#669205000000
1!
1%
#669210000000
0!
0%
#669215000000
1!
1%
#669220000000
0!
0%
#669225000000
1!
1%
#669230000000
0!
0%
#669235000000
1!
1%
#669240000000
0!
0%
#669245000000
1!
1%
#669250000000
0!
0%
#669255000000
1!
1%
#669260000000
0!
0%
#669265000000
1!
1%
#669270000000
0!
0%
#669275000000
1!
1%
#669280000000
0!
0%
#669285000000
1!
1%
#669290000000
0!
0%
#669295000000
1!
1%
#669300000000
0!
0%
#669305000000
1!
1%
#669310000000
0!
0%
#669315000000
1!
1%
#669320000000
0!
0%
#669325000000
1!
1%
#669330000000
0!
0%
#669335000000
1!
1%
#669340000000
0!
0%
#669345000000
1!
1%
#669350000000
0!
0%
#669355000000
1!
1%
#669360000000
0!
0%
#669365000000
1!
1%
#669370000000
0!
0%
#669375000000
1!
1%
#669380000000
0!
0%
#669385000000
1!
1%
#669390000000
0!
0%
#669395000000
1!
1%
#669400000000
0!
0%
#669405000000
1!
1%
#669410000000
0!
0%
#669415000000
1!
1%
#669420000000
0!
0%
#669425000000
1!
1%
#669430000000
0!
0%
#669435000000
1!
1%
#669440000000
0!
0%
#669445000000
1!
1%
#669450000000
0!
0%
#669455000000
1!
1%
#669460000000
0!
0%
#669465000000
1!
1%
#669470000000
0!
0%
#669475000000
1!
1%
#669480000000
0!
0%
#669485000000
1!
1%
#669490000000
0!
0%
#669495000000
1!
1%
#669500000000
0!
0%
#669505000000
1!
1%
#669510000000
0!
0%
#669515000000
1!
1%
#669520000000
0!
0%
#669525000000
1!
1%
#669530000000
0!
0%
#669535000000
1!
1%
#669540000000
0!
0%
#669545000000
1!
1%
#669550000000
0!
0%
#669555000000
1!
1%
#669560000000
0!
0%
#669565000000
1!
1%
#669570000000
0!
0%
#669575000000
1!
1%
#669580000000
0!
0%
#669585000000
1!
1%
#669590000000
0!
0%
#669595000000
1!
1%
#669600000000
0!
0%
#669605000000
1!
1%
#669610000000
0!
0%
#669615000000
1!
1%
#669620000000
0!
0%
#669625000000
1!
1%
#669630000000
0!
0%
#669635000000
1!
1%
#669640000000
0!
0%
#669645000000
1!
1%
#669650000000
0!
0%
#669655000000
1!
1%
#669660000000
0!
0%
#669665000000
1!
1%
#669670000000
0!
0%
#669675000000
1!
1%
#669680000000
0!
0%
#669685000000
1!
1%
#669690000000
0!
0%
#669695000000
1!
1%
#669700000000
0!
0%
#669705000000
1!
1%
#669710000000
0!
0%
#669715000000
1!
1%
#669720000000
0!
0%
#669725000000
1!
1%
#669730000000
0!
0%
#669735000000
1!
1%
#669740000000
0!
0%
#669745000000
1!
1%
#669750000000
0!
0%
#669755000000
1!
1%
#669760000000
0!
0%
#669765000000
1!
1%
#669770000000
0!
0%
#669775000000
1!
1%
#669780000000
0!
0%
#669785000000
1!
1%
#669790000000
0!
0%
#669795000000
1!
1%
#669800000000
0!
0%
#669805000000
1!
1%
#669810000000
0!
0%
#669815000000
1!
1%
#669820000000
0!
0%
#669825000000
1!
1%
#669830000000
0!
0%
#669835000000
1!
1%
#669840000000
0!
0%
#669845000000
1!
1%
#669850000000
0!
0%
#669855000000
1!
1%
#669860000000
0!
0%
#669865000000
1!
1%
#669870000000
0!
0%
#669875000000
1!
1%
#669880000000
0!
0%
#669885000000
1!
1%
#669890000000
0!
0%
#669895000000
1!
1%
#669900000000
0!
0%
#669905000000
1!
1%
#669910000000
0!
0%
#669915000000
1!
1%
#669920000000
0!
0%
#669925000000
1!
1%
#669930000000
0!
0%
#669935000000
1!
1%
#669940000000
0!
0%
#669945000000
1!
1%
#669950000000
0!
0%
#669955000000
1!
1%
#669960000000
0!
0%
#669965000000
1!
1%
#669970000000
0!
0%
#669975000000
1!
1%
#669980000000
0!
0%
#669985000000
1!
1%
#669990000000
0!
0%
#669995000000
1!
1%
#670000000000
0!
0%
#670005000000
1!
1%
#670010000000
0!
0%
#670015000000
1!
1%
#670020000000
0!
0%
#670025000000
1!
1%
#670030000000
0!
0%
#670035000000
1!
1%
#670040000000
0!
0%
#670045000000
1!
1%
#670050000000
0!
0%
#670055000000
1!
1%
#670060000000
0!
0%
#670065000000
1!
1%
#670070000000
0!
0%
#670075000000
1!
1%
#670080000000
0!
0%
#670085000000
1!
1%
#670090000000
0!
0%
#670095000000
1!
1%
#670100000000
0!
0%
#670105000000
1!
1%
#670110000000
0!
0%
#670115000000
1!
1%
#670120000000
0!
0%
#670125000000
1!
1%
#670130000000
0!
0%
#670135000000
1!
1%
#670140000000
0!
0%
#670145000000
1!
1%
#670150000000
0!
0%
#670155000000
1!
1%
#670160000000
0!
0%
#670165000000
1!
1%
#670170000000
0!
0%
#670175000000
1!
1%
#670180000000
0!
0%
#670185000000
1!
1%
#670190000000
0!
0%
#670195000000
1!
1%
#670200000000
0!
0%
#670205000000
1!
1%
#670210000000
0!
0%
#670215000000
1!
1%
#670220000000
0!
0%
#670225000000
1!
1%
#670230000000
0!
0%
#670235000000
1!
1%
#670240000000
0!
0%
#670245000000
1!
1%
#670250000000
0!
0%
#670255000000
1!
1%
#670260000000
0!
0%
#670265000000
1!
1%
#670270000000
0!
0%
#670275000000
1!
1%
#670280000000
0!
0%
#670285000000
1!
1%
#670290000000
0!
0%
#670295000000
1!
1%
#670300000000
0!
0%
#670305000000
1!
1%
#670310000000
0!
0%
#670315000000
1!
1%
#670320000000
0!
0%
#670325000000
1!
1%
#670330000000
0!
0%
#670335000000
1!
1%
#670340000000
0!
0%
#670345000000
1!
1%
#670350000000
0!
0%
#670355000000
1!
1%
#670360000000
0!
0%
#670365000000
1!
1%
#670370000000
0!
0%
#670375000000
1!
1%
#670380000000
0!
0%
#670385000000
1!
1%
#670390000000
0!
0%
#670395000000
1!
1%
#670400000000
0!
0%
#670405000000
1!
1%
#670410000000
0!
0%
#670415000000
1!
1%
#670420000000
0!
0%
#670425000000
1!
1%
#670430000000
0!
0%
#670435000000
1!
1%
#670440000000
0!
0%
#670445000000
1!
1%
#670450000000
0!
0%
#670455000000
1!
1%
#670460000000
0!
0%
#670465000000
1!
1%
#670470000000
0!
0%
#670475000000
1!
1%
#670480000000
0!
0%
#670485000000
1!
1%
#670490000000
0!
0%
#670495000000
1!
1%
#670500000000
0!
0%
#670505000000
1!
1%
#670510000000
0!
0%
#670515000000
1!
1%
#670520000000
0!
0%
#670525000000
1!
1%
#670530000000
0!
0%
#670535000000
1!
1%
#670540000000
0!
0%
#670545000000
1!
1%
#670550000000
0!
0%
#670555000000
1!
1%
#670560000000
0!
0%
#670565000000
1!
1%
#670570000000
0!
0%
#670575000000
1!
1%
#670580000000
0!
0%
#670585000000
1!
1%
#670590000000
0!
0%
#670595000000
1!
1%
#670600000000
0!
0%
#670605000000
1!
1%
#670610000000
0!
0%
#670615000000
1!
1%
#670620000000
0!
0%
#670625000000
1!
1%
#670630000000
0!
0%
#670635000000
1!
1%
#670640000000
0!
0%
#670645000000
1!
1%
#670650000000
0!
0%
#670655000000
1!
1%
#670660000000
0!
0%
#670665000000
1!
1%
#670670000000
0!
0%
#670675000000
1!
1%
#670680000000
0!
0%
#670685000000
1!
1%
#670690000000
0!
0%
#670695000000
1!
1%
#670700000000
0!
0%
#670705000000
1!
1%
#670710000000
0!
0%
#670715000000
1!
1%
#670720000000
0!
0%
#670725000000
1!
1%
#670730000000
0!
0%
#670735000000
1!
1%
#670740000000
0!
0%
#670745000000
1!
1%
#670750000000
0!
0%
#670755000000
1!
1%
#670760000000
0!
0%
#670765000000
1!
1%
#670770000000
0!
0%
#670775000000
1!
1%
#670780000000
0!
0%
#670785000000
1!
1%
#670790000000
0!
0%
#670795000000
1!
1%
#670800000000
0!
0%
#670805000000
1!
1%
#670810000000
0!
0%
#670815000000
1!
1%
#670820000000
0!
0%
#670825000000
1!
1%
#670830000000
0!
0%
#670835000000
1!
1%
#670840000000
0!
0%
#670845000000
1!
1%
#670850000000
0!
0%
#670855000000
1!
1%
#670860000000
0!
0%
#670865000000
1!
1%
#670870000000
0!
0%
#670875000000
1!
1%
#670880000000
0!
0%
#670885000000
1!
1%
#670890000000
0!
0%
#670895000000
1!
1%
#670900000000
0!
0%
#670905000000
1!
1%
#670910000000
0!
0%
#670915000000
1!
1%
#670920000000
0!
0%
#670925000000
1!
1%
#670930000000
0!
0%
#670935000000
1!
1%
#670940000000
0!
0%
#670945000000
1!
1%
#670950000000
0!
0%
#670955000000
1!
1%
#670960000000
0!
0%
#670965000000
1!
1%
#670970000000
0!
0%
#670975000000
1!
1%
#670980000000
0!
0%
#670985000000
1!
1%
#670990000000
0!
0%
#670995000000
1!
1%
#671000000000
0!
0%
#671005000000
1!
1%
#671010000000
0!
0%
#671015000000
1!
1%
#671020000000
0!
0%
#671025000000
1!
1%
#671030000000
0!
0%
#671035000000
1!
1%
#671040000000
0!
0%
#671045000000
1!
1%
#671050000000
0!
0%
#671055000000
1!
1%
#671060000000
0!
0%
#671065000000
1!
1%
#671070000000
0!
0%
#671075000000
1!
1%
#671080000000
0!
0%
#671085000000
1!
1%
#671090000000
0!
0%
#671095000000
1!
1%
#671100000000
0!
0%
#671105000000
1!
1%
#671110000000
0!
0%
#671115000000
1!
1%
#671120000000
0!
0%
#671125000000
1!
1%
#671130000000
0!
0%
#671135000000
1!
1%
#671140000000
0!
0%
#671145000000
1!
1%
#671150000000
0!
0%
#671155000000
1!
1%
#671160000000
0!
0%
#671165000000
1!
1%
#671170000000
0!
0%
#671175000000
1!
1%
#671180000000
0!
0%
#671185000000
1!
1%
#671190000000
0!
0%
#671195000000
1!
1%
#671200000000
0!
0%
#671205000000
1!
1%
#671210000000
0!
0%
#671215000000
1!
1%
#671220000000
0!
0%
#671225000000
1!
1%
#671230000000
0!
0%
#671235000000
1!
1%
#671240000000
0!
0%
#671245000000
1!
1%
#671250000000
0!
0%
#671255000000
1!
1%
#671260000000
0!
0%
#671265000000
1!
1%
#671270000000
0!
0%
#671275000000
1!
1%
#671280000000
0!
0%
#671285000000
1!
1%
#671290000000
0!
0%
#671295000000
1!
1%
#671300000000
0!
0%
#671305000000
1!
1%
#671310000000
0!
0%
#671315000000
1!
1%
#671320000000
0!
0%
#671325000000
1!
1%
#671330000000
0!
0%
#671335000000
1!
1%
#671340000000
0!
0%
#671345000000
1!
1%
#671350000000
0!
0%
#671355000000
1!
1%
#671360000000
0!
0%
#671365000000
1!
1%
#671370000000
0!
0%
#671375000000
1!
1%
#671380000000
0!
0%
#671385000000
1!
1%
#671390000000
0!
0%
#671395000000
1!
1%
#671400000000
0!
0%
#671405000000
1!
1%
#671410000000
0!
0%
#671415000000
1!
1%
#671420000000
0!
0%
#671425000000
1!
1%
#671430000000
0!
0%
#671435000000
1!
1%
#671440000000
0!
0%
#671445000000
1!
1%
#671450000000
0!
0%
#671455000000
1!
1%
#671460000000
0!
0%
#671465000000
1!
1%
#671470000000
0!
0%
#671475000000
1!
1%
#671480000000
0!
0%
#671485000000
1!
1%
#671490000000
0!
0%
#671495000000
1!
1%
#671500000000
0!
0%
#671505000000
1!
1%
#671510000000
0!
0%
#671515000000
1!
1%
#671520000000
0!
0%
#671525000000
1!
1%
#671530000000
0!
0%
#671535000000
1!
1%
#671540000000
0!
0%
#671545000000
1!
1%
#671550000000
0!
0%
#671555000000
1!
1%
#671560000000
0!
0%
#671565000000
1!
1%
#671570000000
0!
0%
#671575000000
1!
1%
#671580000000
0!
0%
#671585000000
1!
1%
#671590000000
0!
0%
#671595000000
1!
1%
#671600000000
0!
0%
#671605000000
1!
1%
#671610000000
0!
0%
#671615000000
1!
1%
#671620000000
0!
0%
#671625000000
1!
1%
#671630000000
0!
0%
#671635000000
1!
1%
#671640000000
0!
0%
#671645000000
1!
1%
#671650000000
0!
0%
#671655000000
1!
1%
#671660000000
0!
0%
#671665000000
1!
1%
#671670000000
0!
0%
#671675000000
1!
1%
#671680000000
0!
0%
#671685000000
1!
1%
#671690000000
0!
0%
#671695000000
1!
1%
#671700000000
0!
0%
#671705000000
1!
1%
#671710000000
0!
0%
#671715000000
1!
1%
#671720000000
0!
0%
#671725000000
1!
1%
#671730000000
0!
0%
#671735000000
1!
1%
#671740000000
0!
0%
#671745000000
1!
1%
#671750000000
0!
0%
#671755000000
1!
1%
#671760000000
0!
0%
#671765000000
1!
1%
#671770000000
0!
0%
#671775000000
1!
1%
#671780000000
0!
0%
#671785000000
1!
1%
#671790000000
0!
0%
#671795000000
1!
1%
#671800000000
0!
0%
#671805000000
1!
1%
#671810000000
0!
0%
#671815000000
1!
1%
#671820000000
0!
0%
#671825000000
1!
1%
#671830000000
0!
0%
#671835000000
1!
1%
#671840000000
0!
0%
#671845000000
1!
1%
#671850000000
0!
0%
#671855000000
1!
1%
#671860000000
0!
0%
#671865000000
1!
1%
#671870000000
0!
0%
#671875000000
1!
1%
#671880000000
0!
0%
#671885000000
1!
1%
#671890000000
0!
0%
#671895000000
1!
1%
#671900000000
0!
0%
#671905000000
1!
1%
#671910000000
0!
0%
#671915000000
1!
1%
#671920000000
0!
0%
#671925000000
1!
1%
#671930000000
0!
0%
#671935000000
1!
1%
#671940000000
0!
0%
#671945000000
1!
1%
#671950000000
0!
0%
#671955000000
1!
1%
#671960000000
0!
0%
#671965000000
1!
1%
#671970000000
0!
0%
#671975000000
1!
1%
#671980000000
0!
0%
#671985000000
1!
1%
#671990000000
0!
0%
#671995000000
1!
1%
#672000000000
0!
0%
#672005000000
1!
1%
#672010000000
0!
0%
#672015000000
1!
1%
#672020000000
0!
0%
#672025000000
1!
1%
#672030000000
0!
0%
#672035000000
1!
1%
#672040000000
0!
0%
#672045000000
1!
1%
#672050000000
0!
0%
#672055000000
1!
1%
#672060000000
0!
0%
#672065000000
1!
1%
#672070000000
0!
0%
#672075000000
1!
1%
#672080000000
0!
0%
#672085000000
1!
1%
#672090000000
0!
0%
#672095000000
1!
1%
#672100000000
0!
0%
#672105000000
1!
1%
#672110000000
0!
0%
#672115000000
1!
1%
#672120000000
0!
0%
#672125000000
1!
1%
#672130000000
0!
0%
#672135000000
1!
1%
#672140000000
0!
0%
#672145000000
1!
1%
#672150000000
0!
0%
#672155000000
1!
1%
#672160000000
0!
0%
#672165000000
1!
1%
#672170000000
0!
0%
#672175000000
1!
1%
#672180000000
0!
0%
#672185000000
1!
1%
#672190000000
0!
0%
#672195000000
1!
1%
#672200000000
0!
0%
#672205000000
1!
1%
#672210000000
0!
0%
#672215000000
1!
1%
#672220000000
0!
0%
#672225000000
1!
1%
#672230000000
0!
0%
#672235000000
1!
1%
#672240000000
0!
0%
#672245000000
1!
1%
#672250000000
0!
0%
#672255000000
1!
1%
#672260000000
0!
0%
#672265000000
1!
1%
#672270000000
0!
0%
#672275000000
1!
1%
#672280000000
0!
0%
#672285000000
1!
1%
#672290000000
0!
0%
#672295000000
1!
1%
#672300000000
0!
0%
#672305000000
1!
1%
#672310000000
0!
0%
#672315000000
1!
1%
#672320000000
0!
0%
#672325000000
1!
1%
#672330000000
0!
0%
#672335000000
1!
1%
#672340000000
0!
0%
#672345000000
1!
1%
#672350000000
0!
0%
#672355000000
1!
1%
#672360000000
0!
0%
#672365000000
1!
1%
#672370000000
0!
0%
#672375000000
1!
1%
#672380000000
0!
0%
#672385000000
1!
1%
#672390000000
0!
0%
#672395000000
1!
1%
#672400000000
0!
0%
#672405000000
1!
1%
#672410000000
0!
0%
#672415000000
1!
1%
#672420000000
0!
0%
#672425000000
1!
1%
#672430000000
0!
0%
#672435000000
1!
1%
#672440000000
0!
0%
#672445000000
1!
1%
#672450000000
0!
0%
#672455000000
1!
1%
#672460000000
0!
0%
#672465000000
1!
1%
#672470000000
0!
0%
#672475000000
1!
1%
#672480000000
0!
0%
#672485000000
1!
1%
#672490000000
0!
0%
#672495000000
1!
1%
#672500000000
0!
0%
#672505000000
1!
1%
#672510000000
0!
0%
#672515000000
1!
1%
#672520000000
0!
0%
#672525000000
1!
1%
#672530000000
0!
0%
#672535000000
1!
1%
#672540000000
0!
0%
#672545000000
1!
1%
#672550000000
0!
0%
#672555000000
1!
1%
#672560000000
0!
0%
#672565000000
1!
1%
#672570000000
0!
0%
#672575000000
1!
1%
#672580000000
0!
0%
#672585000000
1!
1%
#672590000000
0!
0%
#672595000000
1!
1%
#672600000000
0!
0%
#672605000000
1!
1%
#672610000000
0!
0%
#672615000000
1!
1%
#672620000000
0!
0%
#672625000000
1!
1%
#672630000000
0!
0%
#672635000000
1!
1%
#672640000000
0!
0%
#672645000000
1!
1%
#672650000000
0!
0%
#672655000000
1!
1%
#672660000000
0!
0%
#672665000000
1!
1%
#672670000000
0!
0%
#672675000000
1!
1%
#672680000000
0!
0%
#672685000000
1!
1%
#672690000000
0!
0%
#672695000000
1!
1%
#672700000000
0!
0%
#672705000000
1!
1%
#672710000000
0!
0%
#672715000000
1!
1%
#672720000000
0!
0%
#672725000000
1!
1%
#672730000000
0!
0%
#672735000000
1!
1%
#672740000000
0!
0%
#672745000000
1!
1%
#672750000000
0!
0%
#672755000000
1!
1%
#672760000000
0!
0%
#672765000000
1!
1%
#672770000000
0!
0%
#672775000000
1!
1%
#672780000000
0!
0%
#672785000000
1!
1%
#672790000000
0!
0%
#672795000000
1!
1%
#672800000000
0!
0%
#672805000000
1!
1%
#672810000000
0!
0%
#672815000000
1!
1%
#672820000000
0!
0%
#672825000000
1!
1%
#672830000000
0!
0%
#672835000000
1!
1%
#672840000000
0!
0%
#672845000000
1!
1%
#672850000000
0!
0%
#672855000000
1!
1%
#672860000000
0!
0%
#672865000000
1!
1%
#672870000000
0!
0%
#672875000000
1!
1%
#672880000000
0!
0%
#672885000000
1!
1%
#672890000000
0!
0%
#672895000000
1!
1%
#672900000000
0!
0%
#672905000000
1!
1%
#672910000000
0!
0%
#672915000000
1!
1%
#672920000000
0!
0%
#672925000000
1!
1%
#672930000000
0!
0%
#672935000000
1!
1%
#672940000000
0!
0%
#672945000000
1!
1%
#672950000000
0!
0%
#672955000000
1!
1%
#672960000000
0!
0%
#672965000000
1!
1%
#672970000000
0!
0%
#672975000000
1!
1%
#672980000000
0!
0%
#672985000000
1!
1%
#672990000000
0!
0%
#672995000000
1!
1%
#673000000000
0!
0%
#673005000000
1!
1%
#673010000000
0!
0%
#673015000000
1!
1%
#673020000000
0!
0%
#673025000000
1!
1%
#673030000000
0!
0%
#673035000000
1!
1%
#673040000000
0!
0%
#673045000000
1!
1%
#673050000000
0!
0%
#673055000000
1!
1%
#673060000000
0!
0%
#673065000000
1!
1%
#673070000000
0!
0%
#673075000000
1!
1%
#673080000000
0!
0%
#673085000000
1!
1%
#673090000000
0!
0%
#673095000000
1!
1%
#673100000000
0!
0%
#673105000000
1!
1%
#673110000000
0!
0%
#673115000000
1!
1%
#673120000000
0!
0%
#673125000000
1!
1%
#673130000000
0!
0%
#673135000000
1!
1%
#673140000000
0!
0%
#673145000000
1!
1%
#673150000000
0!
0%
#673155000000
1!
1%
#673160000000
0!
0%
#673165000000
1!
1%
#673170000000
0!
0%
#673175000000
1!
1%
#673180000000
0!
0%
#673185000000
1!
1%
#673190000000
0!
0%
#673195000000
1!
1%
#673200000000
0!
0%
#673205000000
1!
1%
#673210000000
0!
0%
#673215000000
1!
1%
#673220000000
0!
0%
#673225000000
1!
1%
#673230000000
0!
0%
#673235000000
1!
1%
#673240000000
0!
0%
#673245000000
1!
1%
#673250000000
0!
0%
#673255000000
1!
1%
#673260000000
0!
0%
#673265000000
1!
1%
#673270000000
0!
0%
#673275000000
1!
1%
#673280000000
0!
0%
#673285000000
1!
1%
#673290000000
0!
0%
#673295000000
1!
1%
#673300000000
0!
0%
#673305000000
1!
1%
#673310000000
0!
0%
#673315000000
1!
1%
#673320000000
0!
0%
#673325000000
1!
1%
#673330000000
0!
0%
#673335000000
1!
1%
#673340000000
0!
0%
#673345000000
1!
1%
#673350000000
0!
0%
#673355000000
1!
1%
#673360000000
0!
0%
#673365000000
1!
1%
#673370000000
0!
0%
#673375000000
1!
1%
#673380000000
0!
0%
#673385000000
1!
1%
#673390000000
0!
0%
#673395000000
1!
1%
#673400000000
0!
0%
#673405000000
1!
1%
#673410000000
0!
0%
#673415000000
1!
1%
#673420000000
0!
0%
#673425000000
1!
1%
#673430000000
0!
0%
#673435000000
1!
1%
#673440000000
0!
0%
#673445000000
1!
1%
#673450000000
0!
0%
#673455000000
1!
1%
#673460000000
0!
0%
#673465000000
1!
1%
#673470000000
0!
0%
#673475000000
1!
1%
#673480000000
0!
0%
#673485000000
1!
1%
#673490000000
0!
0%
#673495000000
1!
1%
#673500000000
0!
0%
#673505000000
1!
1%
#673510000000
0!
0%
#673515000000
1!
1%
#673520000000
0!
0%
#673525000000
1!
1%
#673530000000
0!
0%
#673535000000
1!
1%
#673540000000
0!
0%
#673545000000
1!
1%
#673550000000
0!
0%
#673555000000
1!
1%
#673560000000
0!
0%
#673565000000
1!
1%
#673570000000
0!
0%
#673575000000
1!
1%
#673580000000
0!
0%
#673585000000
1!
1%
#673590000000
0!
0%
#673595000000
1!
1%
#673600000000
0!
0%
#673605000000
1!
1%
#673610000000
0!
0%
#673615000000
1!
1%
#673620000000
0!
0%
#673625000000
1!
1%
#673630000000
0!
0%
#673635000000
1!
1%
#673640000000
0!
0%
#673645000000
1!
1%
#673650000000
0!
0%
#673655000000
1!
1%
#673660000000
0!
0%
#673665000000
1!
1%
#673670000000
0!
0%
#673675000000
1!
1%
#673680000000
0!
0%
#673685000000
1!
1%
#673690000000
0!
0%
#673695000000
1!
1%
#673700000000
0!
0%
#673705000000
1!
1%
#673710000000
0!
0%
#673715000000
1!
1%
#673720000000
0!
0%
#673725000000
1!
1%
#673730000000
0!
0%
#673735000000
1!
1%
#673740000000
0!
0%
#673745000000
1!
1%
#673750000000
0!
0%
#673755000000
1!
1%
#673760000000
0!
0%
#673765000000
1!
1%
#673770000000
0!
0%
#673775000000
1!
1%
#673780000000
0!
0%
#673785000000
1!
1%
#673790000000
0!
0%
#673795000000
1!
1%
#673800000000
0!
0%
#673805000000
1!
1%
#673810000000
0!
0%
#673815000000
1!
1%
#673820000000
0!
0%
#673825000000
1!
1%
#673830000000
0!
0%
#673835000000
1!
1%
#673840000000
0!
0%
#673845000000
1!
1%
#673850000000
0!
0%
#673855000000
1!
1%
#673860000000
0!
0%
#673865000000
1!
1%
#673870000000
0!
0%
#673875000000
1!
1%
#673880000000
0!
0%
#673885000000
1!
1%
#673890000000
0!
0%
#673895000000
1!
1%
#673900000000
0!
0%
#673905000000
1!
1%
#673910000000
0!
0%
#673915000000
1!
1%
#673920000000
0!
0%
#673925000000
1!
1%
#673930000000
0!
0%
#673935000000
1!
1%
#673940000000
0!
0%
#673945000000
1!
1%
#673950000000
0!
0%
#673955000000
1!
1%
#673960000000
0!
0%
#673965000000
1!
1%
#673970000000
0!
0%
#673975000000
1!
1%
#673980000000
0!
0%
#673985000000
1!
1%
#673990000000
0!
0%
#673995000000
1!
1%
#674000000000
0!
0%
#674005000000
1!
1%
#674010000000
0!
0%
#674015000000
1!
1%
#674020000000
0!
0%
#674025000000
1!
1%
#674030000000
0!
0%
#674035000000
1!
1%
#674040000000
0!
0%
#674045000000
1!
1%
#674050000000
0!
0%
#674055000000
1!
1%
#674060000000
0!
0%
#674065000000
1!
1%
#674070000000
0!
0%
#674075000000
1!
1%
#674080000000
0!
0%
#674085000000
1!
1%
#674090000000
0!
0%
#674095000000
1!
1%
#674100000000
0!
0%
#674105000000
1!
1%
#674110000000
0!
0%
#674115000000
1!
1%
#674120000000
0!
0%
#674125000000
1!
1%
#674130000000
0!
0%
#674135000000
1!
1%
#674140000000
0!
0%
#674145000000
1!
1%
#674150000000
0!
0%
#674155000000
1!
1%
#674160000000
0!
0%
#674165000000
1!
1%
#674170000000
0!
0%
#674175000000
1!
1%
#674180000000
0!
0%
#674185000000
1!
1%
#674190000000
0!
0%
#674195000000
1!
1%
#674200000000
0!
0%
#674205000000
1!
1%
#674210000000
0!
0%
#674215000000
1!
1%
#674220000000
0!
0%
#674225000000
1!
1%
#674230000000
0!
0%
#674235000000
1!
1%
#674240000000
0!
0%
#674245000000
1!
1%
#674250000000
0!
0%
#674255000000
1!
1%
#674260000000
0!
0%
#674265000000
1!
1%
#674270000000
0!
0%
#674275000000
1!
1%
#674280000000
0!
0%
#674285000000
1!
1%
#674290000000
0!
0%
#674295000000
1!
1%
#674300000000
0!
0%
#674305000000
1!
1%
#674310000000
0!
0%
#674315000000
1!
1%
#674320000000
0!
0%
#674325000000
1!
1%
#674330000000
0!
0%
#674335000000
1!
1%
#674340000000
0!
0%
#674345000000
1!
1%
#674350000000
0!
0%
#674355000000
1!
1%
#674360000000
0!
0%
#674365000000
1!
1%
#674370000000
0!
0%
#674375000000
1!
1%
#674380000000
0!
0%
#674385000000
1!
1%
#674390000000
0!
0%
#674395000000
1!
1%
#674400000000
0!
0%
#674405000000
1!
1%
#674410000000
0!
0%
#674415000000
1!
1%
#674420000000
0!
0%
#674425000000
1!
1%
#674430000000
0!
0%
#674435000000
1!
1%
#674440000000
0!
0%
#674445000000
1!
1%
#674450000000
0!
0%
#674455000000
1!
1%
#674460000000
0!
0%
#674465000000
1!
1%
#674470000000
0!
0%
#674475000000
1!
1%
#674480000000
0!
0%
#674485000000
1!
1%
#674490000000
0!
0%
#674495000000
1!
1%
#674500000000
0!
0%
#674505000000
1!
1%
#674510000000
0!
0%
#674515000000
1!
1%
#674520000000
0!
0%
#674525000000
1!
1%
#674530000000
0!
0%
#674535000000
1!
1%
#674540000000
0!
0%
#674545000000
1!
1%
#674550000000
0!
0%
#674555000000
1!
1%
#674560000000
0!
0%
#674565000000
1!
1%
#674570000000
0!
0%
#674575000000
1!
1%
#674580000000
0!
0%
#674585000000
1!
1%
#674590000000
0!
0%
#674595000000
1!
1%
#674600000000
0!
0%
#674605000000
1!
1%
#674610000000
0!
0%
#674615000000
1!
1%
#674620000000
0!
0%
#674625000000
1!
1%
#674630000000
0!
0%
#674635000000
1!
1%
#674640000000
0!
0%
#674645000000
1!
1%
#674650000000
0!
0%
#674655000000
1!
1%
#674660000000
0!
0%
#674665000000
1!
1%
#674670000000
0!
0%
#674675000000
1!
1%
#674680000000
0!
0%
#674685000000
1!
1%
#674690000000
0!
0%
#674695000000
1!
1%
#674700000000
0!
0%
#674705000000
1!
1%
#674710000000
0!
0%
#674715000000
1!
1%
#674720000000
0!
0%
#674725000000
1!
1%
#674730000000
0!
0%
#674735000000
1!
1%
#674740000000
0!
0%
#674745000000
1!
1%
#674750000000
0!
0%
#674755000000
1!
1%
#674760000000
0!
0%
#674765000000
1!
1%
#674770000000
0!
0%
#674775000000
1!
1%
#674780000000
0!
0%
#674785000000
1!
1%
#674790000000
0!
0%
#674795000000
1!
1%
#674800000000
0!
0%
#674805000000
1!
1%
#674810000000
0!
0%
#674815000000
1!
1%
#674820000000
0!
0%
#674825000000
1!
1%
#674830000000
0!
0%
#674835000000
1!
1%
#674840000000
0!
0%
#674845000000
1!
1%
#674850000000
0!
0%
#674855000000
1!
1%
#674860000000
0!
0%
#674865000000
1!
1%
#674870000000
0!
0%
#674875000000
1!
1%
#674880000000
0!
0%
#674885000000
1!
1%
#674890000000
0!
0%
#674895000000
1!
1%
#674900000000
0!
0%
#674905000000
1!
1%
#674910000000
0!
0%
#674915000000
1!
1%
#674920000000
0!
0%
#674925000000
1!
1%
#674930000000
0!
0%
#674935000000
1!
1%
#674940000000
0!
0%
#674945000000
1!
1%
#674950000000
0!
0%
#674955000000
1!
1%
#674960000000
0!
0%
#674965000000
1!
1%
#674970000000
0!
0%
#674975000000
1!
1%
#674980000000
0!
0%
#674985000000
1!
1%
#674990000000
0!
0%
#674995000000
1!
1%
#675000000000
0!
0%
#675005000000
1!
1%
#675010000000
0!
0%
#675015000000
1!
1%
#675020000000
0!
0%
#675025000000
1!
1%
#675030000000
0!
0%
#675035000000
1!
1%
#675040000000
0!
0%
#675045000000
1!
1%
#675050000000
0!
0%
#675055000000
1!
1%
#675060000000
0!
0%
#675065000000
1!
1%
#675070000000
0!
0%
#675075000000
1!
1%
#675080000000
0!
0%
#675085000000
1!
1%
#675090000000
0!
0%
#675095000000
1!
1%
#675100000000
0!
0%
#675105000000
1!
1%
#675110000000
0!
0%
#675115000000
1!
1%
#675120000000
0!
0%
#675125000000
1!
1%
#675130000000
0!
0%
#675135000000
1!
1%
#675140000000
0!
0%
#675145000000
1!
1%
#675150000000
0!
0%
#675155000000
1!
1%
#675160000000
0!
0%
#675165000000
1!
1%
#675170000000
0!
0%
#675175000000
1!
1%
#675180000000
0!
0%
#675185000000
1!
1%
#675190000000
0!
0%
#675195000000
1!
1%
#675200000000
0!
0%
#675205000000
1!
1%
#675210000000
0!
0%
#675215000000
1!
1%
#675220000000
0!
0%
#675225000000
1!
1%
#675230000000
0!
0%
#675235000000
1!
1%
#675240000000
0!
0%
#675245000000
1!
1%
#675250000000
0!
0%
#675255000000
1!
1%
#675260000000
0!
0%
#675265000000
1!
1%
#675270000000
0!
0%
#675275000000
1!
1%
#675280000000
0!
0%
#675285000000
1!
1%
#675290000000
0!
0%
#675295000000
1!
1%
#675300000000
0!
0%
#675305000000
1!
1%
#675310000000
0!
0%
#675315000000
1!
1%
#675320000000
0!
0%
#675325000000
1!
1%
#675330000000
0!
0%
#675335000000
1!
1%
#675340000000
0!
0%
#675345000000
1!
1%
#675350000000
0!
0%
#675355000000
1!
1%
#675360000000
0!
0%
#675365000000
1!
1%
#675370000000
0!
0%
#675375000000
1!
1%
#675380000000
0!
0%
#675385000000
1!
1%
#675390000000
0!
0%
#675395000000
1!
1%
#675400000000
0!
0%
#675405000000
1!
1%
#675410000000
0!
0%
#675415000000
1!
1%
#675420000000
0!
0%
#675425000000
1!
1%
#675430000000
0!
0%
#675435000000
1!
1%
#675440000000
0!
0%
#675445000000
1!
1%
#675450000000
0!
0%
#675455000000
1!
1%
#675460000000
0!
0%
#675465000000
1!
1%
#675470000000
0!
0%
#675475000000
1!
1%
#675480000000
0!
0%
#675485000000
1!
1%
#675490000000
0!
0%
#675495000000
1!
1%
#675500000000
0!
0%
#675505000000
1!
1%
#675510000000
0!
0%
#675515000000
1!
1%
#675520000000
0!
0%
#675525000000
1!
1%
#675530000000
0!
0%
#675535000000
1!
1%
#675540000000
0!
0%
#675545000000
1!
1%
#675550000000
0!
0%
#675555000000
1!
1%
#675560000000
0!
0%
#675565000000
1!
1%
#675570000000
0!
0%
#675575000000
1!
1%
#675580000000
0!
0%
#675585000000
1!
1%
#675590000000
0!
0%
#675595000000
1!
1%
#675600000000
0!
0%
#675605000000
1!
1%
#675610000000
0!
0%
#675615000000
1!
1%
#675620000000
0!
0%
#675625000000
1!
1%
#675630000000
0!
0%
#675635000000
1!
1%
#675640000000
0!
0%
#675645000000
1!
1%
#675650000000
0!
0%
#675655000000
1!
1%
#675660000000
0!
0%
#675665000000
1!
1%
#675670000000
0!
0%
#675675000000
1!
1%
#675680000000
0!
0%
#675685000000
1!
1%
#675690000000
0!
0%
#675695000000
1!
1%
#675700000000
0!
0%
#675705000000
1!
1%
#675710000000
0!
0%
#675715000000
1!
1%
#675720000000
0!
0%
#675725000000
1!
1%
#675730000000
0!
0%
#675735000000
1!
1%
#675740000000
0!
0%
#675745000000
1!
1%
#675750000000
0!
0%
#675755000000
1!
1%
#675760000000
0!
0%
#675765000000
1!
1%
#675770000000
0!
0%
#675775000000
1!
1%
#675780000000
0!
0%
#675785000000
1!
1%
#675790000000
0!
0%
#675795000000
1!
1%
#675800000000
0!
0%
#675805000000
1!
1%
#675810000000
0!
0%
#675815000000
1!
1%
#675820000000
0!
0%
#675825000000
1!
1%
#675830000000
0!
0%
#675835000000
1!
1%
#675840000000
0!
0%
#675845000000
1!
1%
#675850000000
0!
0%
#675855000000
1!
1%
#675860000000
0!
0%
#675865000000
1!
1%
#675870000000
0!
0%
#675875000000
1!
1%
#675880000000
0!
0%
#675885000000
1!
1%
#675890000000
0!
0%
#675895000000
1!
1%
#675900000000
0!
0%
#675905000000
1!
1%
#675910000000
0!
0%
#675915000000
1!
1%
#675920000000
0!
0%
#675925000000
1!
1%
#675930000000
0!
0%
#675935000000
1!
1%
#675940000000
0!
0%
#675945000000
1!
1%
#675950000000
0!
0%
#675955000000
1!
1%
#675960000000
0!
0%
#675965000000
1!
1%
#675970000000
0!
0%
#675975000000
1!
1%
#675980000000
0!
0%
#675985000000
1!
1%
#675990000000
0!
0%
#675995000000
1!
1%
#676000000000
0!
0%
#676005000000
1!
1%
#676010000000
0!
0%
#676015000000
1!
1%
#676020000000
0!
0%
#676025000000
1!
1%
#676030000000
0!
0%
#676035000000
1!
1%
#676040000000
0!
0%
#676045000000
1!
1%
#676050000000
0!
0%
#676055000000
1!
1%
#676060000000
0!
0%
#676065000000
1!
1%
#676070000000
0!
0%
#676075000000
1!
1%
#676080000000
0!
0%
#676085000000
1!
1%
#676090000000
0!
0%
#676095000000
1!
1%
#676100000000
0!
0%
#676105000000
1!
1%
#676110000000
0!
0%
#676115000000
1!
1%
#676120000000
0!
0%
#676125000000
1!
1%
#676130000000
0!
0%
#676135000000
1!
1%
#676140000000
0!
0%
#676145000000
1!
1%
#676150000000
0!
0%
#676155000000
1!
1%
#676160000000
0!
0%
#676165000000
1!
1%
#676170000000
0!
0%
#676175000000
1!
1%
#676180000000
0!
0%
#676185000000
1!
1%
#676190000000
0!
0%
#676195000000
1!
1%
#676200000000
0!
0%
#676205000000
1!
1%
#676210000000
0!
0%
#676215000000
1!
1%
#676220000000
0!
0%
#676225000000
1!
1%
#676230000000
0!
0%
#676235000000
1!
1%
#676240000000
0!
0%
#676245000000
1!
1%
#676250000000
0!
0%
#676255000000
1!
1%
#676260000000
0!
0%
#676265000000
1!
1%
#676270000000
0!
0%
#676275000000
1!
1%
#676280000000
0!
0%
#676285000000
1!
1%
#676290000000
0!
0%
#676295000000
1!
1%
#676300000000
0!
0%
#676305000000
1!
1%
#676310000000
0!
0%
#676315000000
1!
1%
#676320000000
0!
0%
#676325000000
1!
1%
#676330000000
0!
0%
#676335000000
1!
1%
#676340000000
0!
0%
#676345000000
1!
1%
#676350000000
0!
0%
#676355000000
1!
1%
#676360000000
0!
0%
#676365000000
1!
1%
#676370000000
0!
0%
#676375000000
1!
1%
#676380000000
0!
0%
#676385000000
1!
1%
#676390000000
0!
0%
#676395000000
1!
1%
#676400000000
0!
0%
#676405000000
1!
1%
#676410000000
0!
0%
#676415000000
1!
1%
#676420000000
0!
0%
#676425000000
1!
1%
#676430000000
0!
0%
#676435000000
1!
1%
#676440000000
0!
0%
#676445000000
1!
1%
#676450000000
0!
0%
#676455000000
1!
1%
#676460000000
0!
0%
#676465000000
1!
1%
#676470000000
0!
0%
#676475000000
1!
1%
#676480000000
0!
0%
#676485000000
1!
1%
#676490000000
0!
0%
#676495000000
1!
1%
#676500000000
0!
0%
#676505000000
1!
1%
#676510000000
0!
0%
#676515000000
1!
1%
#676520000000
0!
0%
#676525000000
1!
1%
#676530000000
0!
0%
#676535000000
1!
1%
#676540000000
0!
0%
#676545000000
1!
1%
#676550000000
0!
0%
#676555000000
1!
1%
#676560000000
0!
0%
#676565000000
1!
1%
#676570000000
0!
0%
#676575000000
1!
1%
#676580000000
0!
0%
#676585000000
1!
1%
#676590000000
0!
0%
#676595000000
1!
1%
#676600000000
0!
0%
#676605000000
1!
1%
#676610000000
0!
0%
#676615000000
1!
1%
#676620000000
0!
0%
#676625000000
1!
1%
#676630000000
0!
0%
#676635000000
1!
1%
#676640000000
0!
0%
#676645000000
1!
1%
#676650000000
0!
0%
#676655000000
1!
1%
#676660000000
0!
0%
#676665000000
1!
1%
#676670000000
0!
0%
#676675000000
1!
1%
#676680000000
0!
0%
#676685000000
1!
1%
#676690000000
0!
0%
#676695000000
1!
1%
#676700000000
0!
0%
#676705000000
1!
1%
#676710000000
0!
0%
#676715000000
1!
1%
#676720000000
0!
0%
#676725000000
1!
1%
#676730000000
0!
0%
#676735000000
1!
1%
#676740000000
0!
0%
#676745000000
1!
1%
#676750000000
0!
0%
#676755000000
1!
1%
#676760000000
0!
0%
#676765000000
1!
1%
#676770000000
0!
0%
#676775000000
1!
1%
#676780000000
0!
0%
#676785000000
1!
1%
#676790000000
0!
0%
#676795000000
1!
1%
#676800000000
0!
0%
#676805000000
1!
1%
#676810000000
0!
0%
#676815000000
1!
1%
#676820000000
0!
0%
#676825000000
1!
1%
#676830000000
0!
0%
#676835000000
1!
1%
#676840000000
0!
0%
#676845000000
1!
1%
#676850000000
0!
0%
#676855000000
1!
1%
#676860000000
0!
0%
#676865000000
1!
1%
#676870000000
0!
0%
#676875000000
1!
1%
#676880000000
0!
0%
#676885000000
1!
1%
#676890000000
0!
0%
#676895000000
1!
1%
#676900000000
0!
0%
#676905000000
1!
1%
#676910000000
0!
0%
#676915000000
1!
1%
#676920000000
0!
0%
#676925000000
1!
1%
#676930000000
0!
0%
#676935000000
1!
1%
#676940000000
0!
0%
#676945000000
1!
1%
#676950000000
0!
0%
#676955000000
1!
1%
#676960000000
0!
0%
#676965000000
1!
1%
#676970000000
0!
0%
#676975000000
1!
1%
#676980000000
0!
0%
#676985000000
1!
1%
#676990000000
0!
0%
#676995000000
1!
1%
#677000000000
0!
0%
#677005000000
1!
1%
#677010000000
0!
0%
#677015000000
1!
1%
#677020000000
0!
0%
#677025000000
1!
1%
#677030000000
0!
0%
#677035000000
1!
1%
#677040000000
0!
0%
#677045000000
1!
1%
#677050000000
0!
0%
#677055000000
1!
1%
#677060000000
0!
0%
#677065000000
1!
1%
#677070000000
0!
0%
#677075000000
1!
1%
#677080000000
0!
0%
#677085000000
1!
1%
#677090000000
0!
0%
#677095000000
1!
1%
#677100000000
0!
0%
#677105000000
1!
1%
#677110000000
0!
0%
#677115000000
1!
1%
#677120000000
0!
0%
#677125000000
1!
1%
#677130000000
0!
0%
#677135000000
1!
1%
#677140000000
0!
0%
#677145000000
1!
1%
#677150000000
0!
0%
#677155000000
1!
1%
#677160000000
0!
0%
#677165000000
1!
1%
#677170000000
0!
0%
#677175000000
1!
1%
#677180000000
0!
0%
#677185000000
1!
1%
#677190000000
0!
0%
#677195000000
1!
1%
#677200000000
0!
0%
#677205000000
1!
1%
#677210000000
0!
0%
#677215000000
1!
1%
#677220000000
0!
0%
#677225000000
1!
1%
#677230000000
0!
0%
#677235000000
1!
1%
#677240000000
0!
0%
#677245000000
1!
1%
#677250000000
0!
0%
#677255000000
1!
1%
#677260000000
0!
0%
#677265000000
1!
1%
#677270000000
0!
0%
#677275000000
1!
1%
#677280000000
0!
0%
#677285000000
1!
1%
#677290000000
0!
0%
#677295000000
1!
1%
#677300000000
0!
0%
#677305000000
1!
1%
#677310000000
0!
0%
#677315000000
1!
1%
#677320000000
0!
0%
#677325000000
1!
1%
#677330000000
0!
0%
#677335000000
1!
1%
#677340000000
0!
0%
#677345000000
1!
1%
#677350000000
0!
0%
#677355000000
1!
1%
#677360000000
0!
0%
#677365000000
1!
1%
#677370000000
0!
0%
#677375000000
1!
1%
#677380000000
0!
0%
#677385000000
1!
1%
#677390000000
0!
0%
#677395000000
1!
1%
#677400000000
0!
0%
#677405000000
1!
1%
#677410000000
0!
0%
#677415000000
1!
1%
#677420000000
0!
0%
#677425000000
1!
1%
#677430000000
0!
0%
#677435000000
1!
1%
#677440000000
0!
0%
#677445000000
1!
1%
#677450000000
0!
0%
#677455000000
1!
1%
#677460000000
0!
0%
#677465000000
1!
1%
#677470000000
0!
0%
#677475000000
1!
1%
#677480000000
0!
0%
#677485000000
1!
1%
#677490000000
0!
0%
#677495000000
1!
1%
#677500000000
0!
0%
#677505000000
1!
1%
#677510000000
0!
0%
#677515000000
1!
1%
#677520000000
0!
0%
#677525000000
1!
1%
#677530000000
0!
0%
#677535000000
1!
1%
#677540000000
0!
0%
#677545000000
1!
1%
#677550000000
0!
0%
#677555000000
1!
1%
#677560000000
0!
0%
#677565000000
1!
1%
#677570000000
0!
0%
#677575000000
1!
1%
#677580000000
0!
0%
#677585000000
1!
1%
#677590000000
0!
0%
#677595000000
1!
1%
#677600000000
0!
0%
#677605000000
1!
1%
#677610000000
0!
0%
#677615000000
1!
1%
#677620000000
0!
0%
#677625000000
1!
1%
#677630000000
0!
0%
#677635000000
1!
1%
#677640000000
0!
0%
#677645000000
1!
1%
#677650000000
0!
0%
#677655000000
1!
1%
#677660000000
0!
0%
#677665000000
1!
1%
#677670000000
0!
0%
#677675000000
1!
1%
#677680000000
0!
0%
#677685000000
1!
1%
#677690000000
0!
0%
#677695000000
1!
1%
#677700000000
0!
0%
#677705000000
1!
1%
#677710000000
0!
0%
#677715000000
1!
1%
#677720000000
0!
0%
#677725000000
1!
1%
#677730000000
0!
0%
#677735000000
1!
1%
#677740000000
0!
0%
#677745000000
1!
1%
#677750000000
0!
0%
#677755000000
1!
1%
#677760000000
0!
0%
#677765000000
1!
1%
#677770000000
0!
0%
#677775000000
1!
1%
#677780000000
0!
0%
#677785000000
1!
1%
#677790000000
0!
0%
#677795000000
1!
1%
#677800000000
0!
0%
#677805000000
1!
1%
#677810000000
0!
0%
#677815000000
1!
1%
#677820000000
0!
0%
#677825000000
1!
1%
#677830000000
0!
0%
#677835000000
1!
1%
#677840000000
0!
0%
#677845000000
1!
1%
#677850000000
0!
0%
#677855000000
1!
1%
#677860000000
0!
0%
#677865000000
1!
1%
#677870000000
0!
0%
#677875000000
1!
1%
#677880000000
0!
0%
#677885000000
1!
1%
#677890000000
0!
0%
#677895000000
1!
1%
#677900000000
0!
0%
#677905000000
1!
1%
#677910000000
0!
0%
#677915000000
1!
1%
#677920000000
0!
0%
#677925000000
1!
1%
#677930000000
0!
0%
#677935000000
1!
1%
#677940000000
0!
0%
#677945000000
1!
1%
#677950000000
0!
0%
#677955000000
1!
1%
#677960000000
0!
0%
#677965000000
1!
1%
#677970000000
0!
0%
#677975000000
1!
1%
#677980000000
0!
0%
#677985000000
1!
1%
#677990000000
0!
0%
#677995000000
1!
1%
#678000000000
0!
0%
#678005000000
1!
1%
#678010000000
0!
0%
#678015000000
1!
1%
#678020000000
0!
0%
#678025000000
1!
1%
#678030000000
0!
0%
#678035000000
1!
1%
#678040000000
0!
0%
#678045000000
1!
1%
#678050000000
0!
0%
#678055000000
1!
1%
#678060000000
0!
0%
#678065000000
1!
1%
#678070000000
0!
0%
#678075000000
1!
1%
#678080000000
0!
0%
#678085000000
1!
1%
#678090000000
0!
0%
#678095000000
1!
1%
#678100000000
0!
0%
#678105000000
1!
1%
#678110000000
0!
0%
#678115000000
1!
1%
#678120000000
0!
0%
#678125000000
1!
1%
#678130000000
0!
0%
#678135000000
1!
1%
#678140000000
0!
0%
#678145000000
1!
1%
#678150000000
0!
0%
#678155000000
1!
1%
#678160000000
0!
0%
#678165000000
1!
1%
#678170000000
0!
0%
#678175000000
1!
1%
#678180000000
0!
0%
#678185000000
1!
1%
#678190000000
0!
0%
#678195000000
1!
1%
#678200000000
0!
0%
#678205000000
1!
1%
#678210000000
0!
0%
#678215000000
1!
1%
#678220000000
0!
0%
#678225000000
1!
1%
#678230000000
0!
0%
#678235000000
1!
1%
#678240000000
0!
0%
#678245000000
1!
1%
#678250000000
0!
0%
#678255000000
1!
1%
#678260000000
0!
0%
#678265000000
1!
1%
#678270000000
0!
0%
#678275000000
1!
1%
#678280000000
0!
0%
#678285000000
1!
1%
#678290000000
0!
0%
#678295000000
1!
1%
#678300000000
0!
0%
#678305000000
1!
1%
#678310000000
0!
0%
#678315000000
1!
1%
#678320000000
0!
0%
#678325000000
1!
1%
#678330000000
0!
0%
#678335000000
1!
1%
#678340000000
0!
0%
#678345000000
1!
1%
#678350000000
0!
0%
#678355000000
1!
1%
#678360000000
0!
0%
#678365000000
1!
1%
#678370000000
0!
0%
#678375000000
1!
1%
#678380000000
0!
0%
#678385000000
1!
1%
#678390000000
0!
0%
#678395000000
1!
1%
#678400000000
0!
0%
#678405000000
1!
1%
#678410000000
0!
0%
#678415000000
1!
1%
#678420000000
0!
0%
#678425000000
1!
1%
#678430000000
0!
0%
#678435000000
1!
1%
#678440000000
0!
0%
#678445000000
1!
1%
#678450000000
0!
0%
#678455000000
1!
1%
#678460000000
0!
0%
#678465000000
1!
1%
#678470000000
0!
0%
#678475000000
1!
1%
#678480000000
0!
0%
#678485000000
1!
1%
#678490000000
0!
0%
#678495000000
1!
1%
#678500000000
0!
0%
#678505000000
1!
1%
#678510000000
0!
0%
#678515000000
1!
1%
#678520000000
0!
0%
#678525000000
1!
1%
#678530000000
0!
0%
#678535000000
1!
1%
#678540000000
0!
0%
#678545000000
1!
1%
#678550000000
0!
0%
#678555000000
1!
1%
#678560000000
0!
0%
#678565000000
1!
1%
#678570000000
0!
0%
#678575000000
1!
1%
#678580000000
0!
0%
#678585000000
1!
1%
#678590000000
0!
0%
#678595000000
1!
1%
#678600000000
0!
0%
#678605000000
1!
1%
#678610000000
0!
0%
#678615000000
1!
1%
#678620000000
0!
0%
#678625000000
1!
1%
#678630000000
0!
0%
#678635000000
1!
1%
#678640000000
0!
0%
#678645000000
1!
1%
#678650000000
0!
0%
#678655000000
1!
1%
#678660000000
0!
0%
#678665000000
1!
1%
#678670000000
0!
0%
#678675000000
1!
1%
#678680000000
0!
0%
#678685000000
1!
1%
#678690000000
0!
0%
#678695000000
1!
1%
#678700000000
0!
0%
#678705000000
1!
1%
#678710000000
0!
0%
#678715000000
1!
1%
#678720000000
0!
0%
#678725000000
1!
1%
#678730000000
0!
0%
#678735000000
1!
1%
#678740000000
0!
0%
#678745000000
1!
1%
#678750000000
0!
0%
#678755000000
1!
1%
#678760000000
0!
0%
#678765000000
1!
1%
#678770000000
0!
0%
#678775000000
1!
1%
#678780000000
0!
0%
#678785000000
1!
1%
#678790000000
0!
0%
#678795000000
1!
1%
#678800000000
0!
0%
#678805000000
1!
1%
#678810000000
0!
0%
#678815000000
1!
1%
#678820000000
0!
0%
#678825000000
1!
1%
#678830000000
0!
0%
#678835000000
1!
1%
#678840000000
0!
0%
#678845000000
1!
1%
#678850000000
0!
0%
#678855000000
1!
1%
#678860000000
0!
0%
#678865000000
1!
1%
#678870000000
0!
0%
#678875000000
1!
1%
#678880000000
0!
0%
#678885000000
1!
1%
#678890000000
0!
0%
#678895000000
1!
1%
#678900000000
0!
0%
#678905000000
1!
1%
#678910000000
0!
0%
#678915000000
1!
1%
#678920000000
0!
0%
#678925000000
1!
1%
#678930000000
0!
0%
#678935000000
1!
1%
#678940000000
0!
0%
#678945000000
1!
1%
#678950000000
0!
0%
#678955000000
1!
1%
#678960000000
0!
0%
#678965000000
1!
1%
#678970000000
0!
0%
#678975000000
1!
1%
#678980000000
0!
0%
#678985000000
1!
1%
#678990000000
0!
0%
#678995000000
1!
1%
#679000000000
0!
0%
#679005000000
1!
1%
#679010000000
0!
0%
#679015000000
1!
1%
#679020000000
0!
0%
#679025000000
1!
1%
#679030000000
0!
0%
#679035000000
1!
1%
#679040000000
0!
0%
#679045000000
1!
1%
#679050000000
0!
0%
#679055000000
1!
1%
#679060000000
0!
0%
#679065000000
1!
1%
#679070000000
0!
0%
#679075000000
1!
1%
#679080000000
0!
0%
#679085000000
1!
1%
#679090000000
0!
0%
#679095000000
1!
1%
#679100000000
0!
0%
#679105000000
1!
1%
#679110000000
0!
0%
#679115000000
1!
1%
#679120000000
0!
0%
#679125000000
1!
1%
#679130000000
0!
0%
#679135000000
1!
1%
#679140000000
0!
0%
#679145000000
1!
1%
#679150000000
0!
0%
#679155000000
1!
1%
#679160000000
0!
0%
#679165000000
1!
1%
#679170000000
0!
0%
#679175000000
1!
1%
#679180000000
0!
0%
#679185000000
1!
1%
#679190000000
0!
0%
#679195000000
1!
1%
#679200000000
0!
0%
#679205000000
1!
1%
#679210000000
0!
0%
#679215000000
1!
1%
#679220000000
0!
0%
#679225000000
1!
1%
#679230000000
0!
0%
#679235000000
1!
1%
#679240000000
0!
0%
#679245000000
1!
1%
#679250000000
0!
0%
#679255000000
1!
1%
#679260000000
0!
0%
#679265000000
1!
1%
#679270000000
0!
0%
#679275000000
1!
1%
#679280000000
0!
0%
#679285000000
1!
1%
#679290000000
0!
0%
#679295000000
1!
1%
#679300000000
0!
0%
#679305000000
1!
1%
#679310000000
0!
0%
#679315000000
1!
1%
#679320000000
0!
0%
#679325000000
1!
1%
#679330000000
0!
0%
#679335000000
1!
1%
#679340000000
0!
0%
#679345000000
1!
1%
#679350000000
0!
0%
#679355000000
1!
1%
#679360000000
0!
0%
#679365000000
1!
1%
#679370000000
0!
0%
#679375000000
1!
1%
#679380000000
0!
0%
#679385000000
1!
1%
#679390000000
0!
0%
#679395000000
1!
1%
#679400000000
0!
0%
#679405000000
1!
1%
#679410000000
0!
0%
#679415000000
1!
1%
#679420000000
0!
0%
#679425000000
1!
1%
#679430000000
0!
0%
#679435000000
1!
1%
#679440000000
0!
0%
#679445000000
1!
1%
#679450000000
0!
0%
#679455000000
1!
1%
#679460000000
0!
0%
#679465000000
1!
1%
#679470000000
0!
0%
#679475000000
1!
1%
#679480000000
0!
0%
#679485000000
1!
1%
#679490000000
0!
0%
#679495000000
1!
1%
#679500000000
0!
0%
#679505000000
1!
1%
#679510000000
0!
0%
#679515000000
1!
1%
#679520000000
0!
0%
#679525000000
1!
1%
#679530000000
0!
0%
#679535000000
1!
1%
#679540000000
0!
0%
#679545000000
1!
1%
#679550000000
0!
0%
#679555000000
1!
1%
#679560000000
0!
0%
#679565000000
1!
1%
#679570000000
0!
0%
#679575000000
1!
1%
#679580000000
0!
0%
#679585000000
1!
1%
#679590000000
0!
0%
#679595000000
1!
1%
#679600000000
0!
0%
#679605000000
1!
1%
#679610000000
0!
0%
#679615000000
1!
1%
#679620000000
0!
0%
#679625000000
1!
1%
#679630000000
0!
0%
#679635000000
1!
1%
#679640000000
0!
0%
#679645000000
1!
1%
#679650000000
0!
0%
#679655000000
1!
1%
#679660000000
0!
0%
#679665000000
1!
1%
#679670000000
0!
0%
#679675000000
1!
1%
#679680000000
0!
0%
#679685000000
1!
1%
#679690000000
0!
0%
#679695000000
1!
1%
#679700000000
0!
0%
#679705000000
1!
1%
#679710000000
0!
0%
#679715000000
1!
1%
#679720000000
0!
0%
#679725000000
1!
1%
#679730000000
0!
0%
#679735000000
1!
1%
#679740000000
0!
0%
#679745000000
1!
1%
#679750000000
0!
0%
#679755000000
1!
1%
#679760000000
0!
0%
#679765000000
1!
1%
#679770000000
0!
0%
#679775000000
1!
1%
#679780000000
0!
0%
#679785000000
1!
1%
#679790000000
0!
0%
#679795000000
1!
1%
#679800000000
0!
0%
#679805000000
1!
1%
#679810000000
0!
0%
#679815000000
1!
1%
#679820000000
0!
0%
#679825000000
1!
1%
#679830000000
0!
0%
#679835000000
1!
1%
#679840000000
0!
0%
#679845000000
1!
1%
#679850000000
0!
0%
#679855000000
1!
1%
#679860000000
0!
0%
#679865000000
1!
1%
#679870000000
0!
0%
#679875000000
1!
1%
#679880000000
0!
0%
#679885000000
1!
1%
#679890000000
0!
0%
#679895000000
1!
1%
#679900000000
0!
0%
#679905000000
1!
1%
#679910000000
0!
0%
#679915000000
1!
1%
#679920000000
0!
0%
#679925000000
1!
1%
#679930000000
0!
0%
#679935000000
1!
1%
#679940000000
0!
0%
#679945000000
1!
1%
#679950000000
0!
0%
#679955000000
1!
1%
#679960000000
0!
0%
#679965000000
1!
1%
#679970000000
0!
0%
#679975000000
1!
1%
#679980000000
0!
0%
#679985000000
1!
1%
#679990000000
0!
0%
#679995000000
1!
1%
#680000000000
0!
0%
#680005000000
1!
1%
#680010000000
0!
0%
#680015000000
1!
1%
#680020000000
0!
0%
#680025000000
1!
1%
#680030000000
0!
0%
#680035000000
1!
1%
#680040000000
0!
0%
#680045000000
1!
1%
#680050000000
0!
0%
#680055000000
1!
1%
#680060000000
0!
0%
#680065000000
1!
1%
#680070000000
0!
0%
#680075000000
1!
1%
#680080000000
0!
0%
#680085000000
1!
1%
#680090000000
0!
0%
#680095000000
1!
1%
#680100000000
0!
0%
#680105000000
1!
1%
#680110000000
0!
0%
#680115000000
1!
1%
#680120000000
0!
0%
#680125000000
1!
1%
#680130000000
0!
0%
#680135000000
1!
1%
#680140000000
0!
0%
#680145000000
1!
1%
#680150000000
0!
0%
#680155000000
1!
1%
#680160000000
0!
0%
#680165000000
1!
1%
#680170000000
0!
0%
#680175000000
1!
1%
#680180000000
0!
0%
#680185000000
1!
1%
#680190000000
0!
0%
#680195000000
1!
1%
#680200000000
0!
0%
#680205000000
1!
1%
#680210000000
0!
0%
#680215000000
1!
1%
#680220000000
0!
0%
#680225000000
1!
1%
#680230000000
0!
0%
#680235000000
1!
1%
#680240000000
0!
0%
#680245000000
1!
1%
#680250000000
0!
0%
#680255000000
1!
1%
#680260000000
0!
0%
#680265000000
1!
1%
#680270000000
0!
0%
#680275000000
1!
1%
#680280000000
0!
0%
#680285000000
1!
1%
#680290000000
0!
0%
#680295000000
1!
1%
#680300000000
0!
0%
#680305000000
1!
1%
#680310000000
0!
0%
#680315000000
1!
1%
#680320000000
0!
0%
#680325000000
1!
1%
#680330000000
0!
0%
#680335000000
1!
1%
#680340000000
0!
0%
#680345000000
1!
1%
#680350000000
0!
0%
#680355000000
1!
1%
#680360000000
0!
0%
#680365000000
1!
1%
#680370000000
0!
0%
#680375000000
1!
1%
#680380000000
0!
0%
#680385000000
1!
1%
#680390000000
0!
0%
#680395000000
1!
1%
#680400000000
0!
0%
#680405000000
1!
1%
#680410000000
0!
0%
#680415000000
1!
1%
#680420000000
0!
0%
#680425000000
1!
1%
#680430000000
0!
0%
#680435000000
1!
1%
#680440000000
0!
0%
#680445000000
1!
1%
#680450000000
0!
0%
#680455000000
1!
1%
#680460000000
0!
0%
#680465000000
1!
1%
#680470000000
0!
0%
#680475000000
1!
1%
#680480000000
0!
0%
#680485000000
1!
1%
#680490000000
0!
0%
#680495000000
1!
1%
#680500000000
0!
0%
#680505000000
1!
1%
#680510000000
0!
0%
#680515000000
1!
1%
#680520000000
0!
0%
#680525000000
1!
1%
#680530000000
0!
0%
#680535000000
1!
1%
#680540000000
0!
0%
#680545000000
1!
1%
#680550000000
0!
0%
#680555000000
1!
1%
#680560000000
0!
0%
#680565000000
1!
1%
#680570000000
0!
0%
#680575000000
1!
1%
#680580000000
0!
0%
#680585000000
1!
1%
#680590000000
0!
0%
#680595000000
1!
1%
#680600000000
0!
0%
#680605000000
1!
1%
#680610000000
0!
0%
#680615000000
1!
1%
#680620000000
0!
0%
#680625000000
1!
1%
#680630000000
0!
0%
#680635000000
1!
1%
#680640000000
0!
0%
#680645000000
1!
1%
#680650000000
0!
0%
#680655000000
1!
1%
#680660000000
0!
0%
#680665000000
1!
1%
#680670000000
0!
0%
#680675000000
1!
1%
#680680000000
0!
0%
#680685000000
1!
1%
#680690000000
0!
0%
#680695000000
1!
1%
#680700000000
0!
0%
#680705000000
1!
1%
#680710000000
0!
0%
#680715000000
1!
1%
#680720000000
0!
0%
#680725000000
1!
1%
#680730000000
0!
0%
#680735000000
1!
1%
#680740000000
0!
0%
#680745000000
1!
1%
#680750000000
0!
0%
#680755000000
1!
1%
#680760000000
0!
0%
#680765000000
1!
1%
#680770000000
0!
0%
#680775000000
1!
1%
#680780000000
0!
0%
#680785000000
1!
1%
#680790000000
0!
0%
#680795000000
1!
1%
#680800000000
0!
0%
#680805000000
1!
1%
#680810000000
0!
0%
#680815000000
1!
1%
#680820000000
0!
0%
#680825000000
1!
1%
#680830000000
0!
0%
#680835000000
1!
1%
#680840000000
0!
0%
#680845000000
1!
1%
#680850000000
0!
0%
#680855000000
1!
1%
#680860000000
0!
0%
#680865000000
1!
1%
#680870000000
0!
0%
#680875000000
1!
1%
#680880000000
0!
0%
#680885000000
1!
1%
#680890000000
0!
0%
#680895000000
1!
1%
#680900000000
0!
0%
#680905000000
1!
1%
#680910000000
0!
0%
#680915000000
1!
1%
#680920000000
0!
0%
#680925000000
1!
1%
#680930000000
0!
0%
#680935000000
1!
1%
#680940000000
0!
0%
#680945000000
1!
1%
#680950000000
0!
0%
#680955000000
1!
1%
#680960000000
0!
0%
#680965000000
1!
1%
#680970000000
0!
0%
#680975000000
1!
1%
#680980000000
0!
0%
#680985000000
1!
1%
#680990000000
0!
0%
#680995000000
1!
1%
#681000000000
0!
0%
#681005000000
1!
1%
#681010000000
0!
0%
#681015000000
1!
1%
#681020000000
0!
0%
#681025000000
1!
1%
#681030000000
0!
0%
#681035000000
1!
1%
#681040000000
0!
0%
#681045000000
1!
1%
#681050000000
0!
0%
#681055000000
1!
1%
#681060000000
0!
0%
#681065000000
1!
1%
#681070000000
0!
0%
#681075000000
1!
1%
#681080000000
0!
0%
#681085000000
1!
1%
#681090000000
0!
0%
#681095000000
1!
1%
#681100000000
0!
0%
#681105000000
1!
1%
#681110000000
0!
0%
#681115000000
1!
1%
#681120000000
0!
0%
#681125000000
1!
1%
#681130000000
0!
0%
#681135000000
1!
1%
#681140000000
0!
0%
#681145000000
1!
1%
#681150000000
0!
0%
#681155000000
1!
1%
#681160000000
0!
0%
#681165000000
1!
1%
#681170000000
0!
0%
#681175000000
1!
1%
#681180000000
0!
0%
#681185000000
1!
1%
#681190000000
0!
0%
#681195000000
1!
1%
#681200000000
0!
0%
#681205000000
1!
1%
#681210000000
0!
0%
#681215000000
1!
1%
#681220000000
0!
0%
#681225000000
1!
1%
#681230000000
0!
0%
#681235000000
1!
1%
#681240000000
0!
0%
#681245000000
1!
1%
#681250000000
0!
0%
#681255000000
1!
1%
#681260000000
0!
0%
#681265000000
1!
1%
#681270000000
0!
0%
#681275000000
1!
1%
#681280000000
0!
0%
#681285000000
1!
1%
#681290000000
0!
0%
#681295000000
1!
1%
#681300000000
0!
0%
#681305000000
1!
1%
#681310000000
0!
0%
#681315000000
1!
1%
#681320000000
0!
0%
#681325000000
1!
1%
#681330000000
0!
0%
#681335000000
1!
1%
#681340000000
0!
0%
#681345000000
1!
1%
#681350000000
0!
0%
#681355000000
1!
1%
#681360000000
0!
0%
#681365000000
1!
1%
#681370000000
0!
0%
#681375000000
1!
1%
#681380000000
0!
0%
#681385000000
1!
1%
#681390000000
0!
0%
#681395000000
1!
1%
#681400000000
0!
0%
#681405000000
1!
1%
#681410000000
0!
0%
#681415000000
1!
1%
#681420000000
0!
0%
#681425000000
1!
1%
#681430000000
0!
0%
#681435000000
1!
1%
#681440000000
0!
0%
#681445000000
1!
1%
#681450000000
0!
0%
#681455000000
1!
1%
#681460000000
0!
0%
#681465000000
1!
1%
#681470000000
0!
0%
#681475000000
1!
1%
#681480000000
0!
0%
#681485000000
1!
1%
#681490000000
0!
0%
#681495000000
1!
1%
#681500000000
0!
0%
#681505000000
1!
1%
#681510000000
0!
0%
#681515000000
1!
1%
#681520000000
0!
0%
#681525000000
1!
1%
#681530000000
0!
0%
#681535000000
1!
1%
#681540000000
0!
0%
#681545000000
1!
1%
#681550000000
0!
0%
#681555000000
1!
1%
#681560000000
0!
0%
#681565000000
1!
1%
#681570000000
0!
0%
#681575000000
1!
1%
#681580000000
0!
0%
#681585000000
1!
1%
#681590000000
0!
0%
#681595000000
1!
1%
#681600000000
0!
0%
#681605000000
1!
1%
#681610000000
0!
0%
#681615000000
1!
1%
#681620000000
0!
0%
#681625000000
1!
1%
#681630000000
0!
0%
#681635000000
1!
1%
#681640000000
0!
0%
#681645000000
1!
1%
#681650000000
0!
0%
#681655000000
1!
1%
#681660000000
0!
0%
#681665000000
1!
1%
#681670000000
0!
0%
#681675000000
1!
1%
#681680000000
0!
0%
#681685000000
1!
1%
#681690000000
0!
0%
#681695000000
1!
1%
#681700000000
0!
0%
#681705000000
1!
1%
#681710000000
0!
0%
#681715000000
1!
1%
#681720000000
0!
0%
#681725000000
1!
1%
#681730000000
0!
0%
#681735000000
1!
1%
#681740000000
0!
0%
#681745000000
1!
1%
#681750000000
0!
0%
#681755000000
1!
1%
#681760000000
0!
0%
#681765000000
1!
1%
#681770000000
0!
0%
#681775000000
1!
1%
#681780000000
0!
0%
#681785000000
1!
1%
#681790000000
0!
0%
#681795000000
1!
1%
#681800000000
0!
0%
#681805000000
1!
1%
#681810000000
0!
0%
#681815000000
1!
1%
#681820000000
0!
0%
#681825000000
1!
1%
#681830000000
0!
0%
#681835000000
1!
1%
#681840000000
0!
0%
#681845000000
1!
1%
#681850000000
0!
0%
#681855000000
1!
1%
#681860000000
0!
0%
#681865000000
1!
1%
#681870000000
0!
0%
#681875000000
1!
1%
#681880000000
0!
0%
#681885000000
1!
1%
#681890000000
0!
0%
#681895000000
1!
1%
#681900000000
0!
0%
#681905000000
1!
1%
#681910000000
0!
0%
#681915000000
1!
1%
#681920000000
0!
0%
#681925000000
1!
1%
#681930000000
0!
0%
#681935000000
1!
1%
#681940000000
0!
0%
#681945000000
1!
1%
#681950000000
0!
0%
#681955000000
1!
1%
#681960000000
0!
0%
#681965000000
1!
1%
#681970000000
0!
0%
#681975000000
1!
1%
#681980000000
0!
0%
#681985000000
1!
1%
#681990000000
0!
0%
#681995000000
1!
1%
#682000000000
0!
0%
#682005000000
1!
1%
#682010000000
0!
0%
#682015000000
1!
1%
#682020000000
0!
0%
#682025000000
1!
1%
#682030000000
0!
0%
#682035000000
1!
1%
#682040000000
0!
0%
#682045000000
1!
1%
#682050000000
0!
0%
#682055000000
1!
1%
#682060000000
0!
0%
#682065000000
1!
1%
#682070000000
0!
0%
#682075000000
1!
1%
#682080000000
0!
0%
#682085000000
1!
1%
#682090000000
0!
0%
#682095000000
1!
1%
#682100000000
0!
0%
#682105000000
1!
1%
#682110000000
0!
0%
#682115000000
1!
1%
#682120000000
0!
0%
#682125000000
1!
1%
#682130000000
0!
0%
#682135000000
1!
1%
#682140000000
0!
0%
#682145000000
1!
1%
#682150000000
0!
0%
#682155000000
1!
1%
#682160000000
0!
0%
#682165000000
1!
1%
#682170000000
0!
0%
#682175000000
1!
1%
#682180000000
0!
0%
#682185000000
1!
1%
#682190000000
0!
0%
#682195000000
1!
1%
#682200000000
0!
0%
#682205000000
1!
1%
#682210000000
0!
0%
#682215000000
1!
1%
#682220000000
0!
0%
#682225000000
1!
1%
#682230000000
0!
0%
#682235000000
1!
1%
#682240000000
0!
0%
#682245000000
1!
1%
#682250000000
0!
0%
#682255000000
1!
1%
#682260000000
0!
0%
#682265000000
1!
1%
#682270000000
0!
0%
#682275000000
1!
1%
#682280000000
0!
0%
#682285000000
1!
1%
#682290000000
0!
0%
#682295000000
1!
1%
#682300000000
0!
0%
#682305000000
1!
1%
#682310000000
0!
0%
#682315000000
1!
1%
#682320000000
0!
0%
#682325000000
1!
1%
#682330000000
0!
0%
#682335000000
1!
1%
#682340000000
0!
0%
#682345000000
1!
1%
#682350000000
0!
0%
#682355000000
1!
1%
#682360000000
0!
0%
#682365000000
1!
1%
#682370000000
0!
0%
#682375000000
1!
1%
#682380000000
0!
0%
#682385000000
1!
1%
#682390000000
0!
0%
#682395000000
1!
1%
#682400000000
0!
0%
#682405000000
1!
1%
#682410000000
0!
0%
#682415000000
1!
1%
#682420000000
0!
0%
#682425000000
1!
1%
#682430000000
0!
0%
#682435000000
1!
1%
#682440000000
0!
0%
#682445000000
1!
1%
#682450000000
0!
0%
#682455000000
1!
1%
#682460000000
0!
0%
#682465000000
1!
1%
#682470000000
0!
0%
#682475000000
1!
1%
#682480000000
0!
0%
#682485000000
1!
1%
#682490000000
0!
0%
#682495000000
1!
1%
#682500000000
0!
0%
#682505000000
1!
1%
#682510000000
0!
0%
#682515000000
1!
1%
#682520000000
0!
0%
#682525000000
1!
1%
#682530000000
0!
0%
#682535000000
1!
1%
#682540000000
0!
0%
#682545000000
1!
1%
#682550000000
0!
0%
#682555000000
1!
1%
#682560000000
0!
0%
#682565000000
1!
1%
#682570000000
0!
0%
#682575000000
1!
1%
#682580000000
0!
0%
#682585000000
1!
1%
#682590000000
0!
0%
#682595000000
1!
1%
#682600000000
0!
0%
#682605000000
1!
1%
#682610000000
0!
0%
#682615000000
1!
1%
#682620000000
0!
0%
#682625000000
1!
1%
#682630000000
0!
0%
#682635000000
1!
1%
#682640000000
0!
0%
#682645000000
1!
1%
#682650000000
0!
0%
#682655000000
1!
1%
#682660000000
0!
0%
#682665000000
1!
1%
#682670000000
0!
0%
#682675000000
1!
1%
#682680000000
0!
0%
#682685000000
1!
1%
#682690000000
0!
0%
#682695000000
1!
1%
#682700000000
0!
0%
#682705000000
1!
1%
#682710000000
0!
0%
#682715000000
1!
1%
#682720000000
0!
0%
#682725000000
1!
1%
#682730000000
0!
0%
#682735000000
1!
1%
#682740000000
0!
0%
#682745000000
1!
1%
#682750000000
0!
0%
#682755000000
1!
1%
#682760000000
0!
0%
#682765000000
1!
1%
#682770000000
0!
0%
#682775000000
1!
1%
#682780000000
0!
0%
#682785000000
1!
1%
#682790000000
0!
0%
#682795000000
1!
1%
#682800000000
0!
0%
#682805000000
1!
1%
#682810000000
0!
0%
#682815000000
1!
1%
#682820000000
0!
0%
#682825000000
1!
1%
#682830000000
0!
0%
#682835000000
1!
1%
#682840000000
0!
0%
#682845000000
1!
1%
#682850000000
0!
0%
#682855000000
1!
1%
#682860000000
0!
0%
#682865000000
1!
1%
#682870000000
0!
0%
#682875000000
1!
1%
#682880000000
0!
0%
#682885000000
1!
1%
#682890000000
0!
0%
#682895000000
1!
1%
#682900000000
0!
0%
#682905000000
1!
1%
#682910000000
0!
0%
#682915000000
1!
1%
#682920000000
0!
0%
#682925000000
1!
1%
#682930000000
0!
0%
#682935000000
1!
1%
#682940000000
0!
0%
#682945000000
1!
1%
#682950000000
0!
0%
#682955000000
1!
1%
#682960000000
0!
0%
#682965000000
1!
1%
#682970000000
0!
0%
#682975000000
1!
1%
#682980000000
0!
0%
#682985000000
1!
1%
#682990000000
0!
0%
#682995000000
1!
1%
#683000000000
0!
0%
#683005000000
1!
1%
#683010000000
0!
0%
#683015000000
1!
1%
#683020000000
0!
0%
#683025000000
1!
1%
#683030000000
0!
0%
#683035000000
1!
1%
#683040000000
0!
0%
#683045000000
1!
1%
#683050000000
0!
0%
#683055000000
1!
1%
#683060000000
0!
0%
#683065000000
1!
1%
#683070000000
0!
0%
#683075000000
1!
1%
#683080000000
0!
0%
#683085000000
1!
1%
#683090000000
0!
0%
#683095000000
1!
1%
#683100000000
0!
0%
#683105000000
1!
1%
#683110000000
0!
0%
#683115000000
1!
1%
#683120000000
0!
0%
#683125000000
1!
1%
#683130000000
0!
0%
#683135000000
1!
1%
#683140000000
0!
0%
#683145000000
1!
1%
#683150000000
0!
0%
#683155000000
1!
1%
#683160000000
0!
0%
#683165000000
1!
1%
#683170000000
0!
0%
#683175000000
1!
1%
#683180000000
0!
0%
#683185000000
1!
1%
#683190000000
0!
0%
#683195000000
1!
1%
#683200000000
0!
0%
#683205000000
1!
1%
#683210000000
0!
0%
#683215000000
1!
1%
#683220000000
0!
0%
#683225000000
1!
1%
#683230000000
0!
0%
#683235000000
1!
1%
#683240000000
0!
0%
#683245000000
1!
1%
#683250000000
0!
0%
#683255000000
1!
1%
#683260000000
0!
0%
#683265000000
1!
1%
#683270000000
0!
0%
#683275000000
1!
1%
#683280000000
0!
0%
#683285000000
1!
1%
#683290000000
0!
0%
#683295000000
1!
1%
#683300000000
0!
0%
#683305000000
1!
1%
#683310000000
0!
0%
#683315000000
1!
1%
#683320000000
0!
0%
#683325000000
1!
1%
#683330000000
0!
0%
#683335000000
1!
1%
#683340000000
0!
0%
#683345000000
1!
1%
#683350000000
0!
0%
#683355000000
1!
1%
#683360000000
0!
0%
#683365000000
1!
1%
#683370000000
0!
0%
#683375000000
1!
1%
#683380000000
0!
0%
#683385000000
1!
1%
#683390000000
0!
0%
#683395000000
1!
1%
#683400000000
0!
0%
#683405000000
1!
1%
#683410000000
0!
0%
#683415000000
1!
1%
#683420000000
0!
0%
#683425000000
1!
1%
#683430000000
0!
0%
#683435000000
1!
1%
#683440000000
0!
0%
#683445000000
1!
1%
#683450000000
0!
0%
#683455000000
1!
1%
#683460000000
0!
0%
#683465000000
1!
1%
#683470000000
0!
0%
#683475000000
1!
1%
#683480000000
0!
0%
#683485000000
1!
1%
#683490000000
0!
0%
#683495000000
1!
1%
#683500000000
0!
0%
#683505000000
1!
1%
#683510000000
0!
0%
#683515000000
1!
1%
#683520000000
0!
0%
#683525000000
1!
1%
#683530000000
0!
0%
#683535000000
1!
1%
#683540000000
0!
0%
#683545000000
1!
1%
#683550000000
0!
0%
#683555000000
1!
1%
#683560000000
0!
0%
#683565000000
1!
1%
#683570000000
0!
0%
#683575000000
1!
1%
#683580000000
0!
0%
#683585000000
1!
1%
#683590000000
0!
0%
#683595000000
1!
1%
#683600000000
0!
0%
#683605000000
1!
1%
#683610000000
0!
0%
#683615000000
1!
1%
#683620000000
0!
0%
#683625000000
1!
1%
#683630000000
0!
0%
#683635000000
1!
1%
#683640000000
0!
0%
#683645000000
1!
1%
#683650000000
0!
0%
#683655000000
1!
1%
#683660000000
0!
0%
#683665000000
1!
1%
#683670000000
0!
0%
#683675000000
1!
1%
#683680000000
0!
0%
#683685000000
1!
1%
#683690000000
0!
0%
#683695000000
1!
1%
#683700000000
0!
0%
#683705000000
1!
1%
#683710000000
0!
0%
#683715000000
1!
1%
#683720000000
0!
0%
#683725000000
1!
1%
#683730000000
0!
0%
#683735000000
1!
1%
#683740000000
0!
0%
#683745000000
1!
1%
#683750000000
0!
0%
#683755000000
1!
1%
#683760000000
0!
0%
#683765000000
1!
1%
#683770000000
0!
0%
#683775000000
1!
1%
#683780000000
0!
0%
#683785000000
1!
1%
#683790000000
0!
0%
#683795000000
1!
1%
#683800000000
0!
0%
#683805000000
1!
1%
#683810000000
0!
0%
#683815000000
1!
1%
#683820000000
0!
0%
#683825000000
1!
1%
#683830000000
0!
0%
#683835000000
1!
1%
#683840000000
0!
0%
#683845000000
1!
1%
#683850000000
0!
0%
#683855000000
1!
1%
#683860000000
0!
0%
#683865000000
1!
1%
#683870000000
0!
0%
#683875000000
1!
1%
#683880000000
0!
0%
#683885000000
1!
1%
#683890000000
0!
0%
#683895000000
1!
1%
#683900000000
0!
0%
#683905000000
1!
1%
#683910000000
0!
0%
#683915000000
1!
1%
#683920000000
0!
0%
#683925000000
1!
1%
#683930000000
0!
0%
#683935000000
1!
1%
#683940000000
0!
0%
#683945000000
1!
1%
#683950000000
0!
0%
#683955000000
1!
1%
#683960000000
0!
0%
#683965000000
1!
1%
#683970000000
0!
0%
#683975000000
1!
1%
#683980000000
0!
0%
#683985000000
1!
1%
#683990000000
0!
0%
#683995000000
1!
1%
#684000000000
0!
0%
#684005000000
1!
1%
#684010000000
0!
0%
#684015000000
1!
1%
#684020000000
0!
0%
#684025000000
1!
1%
#684030000000
0!
0%
#684035000000
1!
1%
#684040000000
0!
0%
#684045000000
1!
1%
#684050000000
0!
0%
#684055000000
1!
1%
#684060000000
0!
0%
#684065000000
1!
1%
#684070000000
0!
0%
#684075000000
1!
1%
#684080000000
0!
0%
#684085000000
1!
1%
#684090000000
0!
0%
#684095000000
1!
1%
#684100000000
0!
0%
#684105000000
1!
1%
#684110000000
0!
0%
#684115000000
1!
1%
#684120000000
0!
0%
#684125000000
1!
1%
#684130000000
0!
0%
#684135000000
1!
1%
#684140000000
0!
0%
#684145000000
1!
1%
#684150000000
0!
0%
#684155000000
1!
1%
#684160000000
0!
0%
#684165000000
1!
1%
#684170000000
0!
0%
#684175000000
1!
1%
#684180000000
0!
0%
#684185000000
1!
1%
#684190000000
0!
0%
#684195000000
1!
1%
#684200000000
0!
0%
#684205000000
1!
1%
#684210000000
0!
0%
#684215000000
1!
1%
#684220000000
0!
0%
#684225000000
1!
1%
#684230000000
0!
0%
#684235000000
1!
1%
#684240000000
0!
0%
#684245000000
1!
1%
#684250000000
0!
0%
#684255000000
1!
1%
#684260000000
0!
0%
#684265000000
1!
1%
#684270000000
0!
0%
#684275000000
1!
1%
#684280000000
0!
0%
#684285000000
1!
1%
#684290000000
0!
0%
#684295000000
1!
1%
#684300000000
0!
0%
#684305000000
1!
1%
#684310000000
0!
0%
#684315000000
1!
1%
#684320000000
0!
0%
#684325000000
1!
1%
#684330000000
0!
0%
#684335000000
1!
1%
#684340000000
0!
0%
#684345000000
1!
1%
#684350000000
0!
0%
#684355000000
1!
1%
#684360000000
0!
0%
#684365000000
1!
1%
#684370000000
0!
0%
#684375000000
1!
1%
#684380000000
0!
0%
#684385000000
1!
1%
#684390000000
0!
0%
#684395000000
1!
1%
#684400000000
0!
0%
#684405000000
1!
1%
#684410000000
0!
0%
#684415000000
1!
1%
#684420000000
0!
0%
#684425000000
1!
1%
#684430000000
0!
0%
#684435000000
1!
1%
#684440000000
0!
0%
#684445000000
1!
1%
#684450000000
0!
0%
#684455000000
1!
1%
#684460000000
0!
0%
#684465000000
1!
1%
#684470000000
0!
0%
#684475000000
1!
1%
#684480000000
0!
0%
#684485000000
1!
1%
#684490000000
0!
0%
#684495000000
1!
1%
#684500000000
0!
0%
#684505000000
1!
1%
#684510000000
0!
0%
#684515000000
1!
1%
#684520000000
0!
0%
#684525000000
1!
1%
#684530000000
0!
0%
#684535000000
1!
1%
#684540000000
0!
0%
#684545000000
1!
1%
#684550000000
0!
0%
#684555000000
1!
1%
#684560000000
0!
0%
#684565000000
1!
1%
#684570000000
0!
0%
#684575000000
1!
1%
#684580000000
0!
0%
#684585000000
1!
1%
#684590000000
0!
0%
#684595000000
1!
1%
#684600000000
0!
0%
#684605000000
1!
1%
#684610000000
0!
0%
#684615000000
1!
1%
#684620000000
0!
0%
#684625000000
1!
1%
#684630000000
0!
0%
#684635000000
1!
1%
#684640000000
0!
0%
#684645000000
1!
1%
#684650000000
0!
0%
#684655000000
1!
1%
#684660000000
0!
0%
#684665000000
1!
1%
#684670000000
0!
0%
#684675000000
1!
1%
#684680000000
0!
0%
#684685000000
1!
1%
#684690000000
0!
0%
#684695000000
1!
1%
#684700000000
0!
0%
#684705000000
1!
1%
#684710000000
0!
0%
#684715000000
1!
1%
#684720000000
0!
0%
#684725000000
1!
1%
#684730000000
0!
0%
#684735000000
1!
1%
#684740000000
0!
0%
#684745000000
1!
1%
#684750000000
0!
0%
#684755000000
1!
1%
#684760000000
0!
0%
#684765000000
1!
1%
#684770000000
0!
0%
#684775000000
1!
1%
#684780000000
0!
0%
#684785000000
1!
1%
#684790000000
0!
0%
#684795000000
1!
1%
#684800000000
0!
0%
#684805000000
1!
1%
#684810000000
0!
0%
#684815000000
1!
1%
#684820000000
0!
0%
#684825000000
1!
1%
#684830000000
0!
0%
#684835000000
1!
1%
#684840000000
0!
0%
#684845000000
1!
1%
#684850000000
0!
0%
#684855000000
1!
1%
#684860000000
0!
0%
#684865000000
1!
1%
#684870000000
0!
0%
#684875000000
1!
1%
#684880000000
0!
0%
#684885000000
1!
1%
#684890000000
0!
0%
#684895000000
1!
1%
#684900000000
0!
0%
#684905000000
1!
1%
#684910000000
0!
0%
#684915000000
1!
1%
#684920000000
0!
0%
#684925000000
1!
1%
#684930000000
0!
0%
#684935000000
1!
1%
#684940000000
0!
0%
#684945000000
1!
1%
#684950000000
0!
0%
#684955000000
1!
1%
#684960000000
0!
0%
#684965000000
1!
1%
#684970000000
0!
0%
#684975000000
1!
1%
#684980000000
0!
0%
#684985000000
1!
1%
#684990000000
0!
0%
#684995000000
1!
1%
#685000000000
0!
0%
#685005000000
1!
1%
#685010000000
0!
0%
#685015000000
1!
1%
#685020000000
0!
0%
#685025000000
1!
1%
#685030000000
0!
0%
#685035000000
1!
1%
#685040000000
0!
0%
#685045000000
1!
1%
#685050000000
0!
0%
#685055000000
1!
1%
#685060000000
0!
0%
#685065000000
1!
1%
#685070000000
0!
0%
#685075000000
1!
1%
#685080000000
0!
0%
#685085000000
1!
1%
#685090000000
0!
0%
#685095000000
1!
1%
#685100000000
0!
0%
#685105000000
1!
1%
#685110000000
0!
0%
#685115000000
1!
1%
#685120000000
0!
0%
#685125000000
1!
1%
#685130000000
0!
0%
#685135000000
1!
1%
#685140000000
0!
0%
#685145000000
1!
1%
#685150000000
0!
0%
#685155000000
1!
1%
#685160000000
0!
0%
#685165000000
1!
1%
#685170000000
0!
0%
#685175000000
1!
1%
#685180000000
0!
0%
#685185000000
1!
1%
#685190000000
0!
0%
#685195000000
1!
1%
#685200000000
0!
0%
#685205000000
1!
1%
#685210000000
0!
0%
#685215000000
1!
1%
#685220000000
0!
0%
#685225000000
1!
1%
#685230000000
0!
0%
#685235000000
1!
1%
#685240000000
0!
0%
#685245000000
1!
1%
#685250000000
0!
0%
#685255000000
1!
1%
#685260000000
0!
0%
#685265000000
1!
1%
#685270000000
0!
0%
#685275000000
1!
1%
#685280000000
0!
0%
#685285000000
1!
1%
#685290000000
0!
0%
#685295000000
1!
1%
#685300000000
0!
0%
#685305000000
1!
1%
#685310000000
0!
0%
#685315000000
1!
1%
#685320000000
0!
0%
#685325000000
1!
1%
#685330000000
0!
0%
#685335000000
1!
1%
#685340000000
0!
0%
#685345000000
1!
1%
#685350000000
0!
0%
#685355000000
1!
1%
#685360000000
0!
0%
#685365000000
1!
1%
#685370000000
0!
0%
#685375000000
1!
1%
#685380000000
0!
0%
#685385000000
1!
1%
#685390000000
0!
0%
#685395000000
1!
1%
#685400000000
0!
0%
#685405000000
1!
1%
#685410000000
0!
0%
#685415000000
1!
1%
#685420000000
0!
0%
#685425000000
1!
1%
#685430000000
0!
0%
#685435000000
1!
1%
#685440000000
0!
0%
#685445000000
1!
1%
#685450000000
0!
0%
#685455000000
1!
1%
#685460000000
0!
0%
#685465000000
1!
1%
#685470000000
0!
0%
#685475000000
1!
1%
#685480000000
0!
0%
#685485000000
1!
1%
#685490000000
0!
0%
#685495000000
1!
1%
#685500000000
0!
0%
#685505000000
1!
1%
#685510000000
0!
0%
#685515000000
1!
1%
#685520000000
0!
0%
#685525000000
1!
1%
#685530000000
0!
0%
#685535000000
1!
1%
#685540000000
0!
0%
#685545000000
1!
1%
#685550000000
0!
0%
#685555000000
1!
1%
#685560000000
0!
0%
#685565000000
1!
1%
#685570000000
0!
0%
#685575000000
1!
1%
#685580000000
0!
0%
#685585000000
1!
1%
#685590000000
0!
0%
#685595000000
1!
1%
#685600000000
0!
0%
#685605000000
1!
1%
#685610000000
0!
0%
#685615000000
1!
1%
#685620000000
0!
0%
#685625000000
1!
1%
#685630000000
0!
0%
#685635000000
1!
1%
#685640000000
0!
0%
#685645000000
1!
1%
#685650000000
0!
0%
#685655000000
1!
1%
#685660000000
0!
0%
#685665000000
1!
1%
#685670000000
0!
0%
#685675000000
1!
1%
#685680000000
0!
0%
#685685000000
1!
1%
#685690000000
0!
0%
#685695000000
1!
1%
#685700000000
0!
0%
#685705000000
1!
1%
#685710000000
0!
0%
#685715000000
1!
1%
#685720000000
0!
0%
#685725000000
1!
1%
#685730000000
0!
0%
#685735000000
1!
1%
#685740000000
0!
0%
#685745000000
1!
1%
#685750000000
0!
0%
#685755000000
1!
1%
#685760000000
0!
0%
#685765000000
1!
1%
#685770000000
0!
0%
#685775000000
1!
1%
#685780000000
0!
0%
#685785000000
1!
1%
#685790000000
0!
0%
#685795000000
1!
1%
#685800000000
0!
0%
#685805000000
1!
1%
#685810000000
0!
0%
#685815000000
1!
1%
#685820000000
0!
0%
#685825000000
1!
1%
#685830000000
0!
0%
#685835000000
1!
1%
#685840000000
0!
0%
#685845000000
1!
1%
#685850000000
0!
0%
#685855000000
1!
1%
#685860000000
0!
0%
#685865000000
1!
1%
#685870000000
0!
0%
#685875000000
1!
1%
#685880000000
0!
0%
#685885000000
1!
1%
#685890000000
0!
0%
#685895000000
1!
1%
#685900000000
0!
0%
#685905000000
1!
1%
#685910000000
0!
0%
#685915000000
1!
1%
#685920000000
0!
0%
#685925000000
1!
1%
#685930000000
0!
0%
#685935000000
1!
1%
#685940000000
0!
0%
#685945000000
1!
1%
#685950000000
0!
0%
#685955000000
1!
1%
#685960000000
0!
0%
#685965000000
1!
1%
#685970000000
0!
0%
#685975000000
1!
1%
#685980000000
0!
0%
#685985000000
1!
1%
#685990000000
0!
0%
#685995000000
1!
1%
#686000000000
0!
0%
#686005000000
1!
1%
#686010000000
0!
0%
#686015000000
1!
1%
#686020000000
0!
0%
#686025000000
1!
1%
#686030000000
0!
0%
#686035000000
1!
1%
#686040000000
0!
0%
#686045000000
1!
1%
#686050000000
0!
0%
#686055000000
1!
1%
#686060000000
0!
0%
#686065000000
1!
1%
#686070000000
0!
0%
#686075000000
1!
1%
#686080000000
0!
0%
#686085000000
1!
1%
#686090000000
0!
0%
#686095000000
1!
1%
#686100000000
0!
0%
#686105000000
1!
1%
#686110000000
0!
0%
#686115000000
1!
1%
#686120000000
0!
0%
#686125000000
1!
1%
#686130000000
0!
0%
#686135000000
1!
1%
#686140000000
0!
0%
#686145000000
1!
1%
#686150000000
0!
0%
#686155000000
1!
1%
#686160000000
0!
0%
#686165000000
1!
1%
#686170000000
0!
0%
#686175000000
1!
1%
#686180000000
0!
0%
#686185000000
1!
1%
#686190000000
0!
0%
#686195000000
1!
1%
#686200000000
0!
0%
#686205000000
1!
1%
#686210000000
0!
0%
#686215000000
1!
1%
#686220000000
0!
0%
#686225000000
1!
1%
#686230000000
0!
0%
#686235000000
1!
1%
#686240000000
0!
0%
#686245000000
1!
1%
#686250000000
0!
0%
#686255000000
1!
1%
#686260000000
0!
0%
#686265000000
1!
1%
#686270000000
0!
0%
#686275000000
1!
1%
#686280000000
0!
0%
#686285000000
1!
1%
#686290000000
0!
0%
#686295000000
1!
1%
#686300000000
0!
0%
#686305000000
1!
1%
#686310000000
0!
0%
#686315000000
1!
1%
#686320000000
0!
0%
#686325000000
1!
1%
#686330000000
0!
0%
#686335000000
1!
1%
#686340000000
0!
0%
#686345000000
1!
1%
#686350000000
0!
0%
#686355000000
1!
1%
#686360000000
0!
0%
#686365000000
1!
1%
#686370000000
0!
0%
#686375000000
1!
1%
#686380000000
0!
0%
#686385000000
1!
1%
#686390000000
0!
0%
#686395000000
1!
1%
#686400000000
0!
0%
#686405000000
1!
1%
#686410000000
0!
0%
#686415000000
1!
1%
#686420000000
0!
0%
#686425000000
1!
1%
#686430000000
0!
0%
#686435000000
1!
1%
#686440000000
0!
0%
#686445000000
1!
1%
#686450000000
0!
0%
#686455000000
1!
1%
#686460000000
0!
0%
#686465000000
1!
1%
#686470000000
0!
0%
#686475000000
1!
1%
#686480000000
0!
0%
#686485000000
1!
1%
#686490000000
0!
0%
#686495000000
1!
1%
#686500000000
0!
0%
#686505000000
1!
1%
#686510000000
0!
0%
#686515000000
1!
1%
#686520000000
0!
0%
#686525000000
1!
1%
#686530000000
0!
0%
#686535000000
1!
1%
#686540000000
0!
0%
#686545000000
1!
1%
#686550000000
0!
0%
#686555000000
1!
1%
#686560000000
0!
0%
#686565000000
1!
1%
#686570000000
0!
0%
#686575000000
1!
1%
#686580000000
0!
0%
#686585000000
1!
1%
#686590000000
0!
0%
#686595000000
1!
1%
#686600000000
0!
0%
#686605000000
1!
1%
#686610000000
0!
0%
#686615000000
1!
1%
#686620000000
0!
0%
#686625000000
1!
1%
#686630000000
0!
0%
#686635000000
1!
1%
#686640000000
0!
0%
#686645000000
1!
1%
#686650000000
0!
0%
#686655000000
1!
1%
#686660000000
0!
0%
#686665000000
1!
1%
#686670000000
0!
0%
#686675000000
1!
1%
#686680000000
0!
0%
#686685000000
1!
1%
#686690000000
0!
0%
#686695000000
1!
1%
#686700000000
0!
0%
#686705000000
1!
1%
#686710000000
0!
0%
#686715000000
1!
1%
#686720000000
0!
0%
#686725000000
1!
1%
#686730000000
0!
0%
#686735000000
1!
1%
#686740000000
0!
0%
#686745000000
1!
1%
#686750000000
0!
0%
#686755000000
1!
1%
#686760000000
0!
0%
#686765000000
1!
1%
#686770000000
0!
0%
#686775000000
1!
1%
#686780000000
0!
0%
#686785000000
1!
1%
#686790000000
0!
0%
#686795000000
1!
1%
#686800000000
0!
0%
#686805000000
1!
1%
#686810000000
0!
0%
#686815000000
1!
1%
#686820000000
0!
0%
#686825000000
1!
1%
#686830000000
0!
0%
#686835000000
1!
1%
#686840000000
0!
0%
#686845000000
1!
1%
#686850000000
0!
0%
#686855000000
1!
1%
#686860000000
0!
0%
#686865000000
1!
1%
#686870000000
0!
0%
#686875000000
1!
1%
#686880000000
0!
0%
#686885000000
1!
1%
#686890000000
0!
0%
#686895000000
1!
1%
#686900000000
0!
0%
#686905000000
1!
1%
#686910000000
0!
0%
#686915000000
1!
1%
#686920000000
0!
0%
#686925000000
1!
1%
#686930000000
0!
0%
#686935000000
1!
1%
#686940000000
0!
0%
#686945000000
1!
1%
#686950000000
0!
0%
#686955000000
1!
1%
#686960000000
0!
0%
#686965000000
1!
1%
#686970000000
0!
0%
#686975000000
1!
1%
#686980000000
0!
0%
#686985000000
1!
1%
#686990000000
0!
0%
#686995000000
1!
1%
#687000000000
0!
0%
#687005000000
1!
1%
#687010000000
0!
0%
#687015000000
1!
1%
#687020000000
0!
0%
#687025000000
1!
1%
#687030000000
0!
0%
#687035000000
1!
1%
#687040000000
0!
0%
#687045000000
1!
1%
#687050000000
0!
0%
#687055000000
1!
1%
#687060000000
0!
0%
#687065000000
1!
1%
#687070000000
0!
0%
#687075000000
1!
1%
#687080000000
0!
0%
#687085000000
1!
1%
#687090000000
0!
0%
#687095000000
1!
1%
#687100000000
0!
0%
#687105000000
1!
1%
#687110000000
0!
0%
#687115000000
1!
1%
#687120000000
0!
0%
#687125000000
1!
1%
#687130000000
0!
0%
#687135000000
1!
1%
#687140000000
0!
0%
#687145000000
1!
1%
#687150000000
0!
0%
#687155000000
1!
1%
#687160000000
0!
0%
#687165000000
1!
1%
#687170000000
0!
0%
#687175000000
1!
1%
#687180000000
0!
0%
#687185000000
1!
1%
#687190000000
0!
0%
#687195000000
1!
1%
#687200000000
0!
0%
#687205000000
1!
1%
#687210000000
0!
0%
#687215000000
1!
1%
#687220000000
0!
0%
#687225000000
1!
1%
#687230000000
0!
0%
#687235000000
1!
1%
#687240000000
0!
0%
#687245000000
1!
1%
#687250000000
0!
0%
#687255000000
1!
1%
#687260000000
0!
0%
#687265000000
1!
1%
#687270000000
0!
0%
#687275000000
1!
1%
#687280000000
0!
0%
#687285000000
1!
1%
#687290000000
0!
0%
#687295000000
1!
1%
#687300000000
0!
0%
#687305000000
1!
1%
#687310000000
0!
0%
#687315000000
1!
1%
#687320000000
0!
0%
#687325000000
1!
1%
#687330000000
0!
0%
#687335000000
1!
1%
#687340000000
0!
0%
#687345000000
1!
1%
#687350000000
0!
0%
#687355000000
1!
1%
#687360000000
0!
0%
#687365000000
1!
1%
#687370000000
0!
0%
#687375000000
1!
1%
#687380000000
0!
0%
#687385000000
1!
1%
#687390000000
0!
0%
#687395000000
1!
1%
#687400000000
0!
0%
#687405000000
1!
1%
#687410000000
0!
0%
#687415000000
1!
1%
#687420000000
0!
0%
#687425000000
1!
1%
#687430000000
0!
0%
#687435000000
1!
1%
#687440000000
0!
0%
#687445000000
1!
1%
#687450000000
0!
0%
#687455000000
1!
1%
#687460000000
0!
0%
#687465000000
1!
1%
#687470000000
0!
0%
#687475000000
1!
1%
#687480000000
0!
0%
#687485000000
1!
1%
#687490000000
0!
0%
#687495000000
1!
1%
#687500000000
0!
0%
#687505000000
1!
1%
#687510000000
0!
0%
#687515000000
1!
1%
#687520000000
0!
0%
#687525000000
1!
1%
#687530000000
0!
0%
#687535000000
1!
1%
#687540000000
0!
0%
#687545000000
1!
1%
#687550000000
0!
0%
#687555000000
1!
1%
#687560000000
0!
0%
#687565000000
1!
1%
#687570000000
0!
0%
#687575000000
1!
1%
#687580000000
0!
0%
#687585000000
1!
1%
#687590000000
0!
0%
#687595000000
1!
1%
#687600000000
0!
0%
#687605000000
1!
1%
#687610000000
0!
0%
#687615000000
1!
1%
#687620000000
0!
0%
#687625000000
1!
1%
#687630000000
0!
0%
#687635000000
1!
1%
#687640000000
0!
0%
#687645000000
1!
1%
#687650000000
0!
0%
#687655000000
1!
1%
#687660000000
0!
0%
#687665000000
1!
1%
#687670000000
0!
0%
#687675000000
1!
1%
#687680000000
0!
0%
#687685000000
1!
1%
#687690000000
0!
0%
#687695000000
1!
1%
#687700000000
0!
0%
#687705000000
1!
1%
#687710000000
0!
0%
#687715000000
1!
1%
#687720000000
0!
0%
#687725000000
1!
1%
#687730000000
0!
0%
#687735000000
1!
1%
#687740000000
0!
0%
#687745000000
1!
1%
#687750000000
0!
0%
#687755000000
1!
1%
#687760000000
0!
0%
#687765000000
1!
1%
#687770000000
0!
0%
#687775000000
1!
1%
#687780000000
0!
0%
#687785000000
1!
1%
#687790000000
0!
0%
#687795000000
1!
1%
#687800000000
0!
0%
#687805000000
1!
1%
#687810000000
0!
0%
#687815000000
1!
1%
#687820000000
0!
0%
#687825000000
1!
1%
#687830000000
0!
0%
#687835000000
1!
1%
#687840000000
0!
0%
#687845000000
1!
1%
#687850000000
0!
0%
#687855000000
1!
1%
#687860000000
0!
0%
#687865000000
1!
1%
#687870000000
0!
0%
#687875000000
1!
1%
#687880000000
0!
0%
#687885000000
1!
1%
#687890000000
0!
0%
#687895000000
1!
1%
#687900000000
0!
0%
#687905000000
1!
1%
#687910000000
0!
0%
#687915000000
1!
1%
#687920000000
0!
0%
#687925000000
1!
1%
#687930000000
0!
0%
#687935000000
1!
1%
#687940000000
0!
0%
#687945000000
1!
1%
#687950000000
0!
0%
#687955000000
1!
1%
#687960000000
0!
0%
#687965000000
1!
1%
#687970000000
0!
0%
#687975000000
1!
1%
#687980000000
0!
0%
#687985000000
1!
1%
#687990000000
0!
0%
#687995000000
1!
1%
#688000000000
0!
0%
#688005000000
1!
1%
#688010000000
0!
0%
#688015000000
1!
1%
#688020000000
0!
0%
#688025000000
1!
1%
#688030000000
0!
0%
#688035000000
1!
1%
#688040000000
0!
0%
#688045000000
1!
1%
#688050000000
0!
0%
#688055000000
1!
1%
#688060000000
0!
0%
#688065000000
1!
1%
#688070000000
0!
0%
#688075000000
1!
1%
#688080000000
0!
0%
#688085000000
1!
1%
#688090000000
0!
0%
#688095000000
1!
1%
#688100000000
0!
0%
#688105000000
1!
1%
#688110000000
0!
0%
#688115000000
1!
1%
#688120000000
0!
0%
#688125000000
1!
1%
#688130000000
0!
0%
#688135000000
1!
1%
#688140000000
0!
0%
#688145000000
1!
1%
#688150000000
0!
0%
#688155000000
1!
1%
#688160000000
0!
0%
#688165000000
1!
1%
#688170000000
0!
0%
#688175000000
1!
1%
#688180000000
0!
0%
#688185000000
1!
1%
#688190000000
0!
0%
#688195000000
1!
1%
#688200000000
0!
0%
#688205000000
1!
1%
#688210000000
0!
0%
#688215000000
1!
1%
#688220000000
0!
0%
#688225000000
1!
1%
#688230000000
0!
0%
#688235000000
1!
1%
#688240000000
0!
0%
#688245000000
1!
1%
#688250000000
0!
0%
#688255000000
1!
1%
#688260000000
0!
0%
#688265000000
1!
1%
#688270000000
0!
0%
#688275000000
1!
1%
#688280000000
0!
0%
#688285000000
1!
1%
#688290000000
0!
0%
#688295000000
1!
1%
#688300000000
0!
0%
#688305000000
1!
1%
#688310000000
0!
0%
#688315000000
1!
1%
#688320000000
0!
0%
#688325000000
1!
1%
#688330000000
0!
0%
#688335000000
1!
1%
#688340000000
0!
0%
#688345000000
1!
1%
#688350000000
0!
0%
#688355000000
1!
1%
#688360000000
0!
0%
#688365000000
1!
1%
#688370000000
0!
0%
#688375000000
1!
1%
#688380000000
0!
0%
#688385000000
1!
1%
#688390000000
0!
0%
#688395000000
1!
1%
#688400000000
0!
0%
#688405000000
1!
1%
#688410000000
0!
0%
#688415000000
1!
1%
#688420000000
0!
0%
#688425000000
1!
1%
#688430000000
0!
0%
#688435000000
1!
1%
#688440000000
0!
0%
#688445000000
1!
1%
#688450000000
0!
0%
#688455000000
1!
1%
#688460000000
0!
0%
#688465000000
1!
1%
#688470000000
0!
0%
#688475000000
1!
1%
#688480000000
0!
0%
#688485000000
1!
1%
#688490000000
0!
0%
#688495000000
1!
1%
#688500000000
0!
0%
#688505000000
1!
1%
#688510000000
0!
0%
#688515000000
1!
1%
#688520000000
0!
0%
#688525000000
1!
1%
#688530000000
0!
0%
#688535000000
1!
1%
#688540000000
0!
0%
#688545000000
1!
1%
#688550000000
0!
0%
#688555000000
1!
1%
#688560000000
0!
0%
#688565000000
1!
1%
#688570000000
0!
0%
#688575000000
1!
1%
#688580000000
0!
0%
#688585000000
1!
1%
#688590000000
0!
0%
#688595000000
1!
1%
#688600000000
0!
0%
#688605000000
1!
1%
#688610000000
0!
0%
#688615000000
1!
1%
#688620000000
0!
0%
#688625000000
1!
1%
#688630000000
0!
0%
#688635000000
1!
1%
#688640000000
0!
0%
#688645000000
1!
1%
#688650000000
0!
0%
#688655000000
1!
1%
#688660000000
0!
0%
#688665000000
1!
1%
#688670000000
0!
0%
#688675000000
1!
1%
#688680000000
0!
0%
#688685000000
1!
1%
#688690000000
0!
0%
#688695000000
1!
1%
#688700000000
0!
0%
#688705000000
1!
1%
#688710000000
0!
0%
#688715000000
1!
1%
#688720000000
0!
0%
#688725000000
1!
1%
#688730000000
0!
0%
#688735000000
1!
1%
#688740000000
0!
0%
#688745000000
1!
1%
#688750000000
0!
0%
#688755000000
1!
1%
#688760000000
0!
0%
#688765000000
1!
1%
#688770000000
0!
0%
#688775000000
1!
1%
#688780000000
0!
0%
#688785000000
1!
1%
#688790000000
0!
0%
#688795000000
1!
1%
#688800000000
0!
0%
#688805000000
1!
1%
#688810000000
0!
0%
#688815000000
1!
1%
#688820000000
0!
0%
#688825000000
1!
1%
#688830000000
0!
0%
#688835000000
1!
1%
#688840000000
0!
0%
#688845000000
1!
1%
#688850000000
0!
0%
#688855000000
1!
1%
#688860000000
0!
0%
#688865000000
1!
1%
#688870000000
0!
0%
#688875000000
1!
1%
#688880000000
0!
0%
#688885000000
1!
1%
#688890000000
0!
0%
#688895000000
1!
1%
#688900000000
0!
0%
#688905000000
1!
1%
#688910000000
0!
0%
#688915000000
1!
1%
#688920000000
0!
0%
#688925000000
1!
1%
#688930000000
0!
0%
#688935000000
1!
1%
#688940000000
0!
0%
#688945000000
1!
1%
#688950000000
0!
0%
#688955000000
1!
1%
#688960000000
0!
0%
#688965000000
1!
1%
#688970000000
0!
0%
#688975000000
1!
1%
#688980000000
0!
0%
#688985000000
1!
1%
#688990000000
0!
0%
#688995000000
1!
1%
#689000000000
0!
0%
#689005000000
1!
1%
#689010000000
0!
0%
#689015000000
1!
1%
#689020000000
0!
0%
#689025000000
1!
1%
#689030000000
0!
0%
#689035000000
1!
1%
#689040000000
0!
0%
#689045000000
1!
1%
#689050000000
0!
0%
#689055000000
1!
1%
#689060000000
0!
0%
#689065000000
1!
1%
#689070000000
0!
0%
#689075000000
1!
1%
#689080000000
0!
0%
#689085000000
1!
1%
#689090000000
0!
0%
#689095000000
1!
1%
#689100000000
0!
0%
#689105000000
1!
1%
#689110000000
0!
0%
#689115000000
1!
1%
#689120000000
0!
0%
#689125000000
1!
1%
#689130000000
0!
0%
#689135000000
1!
1%
#689140000000
0!
0%
#689145000000
1!
1%
#689150000000
0!
0%
#689155000000
1!
1%
#689160000000
0!
0%
#689165000000
1!
1%
#689170000000
0!
0%
#689175000000
1!
1%
#689180000000
0!
0%
#689185000000
1!
1%
#689190000000
0!
0%
#689195000000
1!
1%
#689200000000
0!
0%
#689205000000
1!
1%
#689210000000
0!
0%
#689215000000
1!
1%
#689220000000
0!
0%
#689225000000
1!
1%
#689230000000
0!
0%
#689235000000
1!
1%
#689240000000
0!
0%
#689245000000
1!
1%
#689250000000
0!
0%
#689255000000
1!
1%
#689260000000
0!
0%
#689265000000
1!
1%
#689270000000
0!
0%
#689275000000
1!
1%
#689280000000
0!
0%
#689285000000
1!
1%
#689290000000
0!
0%
#689295000000
1!
1%
#689300000000
0!
0%
#689305000000
1!
1%
#689310000000
0!
0%
#689315000000
1!
1%
#689320000000
0!
0%
#689325000000
1!
1%
#689330000000
0!
0%
#689335000000
1!
1%
#689340000000
0!
0%
#689345000000
1!
1%
#689350000000
0!
0%
#689355000000
1!
1%
#689360000000
0!
0%
#689365000000
1!
1%
#689370000000
0!
0%
#689375000000
1!
1%
#689380000000
0!
0%
#689385000000
1!
1%
#689390000000
0!
0%
#689395000000
1!
1%
#689400000000
0!
0%
#689405000000
1!
1%
#689410000000
0!
0%
#689415000000
1!
1%
#689420000000
0!
0%
#689425000000
1!
1%
#689430000000
0!
0%
#689435000000
1!
1%
#689440000000
0!
0%
#689445000000
1!
1%
#689450000000
0!
0%
#689455000000
1!
1%
#689460000000
0!
0%
#689465000000
1!
1%
#689470000000
0!
0%
#689475000000
1!
1%
#689480000000
0!
0%
#689485000000
1!
1%
#689490000000
0!
0%
#689495000000
1!
1%
#689500000000
0!
0%
#689505000000
1!
1%
#689510000000
0!
0%
#689515000000
1!
1%
#689520000000
0!
0%
#689525000000
1!
1%
#689530000000
0!
0%
#689535000000
1!
1%
#689540000000
0!
0%
#689545000000
1!
1%
#689550000000
0!
0%
#689555000000
1!
1%
#689560000000
0!
0%
#689565000000
1!
1%
#689570000000
0!
0%
#689575000000
1!
1%
#689580000000
0!
0%
#689585000000
1!
1%
#689590000000
0!
0%
#689595000000
1!
1%
#689600000000
0!
0%
#689605000000
1!
1%
#689610000000
0!
0%
#689615000000
1!
1%
#689620000000
0!
0%
#689625000000
1!
1%
#689630000000
0!
0%
#689635000000
1!
1%
#689640000000
0!
0%
#689645000000
1!
1%
#689650000000
0!
0%
#689655000000
1!
1%
#689660000000
0!
0%
#689665000000
1!
1%
#689670000000
0!
0%
#689675000000
1!
1%
#689680000000
0!
0%
#689685000000
1!
1%
#689690000000
0!
0%
#689695000000
1!
1%
#689700000000
0!
0%
#689705000000
1!
1%
#689710000000
0!
0%
#689715000000
1!
1%
#689720000000
0!
0%
#689725000000
1!
1%
#689730000000
0!
0%
#689735000000
1!
1%
#689740000000
0!
0%
#689745000000
1!
1%
#689750000000
0!
0%
#689755000000
1!
1%
#689760000000
0!
0%
#689765000000
1!
1%
#689770000000
0!
0%
#689775000000
1!
1%
#689780000000
0!
0%
#689785000000
1!
1%
#689790000000
0!
0%
#689795000000
1!
1%
#689800000000
0!
0%
#689805000000
1!
1%
#689810000000
0!
0%
#689815000000
1!
1%
#689820000000
0!
0%
#689825000000
1!
1%
#689830000000
0!
0%
#689835000000
1!
1%
#689840000000
0!
0%
#689845000000
1!
1%
#689850000000
0!
0%
#689855000000
1!
1%
#689860000000
0!
0%
#689865000000
1!
1%
#689870000000
0!
0%
#689875000000
1!
1%
#689880000000
0!
0%
#689885000000
1!
1%
#689890000000
0!
0%
#689895000000
1!
1%
#689900000000
0!
0%
#689905000000
1!
1%
#689910000000
0!
0%
#689915000000
1!
1%
#689920000000
0!
0%
#689925000000
1!
1%
#689930000000
0!
0%
#689935000000
1!
1%
#689940000000
0!
0%
#689945000000
1!
1%
#689950000000
0!
0%
#689955000000
1!
1%
#689960000000
0!
0%
#689965000000
1!
1%
#689970000000
0!
0%
#689975000000
1!
1%
#689980000000
0!
0%
#689985000000
1!
1%
#689990000000
0!
0%
#689995000000
1!
1%
#690000000000
0!
0%
#690005000000
1!
1%
#690010000000
0!
0%
#690015000000
1!
1%
#690020000000
0!
0%
#690025000000
1!
1%
#690030000000
0!
0%
#690035000000
1!
1%
#690040000000
0!
0%
#690045000000
1!
1%
#690050000000
0!
0%
#690055000000
1!
1%
#690060000000
0!
0%
#690065000000
1!
1%
#690070000000
0!
0%
#690075000000
1!
1%
#690080000000
0!
0%
#690085000000
1!
1%
#690090000000
0!
0%
#690095000000
1!
1%
#690100000000
0!
0%
#690105000000
1!
1%
#690110000000
0!
0%
#690115000000
1!
1%
#690120000000
0!
0%
#690125000000
1!
1%
#690130000000
0!
0%
#690135000000
1!
1%
#690140000000
0!
0%
#690145000000
1!
1%
#690150000000
0!
0%
#690155000000
1!
1%
#690160000000
0!
0%
#690165000000
1!
1%
#690170000000
0!
0%
#690175000000
1!
1%
#690180000000
0!
0%
#690185000000
1!
1%
#690190000000
0!
0%
#690195000000
1!
1%
#690200000000
0!
0%
#690205000000
1!
1%
#690210000000
0!
0%
#690215000000
1!
1%
#690220000000
0!
0%
#690225000000
1!
1%
#690230000000
0!
0%
#690235000000
1!
1%
#690240000000
0!
0%
#690245000000
1!
1%
#690250000000
0!
0%
#690255000000
1!
1%
#690260000000
0!
0%
#690265000000
1!
1%
#690270000000
0!
0%
#690275000000
1!
1%
#690280000000
0!
0%
#690285000000
1!
1%
#690290000000
0!
0%
#690295000000
1!
1%
#690300000000
0!
0%
#690305000000
1!
1%
#690310000000
0!
0%
#690315000000
1!
1%
#690320000000
0!
0%
#690325000000
1!
1%
#690330000000
0!
0%
#690335000000
1!
1%
#690340000000
0!
0%
#690345000000
1!
1%
#690350000000
0!
0%
#690355000000
1!
1%
#690360000000
0!
0%
#690365000000
1!
1%
#690370000000
0!
0%
#690375000000
1!
1%
#690380000000
0!
0%
#690385000000
1!
1%
#690390000000
0!
0%
#690395000000
1!
1%
#690400000000
0!
0%
#690405000000
1!
1%
#690410000000
0!
0%
#690415000000
1!
1%
#690420000000
0!
0%
#690425000000
1!
1%
#690430000000
0!
0%
#690435000000
1!
1%
#690440000000
0!
0%
#690445000000
1!
1%
#690450000000
0!
0%
#690455000000
1!
1%
#690460000000
0!
0%
#690465000000
1!
1%
#690470000000
0!
0%
#690475000000
1!
1%
#690480000000
0!
0%
#690485000000
1!
1%
#690490000000
0!
0%
#690495000000
1!
1%
#690500000000
0!
0%
#690505000000
1!
1%
#690510000000
0!
0%
#690515000000
1!
1%
#690520000000
0!
0%
#690525000000
1!
1%
#690530000000
0!
0%
#690535000000
1!
1%
#690540000000
0!
0%
#690545000000
1!
1%
#690550000000
0!
0%
#690555000000
1!
1%
#690560000000
0!
0%
#690565000000
1!
1%
#690570000000
0!
0%
#690575000000
1!
1%
#690580000000
0!
0%
#690585000000
1!
1%
#690590000000
0!
0%
#690595000000
1!
1%
#690600000000
0!
0%
#690605000000
1!
1%
#690610000000
0!
0%
#690615000000
1!
1%
#690620000000
0!
0%
#690625000000
1!
1%
#690630000000
0!
0%
#690635000000
1!
1%
#690640000000
0!
0%
#690645000000
1!
1%
#690650000000
0!
0%
#690655000000
1!
1%
#690660000000
0!
0%
#690665000000
1!
1%
#690670000000
0!
0%
#690675000000
1!
1%
#690680000000
0!
0%
#690685000000
1!
1%
#690690000000
0!
0%
#690695000000
1!
1%
#690700000000
0!
0%
#690705000000
1!
1%
#690710000000
0!
0%
#690715000000
1!
1%
#690720000000
0!
0%
#690725000000
1!
1%
#690730000000
0!
0%
#690735000000
1!
1%
#690740000000
0!
0%
#690745000000
1!
1%
#690750000000
0!
0%
#690755000000
1!
1%
#690760000000
0!
0%
#690765000000
1!
1%
#690770000000
0!
0%
#690775000000
1!
1%
#690780000000
0!
0%
#690785000000
1!
1%
#690790000000
0!
0%
#690795000000
1!
1%
#690800000000
0!
0%
#690805000000
1!
1%
#690810000000
0!
0%
#690815000000
1!
1%
#690820000000
0!
0%
#690825000000
1!
1%
#690830000000
0!
0%
#690835000000
1!
1%
#690840000000
0!
0%
#690845000000
1!
1%
#690850000000
0!
0%
#690855000000
1!
1%
#690860000000
0!
0%
#690865000000
1!
1%
#690870000000
0!
0%
#690875000000
1!
1%
#690880000000
0!
0%
#690885000000
1!
1%
#690890000000
0!
0%
#690895000000
1!
1%
#690900000000
0!
0%
#690905000000
1!
1%
#690910000000
0!
0%
#690915000000
1!
1%
#690920000000
0!
0%
#690925000000
1!
1%
#690930000000
0!
0%
#690935000000
1!
1%
#690940000000
0!
0%
#690945000000
1!
1%
#690950000000
0!
0%
#690955000000
1!
1%
#690960000000
0!
0%
#690965000000
1!
1%
#690970000000
0!
0%
#690975000000
1!
1%
#690980000000
0!
0%
#690985000000
1!
1%
#690990000000
0!
0%
#690995000000
1!
1%
#691000000000
0!
0%
#691005000000
1!
1%
#691010000000
0!
0%
#691015000000
1!
1%
#691020000000
0!
0%
#691025000000
1!
1%
#691030000000
0!
0%
#691035000000
1!
1%
#691040000000
0!
0%
#691045000000
1!
1%
#691050000000
0!
0%
#691055000000
1!
1%
#691060000000
0!
0%
#691065000000
1!
1%
#691070000000
0!
0%
#691075000000
1!
1%
#691080000000
0!
0%
#691085000000
1!
1%
#691090000000
0!
0%
#691095000000
1!
1%
#691100000000
0!
0%
#691105000000
1!
1%
#691110000000
0!
0%
#691115000000
1!
1%
#691120000000
0!
0%
#691125000000
1!
1%
#691130000000
0!
0%
#691135000000
1!
1%
#691140000000
0!
0%
#691145000000
1!
1%
#691150000000
0!
0%
#691155000000
1!
1%
#691160000000
0!
0%
#691165000000
1!
1%
#691170000000
0!
0%
#691175000000
1!
1%
#691180000000
0!
0%
#691185000000
1!
1%
#691190000000
0!
0%
#691195000000
1!
1%
#691200000000
0!
0%
#691205000000
1!
1%
#691210000000
0!
0%
#691215000000
1!
1%
#691220000000
0!
0%
#691225000000
1!
1%
#691230000000
0!
0%
#691235000000
1!
1%
#691240000000
0!
0%
#691245000000
1!
1%
#691250000000
0!
0%
#691255000000
1!
1%
#691260000000
0!
0%
#691265000000
1!
1%
#691270000000
0!
0%
#691275000000
1!
1%
#691280000000
0!
0%
#691285000000
1!
1%
#691290000000
0!
0%
#691295000000
1!
1%
#691300000000
0!
0%
#691305000000
1!
1%
#691310000000
0!
0%
#691315000000
1!
1%
#691320000000
0!
0%
#691325000000
1!
1%
#691330000000
0!
0%
#691335000000
1!
1%
#691340000000
0!
0%
#691345000000
1!
1%
#691350000000
0!
0%
#691355000000
1!
1%
#691360000000
0!
0%
#691365000000
1!
1%
#691370000000
0!
0%
#691375000000
1!
1%
#691380000000
0!
0%
#691385000000
1!
1%
#691390000000
0!
0%
#691395000000
1!
1%
#691400000000
0!
0%
#691405000000
1!
1%
#691410000000
0!
0%
#691415000000
1!
1%
#691420000000
0!
0%
#691425000000
1!
1%
#691430000000
0!
0%
#691435000000
1!
1%
#691440000000
0!
0%
#691445000000
1!
1%
#691450000000
0!
0%
#691455000000
1!
1%
#691460000000
0!
0%
#691465000000
1!
1%
#691470000000
0!
0%
#691475000000
1!
1%
#691480000000
0!
0%
#691485000000
1!
1%
#691490000000
0!
0%
#691495000000
1!
1%
#691500000000
0!
0%
#691505000000
1!
1%
#691510000000
0!
0%
#691515000000
1!
1%
#691520000000
0!
0%
#691525000000
1!
1%
#691530000000
0!
0%
#691535000000
1!
1%
#691540000000
0!
0%
#691545000000
1!
1%
#691550000000
0!
0%
#691555000000
1!
1%
#691560000000
0!
0%
#691565000000
1!
1%
#691570000000
0!
0%
#691575000000
1!
1%
#691580000000
0!
0%
#691585000000
1!
1%
#691590000000
0!
0%
#691595000000
1!
1%
#691600000000
0!
0%
#691605000000
1!
1%
#691610000000
0!
0%
#691615000000
1!
1%
#691620000000
0!
0%
#691625000000
1!
1%
#691630000000
0!
0%
#691635000000
1!
1%
#691640000000
0!
0%
#691645000000
1!
1%
#691650000000
0!
0%
#691655000000
1!
1%
#691660000000
0!
0%
#691665000000
1!
1%
#691670000000
0!
0%
#691675000000
1!
1%
#691680000000
0!
0%
#691685000000
1!
1%
#691690000000
0!
0%
#691695000000
1!
1%
#691700000000
0!
0%
#691705000000
1!
1%
#691710000000
0!
0%
#691715000000
1!
1%
#691720000000
0!
0%
#691725000000
1!
1%
#691730000000
0!
0%
#691735000000
1!
1%
#691740000000
0!
0%
#691745000000
1!
1%
#691750000000
0!
0%
#691755000000
1!
1%
#691760000000
0!
0%
#691765000000
1!
1%
#691770000000
0!
0%
#691775000000
1!
1%
#691780000000
0!
0%
#691785000000
1!
1%
#691790000000
0!
0%
#691795000000
1!
1%
#691800000000
0!
0%
#691805000000
1!
1%
#691810000000
0!
0%
#691815000000
1!
1%
#691820000000
0!
0%
#691825000000
1!
1%
#691830000000
0!
0%
#691835000000
1!
1%
#691840000000
0!
0%
#691845000000
1!
1%
#691850000000
0!
0%
#691855000000
1!
1%
#691860000000
0!
0%
#691865000000
1!
1%
#691870000000
0!
0%
#691875000000
1!
1%
#691880000000
0!
0%
#691885000000
1!
1%
#691890000000
0!
0%
#691895000000
1!
1%
#691900000000
0!
0%
#691905000000
1!
1%
#691910000000
0!
0%
#691915000000
1!
1%
#691920000000
0!
0%
#691925000000
1!
1%
#691930000000
0!
0%
#691935000000
1!
1%
#691940000000
0!
0%
#691945000000
1!
1%
#691950000000
0!
0%
#691955000000
1!
1%
#691960000000
0!
0%
#691965000000
1!
1%
#691970000000
0!
0%
#691975000000
1!
1%
#691980000000
0!
0%
#691985000000
1!
1%
#691990000000
0!
0%
#691995000000
1!
1%
#692000000000
0!
0%
#692005000000
1!
1%
#692010000000
0!
0%
#692015000000
1!
1%
#692020000000
0!
0%
#692025000000
1!
1%
#692030000000
0!
0%
#692035000000
1!
1%
#692040000000
0!
0%
#692045000000
1!
1%
#692050000000
0!
0%
#692055000000
1!
1%
#692060000000
0!
0%
#692065000000
1!
1%
#692070000000
0!
0%
#692075000000
1!
1%
#692080000000
0!
0%
#692085000000
1!
1%
#692090000000
0!
0%
#692095000000
1!
1%
#692100000000
0!
0%
#692105000000
1!
1%
#692110000000
0!
0%
#692115000000
1!
1%
#692120000000
0!
0%
#692125000000
1!
1%
#692130000000
0!
0%
#692135000000
1!
1%
#692140000000
0!
0%
#692145000000
1!
1%
#692150000000
0!
0%
#692155000000
1!
1%
#692160000000
0!
0%
#692165000000
1!
1%
#692170000000
0!
0%
#692175000000
1!
1%
#692180000000
0!
0%
#692185000000
1!
1%
#692190000000
0!
0%
#692195000000
1!
1%
#692200000000
0!
0%
#692205000000
1!
1%
#692210000000
0!
0%
#692215000000
1!
1%
#692220000000
0!
0%
#692225000000
1!
1%
#692230000000
0!
0%
#692235000000
1!
1%
#692240000000
0!
0%
#692245000000
1!
1%
#692250000000
0!
0%
#692255000000
1!
1%
#692260000000
0!
0%
#692265000000
1!
1%
#692270000000
0!
0%
#692275000000
1!
1%
#692280000000
0!
0%
#692285000000
1!
1%
#692290000000
0!
0%
#692295000000
1!
1%
#692300000000
0!
0%
#692305000000
1!
1%
#692310000000
0!
0%
#692315000000
1!
1%
#692320000000
0!
0%
#692325000000
1!
1%
#692330000000
0!
0%
#692335000000
1!
1%
#692340000000
0!
0%
#692345000000
1!
1%
#692350000000
0!
0%
#692355000000
1!
1%
#692360000000
0!
0%
#692365000000
1!
1%
#692370000000
0!
0%
#692375000000
1!
1%
#692380000000
0!
0%
#692385000000
1!
1%
#692390000000
0!
0%
#692395000000
1!
1%
#692400000000
0!
0%
#692405000000
1!
1%
#692410000000
0!
0%
#692415000000
1!
1%
#692420000000
0!
0%
#692425000000
1!
1%
#692430000000
0!
0%
#692435000000
1!
1%
#692440000000
0!
0%
#692445000000
1!
1%
#692450000000
0!
0%
#692455000000
1!
1%
#692460000000
0!
0%
#692465000000
1!
1%
#692470000000
0!
0%
#692475000000
1!
1%
#692480000000
0!
0%
#692485000000
1!
1%
#692490000000
0!
0%
#692495000000
1!
1%
#692500000000
0!
0%
#692505000000
1!
1%
#692510000000
0!
0%
#692515000000
1!
1%
#692520000000
0!
0%
#692525000000
1!
1%
#692530000000
0!
0%
#692535000000
1!
1%
#692540000000
0!
0%
#692545000000
1!
1%
#692550000000
0!
0%
#692555000000
1!
1%
#692560000000
0!
0%
#692565000000
1!
1%
#692570000000
0!
0%
#692575000000
1!
1%
#692580000000
0!
0%
#692585000000
1!
1%
#692590000000
0!
0%
#692595000000
1!
1%
#692600000000
0!
0%
#692605000000
1!
1%
#692610000000
0!
0%
#692615000000
1!
1%
#692620000000
0!
0%
#692625000000
1!
1%
#692630000000
0!
0%
#692635000000
1!
1%
#692640000000
0!
0%
#692645000000
1!
1%
#692650000000
0!
0%
#692655000000
1!
1%
#692660000000
0!
0%
#692665000000
1!
1%
#692670000000
0!
0%
#692675000000
1!
1%
#692680000000
0!
0%
#692685000000
1!
1%
#692690000000
0!
0%
#692695000000
1!
1%
#692700000000
0!
0%
#692705000000
1!
1%
#692710000000
0!
0%
#692715000000
1!
1%
#692720000000
0!
0%
#692725000000
1!
1%
#692730000000
0!
0%
#692735000000
1!
1%
#692740000000
0!
0%
#692745000000
1!
1%
#692750000000
0!
0%
#692755000000
1!
1%
#692760000000
0!
0%
#692765000000
1!
1%
#692770000000
0!
0%
#692775000000
1!
1%
#692780000000
0!
0%
#692785000000
1!
1%
#692790000000
0!
0%
#692795000000
1!
1%
#692800000000
0!
0%
#692805000000
1!
1%
#692810000000
0!
0%
#692815000000
1!
1%
#692820000000
0!
0%
#692825000000
1!
1%
#692830000000
0!
0%
#692835000000
1!
1%
#692840000000
0!
0%
#692845000000
1!
1%
#692850000000
0!
0%
#692855000000
1!
1%
#692860000000
0!
0%
#692865000000
1!
1%
#692870000000
0!
0%
#692875000000
1!
1%
#692880000000
0!
0%
#692885000000
1!
1%
#692890000000
0!
0%
#692895000000
1!
1%
#692900000000
0!
0%
#692905000000
1!
1%
#692910000000
0!
0%
#692915000000
1!
1%
#692920000000
0!
0%
#692925000000
1!
1%
#692930000000
0!
0%
#692935000000
1!
1%
#692940000000
0!
0%
#692945000000
1!
1%
#692950000000
0!
0%
#692955000000
1!
1%
#692960000000
0!
0%
#692965000000
1!
1%
#692970000000
0!
0%
#692975000000
1!
1%
#692980000000
0!
0%
#692985000000
1!
1%
#692990000000
0!
0%
#692995000000
1!
1%
#693000000000
0!
0%
#693005000000
1!
1%
#693010000000
0!
0%
#693015000000
1!
1%
#693020000000
0!
0%
#693025000000
1!
1%
#693030000000
0!
0%
#693035000000
1!
1%
#693040000000
0!
0%
#693045000000
1!
1%
#693050000000
0!
0%
#693055000000
1!
1%
#693060000000
0!
0%
#693065000000
1!
1%
#693070000000
0!
0%
#693075000000
1!
1%
#693080000000
0!
0%
#693085000000
1!
1%
#693090000000
0!
0%
#693095000000
1!
1%
#693100000000
0!
0%
#693105000000
1!
1%
#693110000000
0!
0%
#693115000000
1!
1%
#693120000000
0!
0%
#693125000000
1!
1%
#693130000000
0!
0%
#693135000000
1!
1%
#693140000000
0!
0%
#693145000000
1!
1%
#693150000000
0!
0%
#693155000000
1!
1%
#693160000000
0!
0%
#693165000000
1!
1%
#693170000000
0!
0%
#693175000000
1!
1%
#693180000000
0!
0%
#693185000000
1!
1%
#693190000000
0!
0%
#693195000000
1!
1%
#693200000000
0!
0%
#693205000000
1!
1%
#693210000000
0!
0%
#693215000000
1!
1%
#693220000000
0!
0%
#693225000000
1!
1%
#693230000000
0!
0%
#693235000000
1!
1%
#693240000000
0!
0%
#693245000000
1!
1%
#693250000000
0!
0%
#693255000000
1!
1%
#693260000000
0!
0%
#693265000000
1!
1%
#693270000000
0!
0%
#693275000000
1!
1%
#693280000000
0!
0%
#693285000000
1!
1%
#693290000000
0!
0%
#693295000000
1!
1%
#693300000000
0!
0%
#693305000000
1!
1%
#693310000000
0!
0%
#693315000000
1!
1%
#693320000000
0!
0%
#693325000000
1!
1%
#693330000000
0!
0%
#693335000000
1!
1%
#693340000000
0!
0%
#693345000000
1!
1%
#693350000000
0!
0%
#693355000000
1!
1%
#693360000000
0!
0%
#693365000000
1!
1%
#693370000000
0!
0%
#693375000000
1!
1%
#693380000000
0!
0%
#693385000000
1!
1%
#693390000000
0!
0%
#693395000000
1!
1%
#693400000000
0!
0%
#693405000000
1!
1%
#693410000000
0!
0%
#693415000000
1!
1%
#693420000000
0!
0%
#693425000000
1!
1%
#693430000000
0!
0%
#693435000000
1!
1%
#693440000000
0!
0%
#693445000000
1!
1%
#693450000000
0!
0%
#693455000000
1!
1%
#693460000000
0!
0%
#693465000000
1!
1%
#693470000000
0!
0%
#693475000000
1!
1%
#693480000000
0!
0%
#693485000000
1!
1%
#693490000000
0!
0%
#693495000000
1!
1%
#693500000000
0!
0%
#693505000000
1!
1%
#693510000000
0!
0%
#693515000000
1!
1%
#693520000000
0!
0%
#693525000000
1!
1%
#693530000000
0!
0%
#693535000000
1!
1%
#693540000000
0!
0%
#693545000000
1!
1%
#693550000000
0!
0%
#693555000000
1!
1%
#693560000000
0!
0%
#693565000000
1!
1%
#693570000000
0!
0%
#693575000000
1!
1%
#693580000000
0!
0%
#693585000000
1!
1%
#693590000000
0!
0%
#693595000000
1!
1%
#693600000000
0!
0%
#693605000000
1!
1%
#693610000000
0!
0%
#693615000000
1!
1%
#693620000000
0!
0%
#693625000000
1!
1%
#693630000000
0!
0%
#693635000000
1!
1%
#693640000000
0!
0%
#693645000000
1!
1%
#693650000000
0!
0%
#693655000000
1!
1%
#693660000000
0!
0%
#693665000000
1!
1%
#693670000000
0!
0%
#693675000000
1!
1%
#693680000000
0!
0%
#693685000000
1!
1%
#693690000000
0!
0%
#693695000000
1!
1%
#693700000000
0!
0%
#693705000000
1!
1%
#693710000000
0!
0%
#693715000000
1!
1%
#693720000000
0!
0%
#693725000000
1!
1%
#693730000000
0!
0%
#693735000000
1!
1%
#693740000000
0!
0%
#693745000000
1!
1%
#693750000000
0!
0%
#693755000000
1!
1%
#693760000000
0!
0%
#693765000000
1!
1%
#693770000000
0!
0%
#693775000000
1!
1%
#693780000000
0!
0%
#693785000000
1!
1%
#693790000000
0!
0%
#693795000000
1!
1%
#693800000000
0!
0%
#693805000000
1!
1%
#693810000000
0!
0%
#693815000000
1!
1%
#693820000000
0!
0%
#693825000000
1!
1%
#693830000000
0!
0%
#693835000000
1!
1%
#693840000000
0!
0%
#693845000000
1!
1%
#693850000000
0!
0%
#693855000000
1!
1%
#693860000000
0!
0%
#693865000000
1!
1%
#693870000000
0!
0%
#693875000000
1!
1%
#693880000000
0!
0%
#693885000000
1!
1%
#693890000000
0!
0%
#693895000000
1!
1%
#693900000000
0!
0%
#693905000000
1!
1%
#693910000000
0!
0%
#693915000000
1!
1%
#693920000000
0!
0%
#693925000000
1!
1%
#693930000000
0!
0%
#693935000000
1!
1%
#693940000000
0!
0%
#693945000000
1!
1%
#693950000000
0!
0%
#693955000000
1!
1%
#693960000000
0!
0%
#693965000000
1!
1%
#693970000000
0!
0%
#693975000000
1!
1%
#693980000000
0!
0%
#693985000000
1!
1%
#693990000000
0!
0%
#693995000000
1!
1%
#694000000000
0!
0%
#694005000000
1!
1%
#694010000000
0!
0%
#694015000000
1!
1%
#694020000000
0!
0%
#694025000000
1!
1%
#694030000000
0!
0%
#694035000000
1!
1%
#694040000000
0!
0%
#694045000000
1!
1%
#694050000000
0!
0%
#694055000000
1!
1%
#694060000000
0!
0%
#694065000000
1!
1%
#694070000000
0!
0%
#694075000000
1!
1%
#694080000000
0!
0%
#694085000000
1!
1%
#694090000000
0!
0%
#694095000000
1!
1%
#694100000000
0!
0%
#694105000000
1!
1%
#694110000000
0!
0%
#694115000000
1!
1%
#694120000000
0!
0%
#694125000000
1!
1%
#694130000000
0!
0%
#694135000000
1!
1%
#694140000000
0!
0%
#694145000000
1!
1%
#694150000000
0!
0%
#694155000000
1!
1%
#694160000000
0!
0%
#694165000000
1!
1%
#694170000000
0!
0%
#694175000000
1!
1%
#694180000000
0!
0%
#694185000000
1!
1%
#694190000000
0!
0%
#694195000000
1!
1%
#694200000000
0!
0%
#694205000000
1!
1%
#694210000000
0!
0%
#694215000000
1!
1%
#694220000000
0!
0%
#694225000000
1!
1%
#694230000000
0!
0%
#694235000000
1!
1%
#694240000000
0!
0%
#694245000000
1!
1%
#694250000000
0!
0%
#694255000000
1!
1%
#694260000000
0!
0%
#694265000000
1!
1%
#694270000000
0!
0%
#694275000000
1!
1%
#694280000000
0!
0%
#694285000000
1!
1%
#694290000000
0!
0%
#694295000000
1!
1%
#694300000000
0!
0%
#694305000000
1!
1%
#694310000000
0!
0%
#694315000000
1!
1%
#694320000000
0!
0%
#694325000000
1!
1%
#694330000000
0!
0%
#694335000000
1!
1%
#694340000000
0!
0%
#694345000000
1!
1%
#694350000000
0!
0%
#694355000000
1!
1%
#694360000000
0!
0%
#694365000000
1!
1%
#694370000000
0!
0%
#694375000000
1!
1%
#694380000000
0!
0%
#694385000000
1!
1%
#694390000000
0!
0%
#694395000000
1!
1%
#694400000000
0!
0%
#694405000000
1!
1%
#694410000000
0!
0%
#694415000000
1!
1%
#694420000000
0!
0%
#694425000000
1!
1%
#694430000000
0!
0%
#694435000000
1!
1%
#694440000000
0!
0%
#694445000000
1!
1%
#694450000000
0!
0%
#694455000000
1!
1%
#694460000000
0!
0%
#694465000000
1!
1%
#694470000000
0!
0%
#694475000000
1!
1%
#694480000000
0!
0%
#694485000000
1!
1%
#694490000000
0!
0%
#694495000000
1!
1%
#694500000000
0!
0%
#694505000000
1!
1%
#694510000000
0!
0%
#694515000000
1!
1%
#694520000000
0!
0%
#694525000000
1!
1%
#694530000000
0!
0%
#694535000000
1!
1%
#694540000000
0!
0%
#694545000000
1!
1%
#694550000000
0!
0%
#694555000000
1!
1%
#694560000000
0!
0%
#694565000000
1!
1%
#694570000000
0!
0%
#694575000000
1!
1%
#694580000000
0!
0%
#694585000000
1!
1%
#694590000000
0!
0%
#694595000000
1!
1%
#694600000000
0!
0%
#694605000000
1!
1%
#694610000000
0!
0%
#694615000000
1!
1%
#694620000000
0!
0%
#694625000000
1!
1%
#694630000000
0!
0%
#694635000000
1!
1%
#694640000000
0!
0%
#694645000000
1!
1%
#694650000000
0!
0%
#694655000000
1!
1%
#694660000000
0!
0%
#694665000000
1!
1%
#694670000000
0!
0%
#694675000000
1!
1%
#694680000000
0!
0%
#694685000000
1!
1%
#694690000000
0!
0%
#694695000000
1!
1%
#694700000000
0!
0%
#694705000000
1!
1%
#694710000000
0!
0%
#694715000000
1!
1%
#694720000000
0!
0%
#694725000000
1!
1%
#694730000000
0!
0%
#694735000000
1!
1%
#694740000000
0!
0%
#694745000000
1!
1%
#694750000000
0!
0%
#694755000000
1!
1%
#694760000000
0!
0%
#694765000000
1!
1%
#694770000000
0!
0%
#694775000000
1!
1%
#694780000000
0!
0%
#694785000000
1!
1%
#694790000000
0!
0%
#694795000000
1!
1%
#694800000000
0!
0%
#694805000000
1!
1%
#694810000000
0!
0%
#694815000000
1!
1%
#694820000000
0!
0%
#694825000000
1!
1%
#694830000000
0!
0%
#694835000000
1!
1%
#694840000000
0!
0%
#694845000000
1!
1%
#694850000000
0!
0%
#694855000000
1!
1%
#694860000000
0!
0%
#694865000000
1!
1%
#694870000000
0!
0%
#694875000000
1!
1%
#694880000000
0!
0%
#694885000000
1!
1%
#694890000000
0!
0%
#694895000000
1!
1%
#694900000000
0!
0%
#694905000000
1!
1%
#694910000000
0!
0%
#694915000000
1!
1%
#694920000000
0!
0%
#694925000000
1!
1%
#694930000000
0!
0%
#694935000000
1!
1%
#694940000000
0!
0%
#694945000000
1!
1%
#694950000000
0!
0%
#694955000000
1!
1%
#694960000000
0!
0%
#694965000000
1!
1%
#694970000000
0!
0%
#694975000000
1!
1%
#694980000000
0!
0%
#694985000000
1!
1%
#694990000000
0!
0%
#694995000000
1!
1%
#695000000000
0!
0%
#695005000000
1!
1%
#695010000000
0!
0%
#695015000000
1!
1%
#695020000000
0!
0%
#695025000000
1!
1%
#695030000000
0!
0%
#695035000000
1!
1%
#695040000000
0!
0%
#695045000000
1!
1%
#695050000000
0!
0%
#695055000000
1!
1%
#695060000000
0!
0%
#695065000000
1!
1%
#695070000000
0!
0%
#695075000000
1!
1%
#695080000000
0!
0%
#695085000000
1!
1%
#695090000000
0!
0%
#695095000000
1!
1%
#695100000000
0!
0%
#695105000000
1!
1%
#695110000000
0!
0%
#695115000000
1!
1%
#695120000000
0!
0%
#695125000000
1!
1%
#695130000000
0!
0%
#695135000000
1!
1%
#695140000000
0!
0%
#695145000000
1!
1%
#695150000000
0!
0%
#695155000000
1!
1%
#695160000000
0!
0%
#695165000000
1!
1%
#695170000000
0!
0%
#695175000000
1!
1%
#695180000000
0!
0%
#695185000000
1!
1%
#695190000000
0!
0%
#695195000000
1!
1%
#695200000000
0!
0%
#695205000000
1!
1%
#695210000000
0!
0%
#695215000000
1!
1%
#695220000000
0!
0%
#695225000000
1!
1%
#695230000000
0!
0%
#695235000000
1!
1%
#695240000000
0!
0%
#695245000000
1!
1%
#695250000000
0!
0%
#695255000000
1!
1%
#695260000000
0!
0%
#695265000000
1!
1%
#695270000000
0!
0%
#695275000000
1!
1%
#695280000000
0!
0%
#695285000000
1!
1%
#695290000000
0!
0%
#695295000000
1!
1%
#695300000000
0!
0%
#695305000000
1!
1%
#695310000000
0!
0%
#695315000000
1!
1%
#695320000000
0!
0%
#695325000000
1!
1%
#695330000000
0!
0%
#695335000000
1!
1%
#695340000000
0!
0%
#695345000000
1!
1%
#695350000000
0!
0%
#695355000000
1!
1%
#695360000000
0!
0%
#695365000000
1!
1%
#695370000000
0!
0%
#695375000000
1!
1%
#695380000000
0!
0%
#695385000000
1!
1%
#695390000000
0!
0%
#695395000000
1!
1%
#695400000000
0!
0%
#695405000000
1!
1%
#695410000000
0!
0%
#695415000000
1!
1%
#695420000000
0!
0%
#695425000000
1!
1%
#695430000000
0!
0%
#695435000000
1!
1%
#695440000000
0!
0%
#695445000000
1!
1%
#695450000000
0!
0%
#695455000000
1!
1%
#695460000000
0!
0%
#695465000000
1!
1%
#695470000000
0!
0%
#695475000000
1!
1%
#695480000000
0!
0%
#695485000000
1!
1%
#695490000000
0!
0%
#695495000000
1!
1%
#695500000000
0!
0%
#695505000000
1!
1%
#695510000000
0!
0%
#695515000000
1!
1%
#695520000000
0!
0%
#695525000000
1!
1%
#695530000000
0!
0%
#695535000000
1!
1%
#695540000000
0!
0%
#695545000000
1!
1%
#695550000000
0!
0%
#695555000000
1!
1%
#695560000000
0!
0%
#695565000000
1!
1%
#695570000000
0!
0%
#695575000000
1!
1%
#695580000000
0!
0%
#695585000000
1!
1%
#695590000000
0!
0%
#695595000000
1!
1%
#695600000000
0!
0%
#695605000000
1!
1%
#695610000000
0!
0%
#695615000000
1!
1%
#695620000000
0!
0%
#695625000000
1!
1%
#695630000000
0!
0%
#695635000000
1!
1%
#695640000000
0!
0%
#695645000000
1!
1%
#695650000000
0!
0%
#695655000000
1!
1%
#695660000000
0!
0%
#695665000000
1!
1%
#695670000000
0!
0%
#695675000000
1!
1%
#695680000000
0!
0%
#695685000000
1!
1%
#695690000000
0!
0%
#695695000000
1!
1%
#695700000000
0!
0%
#695705000000
1!
1%
#695710000000
0!
0%
#695715000000
1!
1%
#695720000000
0!
0%
#695725000000
1!
1%
#695730000000
0!
0%
#695735000000
1!
1%
#695740000000
0!
0%
#695745000000
1!
1%
#695750000000
0!
0%
#695755000000
1!
1%
#695760000000
0!
0%
#695765000000
1!
1%
#695770000000
0!
0%
#695775000000
1!
1%
#695780000000
0!
0%
#695785000000
1!
1%
#695790000000
0!
0%
#695795000000
1!
1%
#695800000000
0!
0%
#695805000000
1!
1%
#695810000000
0!
0%
#695815000000
1!
1%
#695820000000
0!
0%
#695825000000
1!
1%
#695830000000
0!
0%
#695835000000
1!
1%
#695840000000
0!
0%
#695845000000
1!
1%
#695850000000
0!
0%
#695855000000
1!
1%
#695860000000
0!
0%
#695865000000
1!
1%
#695870000000
0!
0%
#695875000000
1!
1%
#695880000000
0!
0%
#695885000000
1!
1%
#695890000000
0!
0%
#695895000000
1!
1%
#695900000000
0!
0%
#695905000000
1!
1%
#695910000000
0!
0%
#695915000000
1!
1%
#695920000000
0!
0%
#695925000000
1!
1%
#695930000000
0!
0%
#695935000000
1!
1%
#695940000000
0!
0%
#695945000000
1!
1%
#695950000000
0!
0%
#695955000000
1!
1%
#695960000000
0!
0%
#695965000000
1!
1%
#695970000000
0!
0%
#695975000000
1!
1%
#695980000000
0!
0%
#695985000000
1!
1%
#695990000000
0!
0%
#695995000000
1!
1%
#696000000000
0!
0%
#696005000000
1!
1%
#696010000000
0!
0%
#696015000000
1!
1%
#696020000000
0!
0%
#696025000000
1!
1%
#696030000000
0!
0%
#696035000000
1!
1%
#696040000000
0!
0%
#696045000000
1!
1%
#696050000000
0!
0%
#696055000000
1!
1%
#696060000000
0!
0%
#696065000000
1!
1%
#696070000000
0!
0%
#696075000000
1!
1%
#696080000000
0!
0%
#696085000000
1!
1%
#696090000000
0!
0%
#696095000000
1!
1%
#696100000000
0!
0%
#696105000000
1!
1%
#696110000000
0!
0%
#696115000000
1!
1%
#696120000000
0!
0%
#696125000000
1!
1%
#696130000000
0!
0%
#696135000000
1!
1%
#696140000000
0!
0%
#696145000000
1!
1%
#696150000000
0!
0%
#696155000000
1!
1%
#696160000000
0!
0%
#696165000000
1!
1%
#696170000000
0!
0%
#696175000000
1!
1%
#696180000000
0!
0%
#696185000000
1!
1%
#696190000000
0!
0%
#696195000000
1!
1%
#696200000000
0!
0%
#696205000000
1!
1%
#696210000000
0!
0%
#696215000000
1!
1%
#696220000000
0!
0%
#696225000000
1!
1%
#696230000000
0!
0%
#696235000000
1!
1%
#696240000000
0!
0%
#696245000000
1!
1%
#696250000000
0!
0%
#696255000000
1!
1%
#696260000000
0!
0%
#696265000000
1!
1%
#696270000000
0!
0%
#696275000000
1!
1%
#696280000000
0!
0%
#696285000000
1!
1%
#696290000000
0!
0%
#696295000000
1!
1%
#696300000000
0!
0%
#696305000000
1!
1%
#696310000000
0!
0%
#696315000000
1!
1%
#696320000000
0!
0%
#696325000000
1!
1%
#696330000000
0!
0%
#696335000000
1!
1%
#696340000000
0!
0%
#696345000000
1!
1%
#696350000000
0!
0%
#696355000000
1!
1%
#696360000000
0!
0%
#696365000000
1!
1%
#696370000000
0!
0%
#696375000000
1!
1%
#696380000000
0!
0%
#696385000000
1!
1%
#696390000000
0!
0%
#696395000000
1!
1%
#696400000000
0!
0%
#696405000000
1!
1%
#696410000000
0!
0%
#696415000000
1!
1%
#696420000000
0!
0%
#696425000000
1!
1%
#696430000000
0!
0%
#696435000000
1!
1%
#696440000000
0!
0%
#696445000000
1!
1%
#696450000000
0!
0%
#696455000000
1!
1%
#696460000000
0!
0%
#696465000000
1!
1%
#696470000000
0!
0%
#696475000000
1!
1%
#696480000000
0!
0%
#696485000000
1!
1%
#696490000000
0!
0%
#696495000000
1!
1%
#696500000000
0!
0%
#696505000000
1!
1%
#696510000000
0!
0%
#696515000000
1!
1%
#696520000000
0!
0%
#696525000000
1!
1%
#696530000000
0!
0%
#696535000000
1!
1%
#696540000000
0!
0%
#696545000000
1!
1%
#696550000000
0!
0%
#696555000000
1!
1%
#696560000000
0!
0%
#696565000000
1!
1%
#696570000000
0!
0%
#696575000000
1!
1%
#696580000000
0!
0%
#696585000000
1!
1%
#696590000000
0!
0%
#696595000000
1!
1%
#696600000000
0!
0%
#696605000000
1!
1%
#696610000000
0!
0%
#696615000000
1!
1%
#696620000000
0!
0%
#696625000000
1!
1%
#696630000000
0!
0%
#696635000000
1!
1%
#696640000000
0!
0%
#696645000000
1!
1%
#696650000000
0!
0%
#696655000000
1!
1%
#696660000000
0!
0%
#696665000000
1!
1%
#696670000000
0!
0%
#696675000000
1!
1%
#696680000000
0!
0%
#696685000000
1!
1%
#696690000000
0!
0%
#696695000000
1!
1%
#696700000000
0!
0%
#696705000000
1!
1%
#696710000000
0!
0%
#696715000000
1!
1%
#696720000000
0!
0%
#696725000000
1!
1%
#696730000000
0!
0%
#696735000000
1!
1%
#696740000000
0!
0%
#696745000000
1!
1%
#696750000000
0!
0%
#696755000000
1!
1%
#696760000000
0!
0%
#696765000000
1!
1%
#696770000000
0!
0%
#696775000000
1!
1%
#696780000000
0!
0%
#696785000000
1!
1%
#696790000000
0!
0%
#696795000000
1!
1%
#696800000000
0!
0%
#696805000000
1!
1%
#696810000000
0!
0%
#696815000000
1!
1%
#696820000000
0!
0%
#696825000000
1!
1%
#696830000000
0!
0%
#696835000000
1!
1%
#696840000000
0!
0%
#696845000000
1!
1%
#696850000000
0!
0%
#696855000000
1!
1%
#696860000000
0!
0%
#696865000000
1!
1%
#696870000000
0!
0%
#696875000000
1!
1%
#696880000000
0!
0%
#696885000000
1!
1%
#696890000000
0!
0%
#696895000000
1!
1%
#696900000000
0!
0%
#696905000000
1!
1%
#696910000000
0!
0%
#696915000000
1!
1%
#696920000000
0!
0%
#696925000000
1!
1%
#696930000000
0!
0%
#696935000000
1!
1%
#696940000000
0!
0%
#696945000000
1!
1%
#696950000000
0!
0%
#696955000000
1!
1%
#696960000000
0!
0%
#696965000000
1!
1%
#696970000000
0!
0%
#696975000000
1!
1%
#696980000000
0!
0%
#696985000000
1!
1%
#696990000000
0!
0%
#696995000000
1!
1%
#697000000000
0!
0%
#697005000000
1!
1%
#697010000000
0!
0%
#697015000000
1!
1%
#697020000000
0!
0%
#697025000000
1!
1%
#697030000000
0!
0%
#697035000000
1!
1%
#697040000000
0!
0%
#697045000000
1!
1%
#697050000000
0!
0%
#697055000000
1!
1%
#697060000000
0!
0%
#697065000000
1!
1%
#697070000000
0!
0%
#697075000000
1!
1%
#697080000000
0!
0%
#697085000000
1!
1%
#697090000000
0!
0%
#697095000000
1!
1%
#697100000000
0!
0%
#697105000000
1!
1%
#697110000000
0!
0%
#697115000000
1!
1%
#697120000000
0!
0%
#697125000000
1!
1%
#697130000000
0!
0%
#697135000000
1!
1%
#697140000000
0!
0%
#697145000000
1!
1%
#697150000000
0!
0%
#697155000000
1!
1%
#697160000000
0!
0%
#697165000000
1!
1%
#697170000000
0!
0%
#697175000000
1!
1%
#697180000000
0!
0%
#697185000000
1!
1%
#697190000000
0!
0%
#697195000000
1!
1%
#697200000000
0!
0%
#697205000000
1!
1%
#697210000000
0!
0%
#697215000000
1!
1%
#697220000000
0!
0%
#697225000000
1!
1%
#697230000000
0!
0%
#697235000000
1!
1%
#697240000000
0!
0%
#697245000000
1!
1%
#697250000000
0!
0%
#697255000000
1!
1%
#697260000000
0!
0%
#697265000000
1!
1%
#697270000000
0!
0%
#697275000000
1!
1%
#697280000000
0!
0%
#697285000000
1!
1%
#697290000000
0!
0%
#697295000000
1!
1%
#697300000000
0!
0%
#697305000000
1!
1%
#697310000000
0!
0%
#697315000000
1!
1%
#697320000000
0!
0%
#697325000000
1!
1%
#697330000000
0!
0%
#697335000000
1!
1%
#697340000000
0!
0%
#697345000000
1!
1%
#697350000000
0!
0%
#697355000000
1!
1%
#697360000000
0!
0%
#697365000000
1!
1%
#697370000000
0!
0%
#697375000000
1!
1%
#697380000000
0!
0%
#697385000000
1!
1%
#697390000000
0!
0%
#697395000000
1!
1%
#697400000000
0!
0%
#697405000000
1!
1%
#697410000000
0!
0%
#697415000000
1!
1%
#697420000000
0!
0%
#697425000000
1!
1%
#697430000000
0!
0%
#697435000000
1!
1%
#697440000000
0!
0%
#697445000000
1!
1%
#697450000000
0!
0%
#697455000000
1!
1%
#697460000000
0!
0%
#697465000000
1!
1%
#697470000000
0!
0%
#697475000000
1!
1%
#697480000000
0!
0%
#697485000000
1!
1%
#697490000000
0!
0%
#697495000000
1!
1%
#697500000000
0!
0%
#697505000000
1!
1%
#697510000000
0!
0%
#697515000000
1!
1%
#697520000000
0!
0%
#697525000000
1!
1%
#697530000000
0!
0%
#697535000000
1!
1%
#697540000000
0!
0%
#697545000000
1!
1%
#697550000000
0!
0%
#697555000000
1!
1%
#697560000000
0!
0%
#697565000000
1!
1%
#697570000000
0!
0%
#697575000000
1!
1%
#697580000000
0!
0%
#697585000000
1!
1%
#697590000000
0!
0%
#697595000000
1!
1%
#697600000000
0!
0%
#697605000000
1!
1%
#697610000000
0!
0%
#697615000000
1!
1%
#697620000000
0!
0%
#697625000000
1!
1%
#697630000000
0!
0%
#697635000000
1!
1%
#697640000000
0!
0%
#697645000000
1!
1%
#697650000000
0!
0%
#697655000000
1!
1%
#697660000000
0!
0%
#697665000000
1!
1%
#697670000000
0!
0%
#697675000000
1!
1%
#697680000000
0!
0%
#697685000000
1!
1%
#697690000000
0!
0%
#697695000000
1!
1%
#697700000000
0!
0%
#697705000000
1!
1%
#697710000000
0!
0%
#697715000000
1!
1%
#697720000000
0!
0%
#697725000000
1!
1%
#697730000000
0!
0%
#697735000000
1!
1%
#697740000000
0!
0%
#697745000000
1!
1%
#697750000000
0!
0%
#697755000000
1!
1%
#697760000000
0!
0%
#697765000000
1!
1%
#697770000000
0!
0%
#697775000000
1!
1%
#697780000000
0!
0%
#697785000000
1!
1%
#697790000000
0!
0%
#697795000000
1!
1%
#697800000000
0!
0%
#697805000000
1!
1%
#697810000000
0!
0%
#697815000000
1!
1%
#697820000000
0!
0%
#697825000000
1!
1%
#697830000000
0!
0%
#697835000000
1!
1%
#697840000000
0!
0%
#697845000000
1!
1%
#697850000000
0!
0%
#697855000000
1!
1%
#697860000000
0!
0%
#697865000000
1!
1%
#697870000000
0!
0%
#697875000000
1!
1%
#697880000000
0!
0%
#697885000000
1!
1%
#697890000000
0!
0%
#697895000000
1!
1%
#697900000000
0!
0%
#697905000000
1!
1%
#697910000000
0!
0%
#697915000000
1!
1%
#697920000000
0!
0%
#697925000000
1!
1%
#697930000000
0!
0%
#697935000000
1!
1%
#697940000000
0!
0%
#697945000000
1!
1%
#697950000000
0!
0%
#697955000000
1!
1%
#697960000000
0!
0%
#697965000000
1!
1%
#697970000000
0!
0%
#697975000000
1!
1%
#697980000000
0!
0%
#697985000000
1!
1%
#697990000000
0!
0%
#697995000000
1!
1%
#698000000000
0!
0%
#698005000000
1!
1%
#698010000000
0!
0%
#698015000000
1!
1%
#698020000000
0!
0%
#698025000000
1!
1%
#698030000000
0!
0%
#698035000000
1!
1%
#698040000000
0!
0%
#698045000000
1!
1%
#698050000000
0!
0%
#698055000000
1!
1%
#698060000000
0!
0%
#698065000000
1!
1%
#698070000000
0!
0%
#698075000000
1!
1%
#698080000000
0!
0%
#698085000000
1!
1%
#698090000000
0!
0%
#698095000000
1!
1%
#698100000000
0!
0%
#698105000000
1!
1%
#698110000000
0!
0%
#698115000000
1!
1%
#698120000000
0!
0%
#698125000000
1!
1%
#698130000000
0!
0%
#698135000000
1!
1%
#698140000000
0!
0%
#698145000000
1!
1%
#698150000000
0!
0%
#698155000000
1!
1%
#698160000000
0!
0%
#698165000000
1!
1%
#698170000000
0!
0%
#698175000000
1!
1%
#698180000000
0!
0%
#698185000000
1!
1%
#698190000000
0!
0%
#698195000000
1!
1%
#698200000000
0!
0%
#698205000000
1!
1%
#698210000000
0!
0%
#698215000000
1!
1%
#698220000000
0!
0%
#698225000000
1!
1%
#698230000000
0!
0%
#698235000000
1!
1%
#698240000000
0!
0%
#698245000000
1!
1%
#698250000000
0!
0%
#698255000000
1!
1%
#698260000000
0!
0%
#698265000000
1!
1%
#698270000000
0!
0%
#698275000000
1!
1%
#698280000000
0!
0%
#698285000000
1!
1%
#698290000000
0!
0%
#698295000000
1!
1%
#698300000000
0!
0%
#698305000000
1!
1%
#698310000000
0!
0%
#698315000000
1!
1%
#698320000000
0!
0%
#698325000000
1!
1%
#698330000000
0!
0%
#698335000000
1!
1%
#698340000000
0!
0%
#698345000000
1!
1%
#698350000000
0!
0%
#698355000000
1!
1%
#698360000000
0!
0%
#698365000000
1!
1%
#698370000000
0!
0%
#698375000000
1!
1%
#698380000000
0!
0%
#698385000000
1!
1%
#698390000000
0!
0%
#698395000000
1!
1%
#698400000000
0!
0%
#698405000000
1!
1%
#698410000000
0!
0%
#698415000000
1!
1%
#698420000000
0!
0%
#698425000000
1!
1%
#698430000000
0!
0%
#698435000000
1!
1%
#698440000000
0!
0%
#698445000000
1!
1%
#698450000000
0!
0%
#698455000000
1!
1%
#698460000000
0!
0%
#698465000000
1!
1%
#698470000000
0!
0%
#698475000000
1!
1%
#698480000000
0!
0%
#698485000000
1!
1%
#698490000000
0!
0%
#698495000000
1!
1%
#698500000000
0!
0%
#698505000000
1!
1%
#698510000000
0!
0%
#698515000000
1!
1%
#698520000000
0!
0%
#698525000000
1!
1%
#698530000000
0!
0%
#698535000000
1!
1%
#698540000000
0!
0%
#698545000000
1!
1%
#698550000000
0!
0%
#698555000000
1!
1%
#698560000000
0!
0%
#698565000000
1!
1%
#698570000000
0!
0%
#698575000000
1!
1%
#698580000000
0!
0%
#698585000000
1!
1%
#698590000000
0!
0%
#698595000000
1!
1%
#698600000000
0!
0%
#698605000000
1!
1%
#698610000000
0!
0%
#698615000000
1!
1%
#698620000000
0!
0%
#698625000000
1!
1%
#698630000000
0!
0%
#698635000000
1!
1%
#698640000000
0!
0%
#698645000000
1!
1%
#698650000000
0!
0%
#698655000000
1!
1%
#698660000000
0!
0%
#698665000000
1!
1%
#698670000000
0!
0%
#698675000000
1!
1%
#698680000000
0!
0%
#698685000000
1!
1%
#698690000000
0!
0%
#698695000000
1!
1%
#698700000000
0!
0%
#698705000000
1!
1%
#698710000000
0!
0%
#698715000000
1!
1%
#698720000000
0!
0%
#698725000000
1!
1%
#698730000000
0!
0%
#698735000000
1!
1%
#698740000000
0!
0%
#698745000000
1!
1%
#698750000000
0!
0%
#698755000000
1!
1%
#698760000000
0!
0%
#698765000000
1!
1%
#698770000000
0!
0%
#698775000000
1!
1%
#698780000000
0!
0%
#698785000000
1!
1%
#698790000000
0!
0%
#698795000000
1!
1%
#698800000000
0!
0%
#698805000000
1!
1%
#698810000000
0!
0%
#698815000000
1!
1%
#698820000000
0!
0%
#698825000000
1!
1%
#698830000000
0!
0%
#698835000000
1!
1%
#698840000000
0!
0%
#698845000000
1!
1%
#698850000000
0!
0%
#698855000000
1!
1%
#698860000000
0!
0%
#698865000000
1!
1%
#698870000000
0!
0%
#698875000000
1!
1%
#698880000000
0!
0%
#698885000000
1!
1%
#698890000000
0!
0%
#698895000000
1!
1%
#698900000000
0!
0%
#698905000000
1!
1%
#698910000000
0!
0%
#698915000000
1!
1%
#698920000000
0!
0%
#698925000000
1!
1%
#698930000000
0!
0%
#698935000000
1!
1%
#698940000000
0!
0%
#698945000000
1!
1%
#698950000000
0!
0%
#698955000000
1!
1%
#698960000000
0!
0%
#698965000000
1!
1%
#698970000000
0!
0%
#698975000000
1!
1%
#698980000000
0!
0%
#698985000000
1!
1%
#698990000000
0!
0%
#698995000000
1!
1%
#699000000000
0!
0%
#699005000000
1!
1%
#699010000000
0!
0%
#699015000000
1!
1%
#699020000000
0!
0%
#699025000000
1!
1%
#699030000000
0!
0%
#699035000000
1!
1%
#699040000000
0!
0%
#699045000000
1!
1%
#699050000000
0!
0%
#699055000000
1!
1%
#699060000000
0!
0%
#699065000000
1!
1%
#699070000000
0!
0%
#699075000000
1!
1%
#699080000000
0!
0%
#699085000000
1!
1%
#699090000000
0!
0%
#699095000000
1!
1%
#699100000000
0!
0%
#699105000000
1!
1%
#699110000000
0!
0%
#699115000000
1!
1%
#699120000000
0!
0%
#699125000000
1!
1%
#699130000000
0!
0%
#699135000000
1!
1%
#699140000000
0!
0%
#699145000000
1!
1%
#699150000000
0!
0%
#699155000000
1!
1%
#699160000000
0!
0%
#699165000000
1!
1%
#699170000000
0!
0%
#699175000000
1!
1%
#699180000000
0!
0%
#699185000000
1!
1%
#699190000000
0!
0%
#699195000000
1!
1%
#699200000000
0!
0%
#699205000000
1!
1%
#699210000000
0!
0%
#699215000000
1!
1%
#699220000000
0!
0%
#699225000000
1!
1%
#699230000000
0!
0%
#699235000000
1!
1%
#699240000000
0!
0%
#699245000000
1!
1%
#699250000000
0!
0%
#699255000000
1!
1%
#699260000000
0!
0%
#699265000000
1!
1%
#699270000000
0!
0%
#699275000000
1!
1%
#699280000000
0!
0%
#699285000000
1!
1%
#699290000000
0!
0%
#699295000000
1!
1%
#699300000000
0!
0%
#699305000000
1!
1%
#699310000000
0!
0%
#699315000000
1!
1%
#699320000000
0!
0%
#699325000000
1!
1%
#699330000000
0!
0%
#699335000000
1!
1%
#699340000000
0!
0%
#699345000000
1!
1%
#699350000000
0!
0%
#699355000000
1!
1%
#699360000000
0!
0%
#699365000000
1!
1%
#699370000000
0!
0%
#699375000000
1!
1%
#699380000000
0!
0%
#699385000000
1!
1%
#699390000000
0!
0%
#699395000000
1!
1%
#699400000000
0!
0%
#699405000000
1!
1%
#699410000000
0!
0%
#699415000000
1!
1%
#699420000000
0!
0%
#699425000000
1!
1%
#699430000000
0!
0%
#699435000000
1!
1%
#699440000000
0!
0%
#699445000000
1!
1%
#699450000000
0!
0%
#699455000000
1!
1%
#699460000000
0!
0%
#699465000000
1!
1%
#699470000000
0!
0%
#699475000000
1!
1%
#699480000000
0!
0%
#699485000000
1!
1%
#699490000000
0!
0%
#699495000000
1!
1%
#699500000000
0!
0%
#699505000000
1!
1%
#699510000000
0!
0%
#699515000000
1!
1%
#699520000000
0!
0%
#699525000000
1!
1%
#699530000000
0!
0%
#699535000000
1!
1%
#699540000000
0!
0%
#699545000000
1!
1%
#699550000000
0!
0%
#699555000000
1!
1%
#699560000000
0!
0%
#699565000000
1!
1%
#699570000000
0!
0%
#699575000000
1!
1%
#699580000000
0!
0%
#699585000000
1!
1%
#699590000000
0!
0%
#699595000000
1!
1%
#699600000000
0!
0%
#699605000000
1!
1%
#699610000000
0!
0%
#699615000000
1!
1%
#699620000000
0!
0%
#699625000000
1!
1%
#699630000000
0!
0%
#699635000000
1!
1%
#699640000000
0!
0%
#699645000000
1!
1%
#699650000000
0!
0%
#699655000000
1!
1%
#699660000000
0!
0%
#699665000000
1!
1%
#699670000000
0!
0%
#699675000000
1!
1%
#699680000000
0!
0%
#699685000000
1!
1%
#699690000000
0!
0%
#699695000000
1!
1%
#699700000000
0!
0%
#699705000000
1!
1%
#699710000000
0!
0%
#699715000000
1!
1%
#699720000000
0!
0%
#699725000000
1!
1%
#699730000000
0!
0%
#699735000000
1!
1%
#699740000000
0!
0%
#699745000000
1!
1%
#699750000000
0!
0%
#699755000000
1!
1%
#699760000000
0!
0%
#699765000000
1!
1%
#699770000000
0!
0%
#699775000000
1!
1%
#699780000000
0!
0%
#699785000000
1!
1%
#699790000000
0!
0%
#699795000000
1!
1%
#699800000000
0!
0%
#699805000000
1!
1%
#699810000000
0!
0%
#699815000000
1!
1%
#699820000000
0!
0%
#699825000000
1!
1%
#699830000000
0!
0%
#699835000000
1!
1%
#699840000000
0!
0%
#699845000000
1!
1%
#699850000000
0!
0%
#699855000000
1!
1%
#699860000000
0!
0%
#699865000000
1!
1%
#699870000000
0!
0%
#699875000000
1!
1%
#699880000000
0!
0%
#699885000000
1!
1%
#699890000000
0!
0%
#699895000000
1!
1%
#699900000000
0!
0%
#699905000000
1!
1%
#699910000000
0!
0%
#699915000000
1!
1%
#699920000000
0!
0%
#699925000000
1!
1%
#699930000000
0!
0%
#699935000000
1!
1%
#699940000000
0!
0%
#699945000000
1!
1%
#699950000000
0!
0%
#699955000000
1!
1%
#699960000000
0!
0%
#699965000000
1!
1%
#699970000000
0!
0%
#699975000000
1!
1%
#699980000000
0!
0%
#699985000000
1!
1%
#699990000000
0!
0%
#699995000000
1!
1%
#700000000000
0!
0%
#700005000000
1!
1%
#700010000000
0!
0%
#700015000000
1!
1%
#700020000000
0!
0%
#700025000000
1!
1%
#700030000000
0!
0%
#700035000000
1!
1%
#700040000000
0!
0%
#700045000000
1!
1%
#700050000000
0!
0%
#700055000000
1!
1%
#700060000000
0!
0%
#700065000000
1!
1%
#700070000000
0!
0%
#700075000000
1!
1%
#700080000000
0!
0%
#700085000000
1!
1%
#700090000000
0!
0%
#700095000000
1!
1%
#700100000000
0!
0%
#700105000000
1!
1%
#700110000000
0!
0%
#700115000000
1!
1%
#700120000000
0!
0%
#700125000000
1!
1%
#700130000000
0!
0%
#700135000000
1!
1%
#700140000000
0!
0%
#700145000000
1!
1%
#700150000000
0!
0%
#700155000000
1!
1%
#700160000000
0!
0%
#700165000000
1!
1%
#700170000000
0!
0%
#700175000000
1!
1%
#700180000000
0!
0%
#700185000000
1!
1%
#700190000000
0!
0%
#700195000000
1!
1%
#700200000000
0!
0%
#700205000000
1!
1%
#700210000000
0!
0%
#700215000000
1!
1%
#700220000000
0!
0%
#700225000000
1!
1%
#700230000000
0!
0%
#700235000000
1!
1%
#700240000000
0!
0%
#700245000000
1!
1%
#700250000000
0!
0%
#700255000000
1!
1%
#700260000000
0!
0%
#700265000000
1!
1%
#700270000000
0!
0%
#700275000000
1!
1%
#700280000000
0!
0%
#700285000000
1!
1%
#700290000000
0!
0%
#700295000000
1!
1%
#700300000000
0!
0%
#700305000000
1!
1%
#700310000000
0!
0%
#700315000000
1!
1%
#700320000000
0!
0%
#700325000000
1!
1%
#700330000000
0!
0%
#700335000000
1!
1%
#700340000000
0!
0%
#700345000000
1!
1%
#700350000000
0!
0%
#700355000000
1!
1%
#700360000000
0!
0%
#700365000000
1!
1%
#700370000000
0!
0%
#700375000000
1!
1%
#700380000000
0!
0%
#700385000000
1!
1%
#700390000000
0!
0%
#700395000000
1!
1%
#700400000000
0!
0%
#700405000000
1!
1%
#700410000000
0!
0%
#700415000000
1!
1%
#700420000000
0!
0%
#700425000000
1!
1%
#700430000000
0!
0%
#700435000000
1!
1%
#700440000000
0!
0%
#700445000000
1!
1%
#700450000000
0!
0%
#700455000000
1!
1%
#700460000000
0!
0%
#700465000000
1!
1%
#700470000000
0!
0%
#700475000000
1!
1%
#700480000000
0!
0%
#700485000000
1!
1%
#700490000000
0!
0%
#700495000000
1!
1%
#700500000000
0!
0%
#700505000000
1!
1%
#700510000000
0!
0%
#700515000000
1!
1%
#700520000000
0!
0%
#700525000000
1!
1%
#700530000000
0!
0%
#700535000000
1!
1%
#700540000000
0!
0%
#700545000000
1!
1%
#700550000000
0!
0%
#700555000000
1!
1%
#700560000000
0!
0%
#700565000000
1!
1%
#700570000000
0!
0%
#700575000000
1!
1%
#700580000000
0!
0%
#700585000000
1!
1%
#700590000000
0!
0%
#700595000000
1!
1%
#700600000000
0!
0%
#700605000000
1!
1%
#700610000000
0!
0%
#700615000000
1!
1%
#700620000000
0!
0%
#700625000000
1!
1%
#700630000000
0!
0%
#700635000000
1!
1%
#700640000000
0!
0%
#700645000000
1!
1%
#700650000000
0!
0%
#700655000000
1!
1%
#700660000000
0!
0%
#700665000000
1!
1%
#700670000000
0!
0%
#700675000000
1!
1%
#700680000000
0!
0%
#700685000000
1!
1%
#700690000000
0!
0%
#700695000000
1!
1%
#700700000000
0!
0%
#700705000000
1!
1%
#700710000000
0!
0%
#700715000000
1!
1%
#700720000000
0!
0%
#700725000000
1!
1%
#700730000000
0!
0%
#700735000000
1!
1%
#700740000000
0!
0%
#700745000000
1!
1%
#700750000000
0!
0%
#700755000000
1!
1%
#700760000000
0!
0%
#700765000000
1!
1%
#700770000000
0!
0%
#700775000000
1!
1%
#700780000000
0!
0%
#700785000000
1!
1%
#700790000000
0!
0%
#700795000000
1!
1%
#700800000000
0!
0%
#700805000000
1!
1%
#700810000000
0!
0%
#700815000000
1!
1%
#700820000000
0!
0%
#700825000000
1!
1%
#700830000000
0!
0%
#700835000000
1!
1%
#700840000000
0!
0%
#700845000000
1!
1%
#700850000000
0!
0%
#700855000000
1!
1%
#700860000000
0!
0%
#700865000000
1!
1%
#700870000000
0!
0%
#700875000000
1!
1%
#700880000000
0!
0%
#700885000000
1!
1%
#700890000000
0!
0%
#700895000000
1!
1%
#700900000000
0!
0%
#700905000000
1!
1%
#700910000000
0!
0%
#700915000000
1!
1%
#700920000000
0!
0%
#700925000000
1!
1%
#700930000000
0!
0%
#700935000000
1!
1%
#700940000000
0!
0%
#700945000000
1!
1%
#700950000000
0!
0%
#700955000000
1!
1%
#700960000000
0!
0%
#700965000000
1!
1%
#700970000000
0!
0%
#700975000000
1!
1%
#700980000000
0!
0%
#700985000000
1!
1%
#700990000000
0!
0%
#700995000000
1!
1%
#701000000000
0!
0%
#701005000000
1!
1%
#701010000000
0!
0%
#701015000000
1!
1%
#701020000000
0!
0%
#701025000000
1!
1%
#701030000000
0!
0%
#701035000000
1!
1%
#701040000000
0!
0%
#701045000000
1!
1%
#701050000000
0!
0%
#701055000000
1!
1%
#701060000000
0!
0%
#701065000000
1!
1%
#701070000000
0!
0%
#701075000000
1!
1%
#701080000000
0!
0%
#701085000000
1!
1%
#701090000000
0!
0%
#701095000000
1!
1%
#701100000000
0!
0%
#701105000000
1!
1%
#701110000000
0!
0%
#701115000000
1!
1%
#701120000000
0!
0%
#701125000000
1!
1%
#701130000000
0!
0%
#701135000000
1!
1%
#701140000000
0!
0%
#701145000000
1!
1%
#701150000000
0!
0%
#701155000000
1!
1%
#701160000000
0!
0%
#701165000000
1!
1%
#701170000000
0!
0%
#701175000000
1!
1%
#701180000000
0!
0%
#701185000000
1!
1%
#701190000000
0!
0%
#701195000000
1!
1%
#701200000000
0!
0%
#701205000000
1!
1%
#701210000000
0!
0%
#701215000000
1!
1%
#701220000000
0!
0%
#701225000000
1!
1%
#701230000000
0!
0%
#701235000000
1!
1%
#701240000000
0!
0%
#701245000000
1!
1%
#701250000000
0!
0%
#701255000000
1!
1%
#701260000000
0!
0%
#701265000000
1!
1%
#701270000000
0!
0%
#701275000000
1!
1%
#701280000000
0!
0%
#701285000000
1!
1%
#701290000000
0!
0%
#701295000000
1!
1%
#701300000000
0!
0%
#701305000000
1!
1%
#701310000000
0!
0%
#701315000000
1!
1%
#701320000000
0!
0%
#701325000000
1!
1%
#701330000000
0!
0%
#701335000000
1!
1%
#701340000000
0!
0%
#701345000000
1!
1%
#701350000000
0!
0%
#701355000000
1!
1%
#701360000000
0!
0%
#701365000000
1!
1%
#701370000000
0!
0%
#701375000000
1!
1%
#701380000000
0!
0%
#701385000000
1!
1%
#701390000000
0!
0%
#701395000000
1!
1%
#701400000000
0!
0%
#701405000000
1!
1%
#701410000000
0!
0%
#701415000000
1!
1%
#701420000000
0!
0%
#701425000000
1!
1%
#701430000000
0!
0%
#701435000000
1!
1%
#701440000000
0!
0%
#701445000000
1!
1%
#701450000000
0!
0%
#701455000000
1!
1%
#701460000000
0!
0%
#701465000000
1!
1%
#701470000000
0!
0%
#701475000000
1!
1%
#701480000000
0!
0%
#701485000000
1!
1%
#701490000000
0!
0%
#701495000000
1!
1%
#701500000000
0!
0%
#701505000000
1!
1%
#701510000000
0!
0%
#701515000000
1!
1%
#701520000000
0!
0%
#701525000000
1!
1%
#701530000000
0!
0%
#701535000000
1!
1%
#701540000000
0!
0%
#701545000000
1!
1%
#701550000000
0!
0%
#701555000000
1!
1%
#701560000000
0!
0%
#701565000000
1!
1%
#701570000000
0!
0%
#701575000000
1!
1%
#701580000000
0!
0%
#701585000000
1!
1%
#701590000000
0!
0%
#701595000000
1!
1%
#701600000000
0!
0%
#701605000000
1!
1%
#701610000000
0!
0%
#701615000000
1!
1%
#701620000000
0!
0%
#701625000000
1!
1%
#701630000000
0!
0%
#701635000000
1!
1%
#701640000000
0!
0%
#701645000000
1!
1%
#701650000000
0!
0%
#701655000000
1!
1%
#701660000000
0!
0%
#701665000000
1!
1%
#701670000000
0!
0%
#701675000000
1!
1%
#701680000000
0!
0%
#701685000000
1!
1%
#701690000000
0!
0%
#701695000000
1!
1%
#701700000000
0!
0%
#701705000000
1!
1%
#701710000000
0!
0%
#701715000000
1!
1%
#701720000000
0!
0%
#701725000000
1!
1%
#701730000000
0!
0%
#701735000000
1!
1%
#701740000000
0!
0%
#701745000000
1!
1%
#701750000000
0!
0%
#701755000000
1!
1%
#701760000000
0!
0%
#701765000000
1!
1%
#701770000000
0!
0%
#701775000000
1!
1%
#701780000000
0!
0%
#701785000000
1!
1%
#701790000000
0!
0%
#701795000000
1!
1%
#701800000000
0!
0%
#701805000000
1!
1%
#701810000000
0!
0%
#701815000000
1!
1%
#701820000000
0!
0%
#701825000000
1!
1%
#701830000000
0!
0%
#701835000000
1!
1%
#701840000000
0!
0%
#701845000000
1!
1%
#701850000000
0!
0%
#701855000000
1!
1%
#701860000000
0!
0%
#701865000000
1!
1%
#701870000000
0!
0%
#701875000000
1!
1%
#701880000000
0!
0%
#701885000000
1!
1%
#701890000000
0!
0%
#701895000000
1!
1%
#701900000000
0!
0%
#701905000000
1!
1%
#701910000000
0!
0%
#701915000000
1!
1%
#701920000000
0!
0%
#701925000000
1!
1%
#701930000000
0!
0%
#701935000000
1!
1%
#701940000000
0!
0%
#701945000000
1!
1%
#701950000000
0!
0%
#701955000000
1!
1%
#701960000000
0!
0%
#701965000000
1!
1%
#701970000000
0!
0%
#701975000000
1!
1%
#701980000000
0!
0%
#701985000000
1!
1%
#701990000000
0!
0%
#701995000000
1!
1%
#702000000000
0!
0%
#702005000000
1!
1%
#702010000000
0!
0%
#702015000000
1!
1%
#702020000000
0!
0%
#702025000000
1!
1%
#702030000000
0!
0%
#702035000000
1!
1%
#702040000000
0!
0%
#702045000000
1!
1%
#702050000000
0!
0%
#702055000000
1!
1%
#702060000000
0!
0%
#702065000000
1!
1%
#702070000000
0!
0%
#702075000000
1!
1%
#702080000000
0!
0%
#702085000000
1!
1%
#702090000000
0!
0%
#702095000000
1!
1%
#702100000000
0!
0%
#702105000000
1!
1%
#702110000000
0!
0%
#702115000000
1!
1%
#702120000000
0!
0%
#702125000000
1!
1%
#702130000000
0!
0%
#702135000000
1!
1%
#702140000000
0!
0%
#702145000000
1!
1%
#702150000000
0!
0%
#702155000000
1!
1%
#702160000000
0!
0%
#702165000000
1!
1%
#702170000000
0!
0%
#702175000000
1!
1%
#702180000000
0!
0%
#702185000000
1!
1%
#702190000000
0!
0%
#702195000000
1!
1%
#702200000000
0!
0%
#702205000000
1!
1%
#702210000000
0!
0%
#702215000000
1!
1%
#702220000000
0!
0%
#702225000000
1!
1%
#702230000000
0!
0%
#702235000000
1!
1%
#702240000000
0!
0%
#702245000000
1!
1%
#702250000000
0!
0%
#702255000000
1!
1%
#702260000000
0!
0%
#702265000000
1!
1%
#702270000000
0!
0%
#702275000000
1!
1%
#702280000000
0!
0%
#702285000000
1!
1%
#702290000000
0!
0%
#702295000000
1!
1%
#702300000000
0!
0%
#702305000000
1!
1%
#702310000000
0!
0%
#702315000000
1!
1%
#702320000000
0!
0%
#702325000000
1!
1%
#702330000000
0!
0%
#702335000000
1!
1%
#702340000000
0!
0%
#702345000000
1!
1%
#702350000000
0!
0%
#702355000000
1!
1%
#702360000000
0!
0%
#702365000000
1!
1%
#702370000000
0!
0%
#702375000000
1!
1%
#702380000000
0!
0%
#702385000000
1!
1%
#702390000000
0!
0%
#702395000000
1!
1%
#702400000000
0!
0%
#702405000000
1!
1%
#702410000000
0!
0%
#702415000000
1!
1%
#702420000000
0!
0%
#702425000000
1!
1%
#702430000000
0!
0%
#702435000000
1!
1%
#702440000000
0!
0%
#702445000000
1!
1%
#702450000000
0!
0%
#702455000000
1!
1%
#702460000000
0!
0%
#702465000000
1!
1%
#702470000000
0!
0%
#702475000000
1!
1%
#702480000000
0!
0%
#702485000000
1!
1%
#702490000000
0!
0%
#702495000000
1!
1%
#702500000000
0!
0%
#702505000000
1!
1%
#702510000000
0!
0%
#702515000000
1!
1%
#702520000000
0!
0%
#702525000000
1!
1%
#702530000000
0!
0%
#702535000000
1!
1%
#702540000000
0!
0%
#702545000000
1!
1%
#702550000000
0!
0%
#702555000000
1!
1%
#702560000000
0!
0%
#702565000000
1!
1%
#702570000000
0!
0%
#702575000000
1!
1%
#702580000000
0!
0%
#702585000000
1!
1%
#702590000000
0!
0%
#702595000000
1!
1%
#702600000000
0!
0%
#702605000000
1!
1%
#702610000000
0!
0%
#702615000000
1!
1%
#702620000000
0!
0%
#702625000000
1!
1%
#702630000000
0!
0%
#702635000000
1!
1%
#702640000000
0!
0%
#702645000000
1!
1%
#702650000000
0!
0%
#702655000000
1!
1%
#702660000000
0!
0%
#702665000000
1!
1%
#702670000000
0!
0%
#702675000000
1!
1%
#702680000000
0!
0%
#702685000000
1!
1%
#702690000000
0!
0%
#702695000000
1!
1%
#702700000000
0!
0%
#702705000000
1!
1%
#702710000000
0!
0%
#702715000000
1!
1%
#702720000000
0!
0%
#702725000000
1!
1%
#702730000000
0!
0%
#702735000000
1!
1%
#702740000000
0!
0%
#702745000000
1!
1%
#702750000000
0!
0%
#702755000000
1!
1%
#702760000000
0!
0%
#702765000000
1!
1%
#702770000000
0!
0%
#702775000000
1!
1%
#702780000000
0!
0%
#702785000000
1!
1%
#702790000000
0!
0%
#702795000000
1!
1%
#702800000000
0!
0%
#702805000000
1!
1%
#702810000000
0!
0%
#702815000000
1!
1%
#702820000000
0!
0%
#702825000000
1!
1%
#702830000000
0!
0%
#702835000000
1!
1%
#702840000000
0!
0%
#702845000000
1!
1%
#702850000000
0!
0%
#702855000000
1!
1%
#702860000000
0!
0%
#702865000000
1!
1%
#702870000000
0!
0%
#702875000000
1!
1%
#702880000000
0!
0%
#702885000000
1!
1%
#702890000000
0!
0%
#702895000000
1!
1%
#702900000000
0!
0%
#702905000000
1!
1%
#702910000000
0!
0%
#702915000000
1!
1%
#702920000000
0!
0%
#702925000000
1!
1%
#702930000000
0!
0%
#702935000000
1!
1%
#702940000000
0!
0%
#702945000000
1!
1%
#702950000000
0!
0%
#702955000000
1!
1%
#702960000000
0!
0%
#702965000000
1!
1%
#702970000000
0!
0%
#702975000000
1!
1%
#702980000000
0!
0%
#702985000000
1!
1%
#702990000000
0!
0%
#702995000000
1!
1%
#703000000000
0!
0%
#703005000000
1!
1%
#703010000000
0!
0%
#703015000000
1!
1%
#703020000000
0!
0%
#703025000000
1!
1%
#703030000000
0!
0%
#703035000000
1!
1%
#703040000000
0!
0%
#703045000000
1!
1%
#703050000000
0!
0%
#703055000000
1!
1%
#703060000000
0!
0%
#703065000000
1!
1%
#703070000000
0!
0%
#703075000000
1!
1%
#703080000000
0!
0%
#703085000000
1!
1%
#703090000000
0!
0%
#703095000000
1!
1%
#703100000000
0!
0%
#703105000000
1!
1%
#703110000000
0!
0%
#703115000000
1!
1%
#703120000000
0!
0%
#703125000000
1!
1%
#703130000000
0!
0%
#703135000000
1!
1%
#703140000000
0!
0%
#703145000000
1!
1%
#703150000000
0!
0%
#703155000000
1!
1%
#703160000000
0!
0%
#703165000000
1!
1%
#703170000000
0!
0%
#703175000000
1!
1%
#703180000000
0!
0%
#703185000000
1!
1%
#703190000000
0!
0%
#703195000000
1!
1%
#703200000000
0!
0%
#703205000000
1!
1%
#703210000000
0!
0%
#703215000000
1!
1%
#703220000000
0!
0%
#703225000000
1!
1%
#703230000000
0!
0%
#703235000000
1!
1%
#703240000000
0!
0%
#703245000000
1!
1%
#703250000000
0!
0%
#703255000000
1!
1%
#703260000000
0!
0%
#703265000000
1!
1%
#703270000000
0!
0%
#703275000000
1!
1%
#703280000000
0!
0%
#703285000000
1!
1%
#703290000000
0!
0%
#703295000000
1!
1%
#703300000000
0!
0%
#703305000000
1!
1%
#703310000000
0!
0%
#703315000000
1!
1%
#703320000000
0!
0%
#703325000000
1!
1%
#703330000000
0!
0%
#703335000000
1!
1%
#703340000000
0!
0%
#703345000000
1!
1%
#703350000000
0!
0%
#703355000000
1!
1%
#703360000000
0!
0%
#703365000000
1!
1%
#703370000000
0!
0%
#703375000000
1!
1%
#703380000000
0!
0%
#703385000000
1!
1%
#703390000000
0!
0%
#703395000000
1!
1%
#703400000000
0!
0%
#703405000000
1!
1%
#703410000000
0!
0%
#703415000000
1!
1%
#703420000000
0!
0%
#703425000000
1!
1%
#703430000000
0!
0%
#703435000000
1!
1%
#703440000000
0!
0%
#703445000000
1!
1%
#703450000000
0!
0%
#703455000000
1!
1%
#703460000000
0!
0%
#703465000000
1!
1%
#703470000000
0!
0%
#703475000000
1!
1%
#703480000000
0!
0%
#703485000000
1!
1%
#703490000000
0!
0%
#703495000000
1!
1%
#703500000000
0!
0%
#703505000000
1!
1%
#703510000000
0!
0%
#703515000000
1!
1%
#703520000000
0!
0%
#703525000000
1!
1%
#703530000000
0!
0%
#703535000000
1!
1%
#703540000000
0!
0%
#703545000000
1!
1%
#703550000000
0!
0%
#703555000000
1!
1%
#703560000000
0!
0%
#703565000000
1!
1%
#703570000000
0!
0%
#703575000000
1!
1%
#703580000000
0!
0%
#703585000000
1!
1%
#703590000000
0!
0%
#703595000000
1!
1%
#703600000000
0!
0%
#703605000000
1!
1%
#703610000000
0!
0%
#703615000000
1!
1%
#703620000000
0!
0%
#703625000000
1!
1%
#703630000000
0!
0%
#703635000000
1!
1%
#703640000000
0!
0%
#703645000000
1!
1%
#703650000000
0!
0%
#703655000000
1!
1%
#703660000000
0!
0%
#703665000000
1!
1%
#703670000000
0!
0%
#703675000000
1!
1%
#703680000000
0!
0%
#703685000000
1!
1%
#703690000000
0!
0%
#703695000000
1!
1%
#703700000000
0!
0%
#703705000000
1!
1%
#703710000000
0!
0%
#703715000000
1!
1%
#703720000000
0!
0%
#703725000000
1!
1%
#703730000000
0!
0%
#703735000000
1!
1%
#703740000000
0!
0%
#703745000000
1!
1%
#703750000000
0!
0%
#703755000000
1!
1%
#703760000000
0!
0%
#703765000000
1!
1%
#703770000000
0!
0%
#703775000000
1!
1%
#703780000000
0!
0%
#703785000000
1!
1%
#703790000000
0!
0%
#703795000000
1!
1%
#703800000000
0!
0%
#703805000000
1!
1%
#703810000000
0!
0%
#703815000000
1!
1%
#703820000000
0!
0%
#703825000000
1!
1%
#703830000000
0!
0%
#703835000000
1!
1%
#703840000000
0!
0%
#703845000000
1!
1%
#703850000000
0!
0%
#703855000000
1!
1%
#703860000000
0!
0%
#703865000000
1!
1%
#703870000000
0!
0%
#703875000000
1!
1%
#703880000000
0!
0%
#703885000000
1!
1%
#703890000000
0!
0%
#703895000000
1!
1%
#703900000000
0!
0%
#703905000000
1!
1%
#703910000000
0!
0%
#703915000000
1!
1%
#703920000000
0!
0%
#703925000000
1!
1%
#703930000000
0!
0%
#703935000000
1!
1%
#703940000000
0!
0%
#703945000000
1!
1%
#703950000000
0!
0%
#703955000000
1!
1%
#703960000000
0!
0%
#703965000000
1!
1%
#703970000000
0!
0%
#703975000000
1!
1%
#703980000000
0!
0%
#703985000000
1!
1%
#703990000000
0!
0%
#703995000000
1!
1%
#704000000000
0!
0%
#704005000000
1!
1%
#704010000000
0!
0%
#704015000000
1!
1%
#704020000000
0!
0%
#704025000000
1!
1%
#704030000000
0!
0%
#704035000000
1!
1%
#704040000000
0!
0%
#704045000000
1!
1%
#704050000000
0!
0%
#704055000000
1!
1%
#704060000000
0!
0%
#704065000000
1!
1%
#704070000000
0!
0%
#704075000000
1!
1%
#704080000000
0!
0%
#704085000000
1!
1%
#704090000000
0!
0%
#704095000000
1!
1%
#704100000000
0!
0%
#704105000000
1!
1%
#704110000000
0!
0%
#704115000000
1!
1%
#704120000000
0!
0%
#704125000000
1!
1%
#704130000000
0!
0%
#704135000000
1!
1%
#704140000000
0!
0%
#704145000000
1!
1%
#704150000000
0!
0%
#704155000000
1!
1%
#704160000000
0!
0%
#704165000000
1!
1%
#704170000000
0!
0%
#704175000000
1!
1%
#704180000000
0!
0%
#704185000000
1!
1%
#704190000000
0!
0%
#704195000000
1!
1%
#704200000000
0!
0%
#704205000000
1!
1%
#704210000000
0!
0%
#704215000000
1!
1%
#704220000000
0!
0%
#704225000000
1!
1%
#704230000000
0!
0%
#704235000000
1!
1%
#704240000000
0!
0%
#704245000000
1!
1%
#704250000000
0!
0%
#704255000000
1!
1%
#704260000000
0!
0%
#704265000000
1!
1%
#704270000000
0!
0%
#704275000000
1!
1%
#704280000000
0!
0%
#704285000000
1!
1%
#704290000000
0!
0%
#704295000000
1!
1%
#704300000000
0!
0%
#704305000000
1!
1%
#704310000000
0!
0%
#704315000000
1!
1%
#704320000000
0!
0%
#704325000000
1!
1%
#704330000000
0!
0%
#704335000000
1!
1%
#704340000000
0!
0%
#704345000000
1!
1%
#704350000000
0!
0%
#704355000000
1!
1%
#704360000000
0!
0%
#704365000000
1!
1%
#704370000000
0!
0%
#704375000000
1!
1%
#704380000000
0!
0%
#704385000000
1!
1%
#704390000000
0!
0%
#704395000000
1!
1%
#704400000000
0!
0%
#704405000000
1!
1%
#704410000000
0!
0%
#704415000000
1!
1%
#704420000000
0!
0%
#704425000000
1!
1%
#704430000000
0!
0%
#704435000000
1!
1%
#704440000000
0!
0%
#704445000000
1!
1%
#704450000000
0!
0%
#704455000000
1!
1%
#704460000000
0!
0%
#704465000000
1!
1%
#704470000000
0!
0%
#704475000000
1!
1%
#704480000000
0!
0%
#704485000000
1!
1%
#704490000000
0!
0%
#704495000000
1!
1%
#704500000000
0!
0%
#704505000000
1!
1%
#704510000000
0!
0%
#704515000000
1!
1%
#704520000000
0!
0%
#704525000000
1!
1%
#704530000000
0!
0%
#704535000000
1!
1%
#704540000000
0!
0%
#704545000000
1!
1%
#704550000000
0!
0%
#704555000000
1!
1%
#704560000000
0!
0%
#704565000000
1!
1%
#704570000000
0!
0%
#704575000000
1!
1%
#704580000000
0!
0%
#704585000000
1!
1%
#704590000000
0!
0%
#704595000000
1!
1%
#704600000000
0!
0%
#704605000000
1!
1%
#704610000000
0!
0%
#704615000000
1!
1%
#704620000000
0!
0%
#704625000000
1!
1%
#704630000000
0!
0%
#704635000000
1!
1%
#704640000000
0!
0%
#704645000000
1!
1%
#704650000000
0!
0%
#704655000000
1!
1%
#704660000000
0!
0%
#704665000000
1!
1%
#704670000000
0!
0%
#704675000000
1!
1%
#704680000000
0!
0%
#704685000000
1!
1%
#704690000000
0!
0%
#704695000000
1!
1%
#704700000000
0!
0%
#704705000000
1!
1%
#704710000000
0!
0%
#704715000000
1!
1%
#704720000000
0!
0%
#704725000000
1!
1%
#704730000000
0!
0%
#704735000000
1!
1%
#704740000000
0!
0%
#704745000000
1!
1%
#704750000000
0!
0%
#704755000000
1!
1%
#704760000000
0!
0%
#704765000000
1!
1%
#704770000000
0!
0%
#704775000000
1!
1%
#704780000000
0!
0%
#704785000000
1!
1%
#704790000000
0!
0%
#704795000000
1!
1%
#704800000000
0!
0%
#704805000000
1!
1%
#704810000000
0!
0%
#704815000000
1!
1%
#704820000000
0!
0%
#704825000000
1!
1%
#704830000000
0!
0%
#704835000000
1!
1%
#704840000000
0!
0%
#704845000000
1!
1%
#704850000000
0!
0%
#704855000000
1!
1%
#704860000000
0!
0%
#704865000000
1!
1%
#704870000000
0!
0%
#704875000000
1!
1%
#704880000000
0!
0%
#704885000000
1!
1%
#704890000000
0!
0%
#704895000000
1!
1%
#704900000000
0!
0%
#704905000000
1!
1%
#704910000000
0!
0%
#704915000000
1!
1%
#704920000000
0!
0%
#704925000000
1!
1%
#704930000000
0!
0%
#704935000000
1!
1%
#704940000000
0!
0%
#704945000000
1!
1%
#704950000000
0!
0%
#704955000000
1!
1%
#704960000000
0!
0%
#704965000000
1!
1%
#704970000000
0!
0%
#704975000000
1!
1%
#704980000000
0!
0%
#704985000000
1!
1%
#704990000000
0!
0%
#704995000000
1!
1%
#705000000000
0!
0%
#705005000000
1!
1%
#705010000000
0!
0%
#705015000000
1!
1%
#705020000000
0!
0%
#705025000000
1!
1%
#705030000000
0!
0%
#705035000000
1!
1%
#705040000000
0!
0%
#705045000000
1!
1%
#705050000000
0!
0%
#705055000000
1!
1%
#705060000000
0!
0%
#705065000000
1!
1%
#705070000000
0!
0%
#705075000000
1!
1%
#705080000000
0!
0%
#705085000000
1!
1%
#705090000000
0!
0%
#705095000000
1!
1%
#705100000000
0!
0%
#705105000000
1!
1%
#705110000000
0!
0%
#705115000000
1!
1%
#705120000000
0!
0%
#705125000000
1!
1%
#705130000000
0!
0%
#705135000000
1!
1%
#705140000000
0!
0%
#705145000000
1!
1%
#705150000000
0!
0%
#705155000000
1!
1%
#705160000000
0!
0%
#705165000000
1!
1%
#705170000000
0!
0%
#705175000000
1!
1%
#705180000000
0!
0%
#705185000000
1!
1%
#705190000000
0!
0%
#705195000000
1!
1%
#705200000000
0!
0%
#705205000000
1!
1%
#705210000000
0!
0%
#705215000000
1!
1%
#705220000000
0!
0%
#705225000000
1!
1%
#705230000000
0!
0%
#705235000000
1!
1%
#705240000000
0!
0%
#705245000000
1!
1%
#705250000000
0!
0%
#705255000000
1!
1%
#705260000000
0!
0%
#705265000000
1!
1%
#705270000000
0!
0%
#705275000000
1!
1%
#705280000000
0!
0%
#705285000000
1!
1%
#705290000000
0!
0%
#705295000000
1!
1%
#705300000000
0!
0%
#705305000000
1!
1%
#705310000000
0!
0%
#705315000000
1!
1%
#705320000000
0!
0%
#705325000000
1!
1%
#705330000000
0!
0%
#705335000000
1!
1%
#705340000000
0!
0%
#705345000000
1!
1%
#705350000000
0!
0%
#705355000000
1!
1%
#705360000000
0!
0%
#705365000000
1!
1%
#705370000000
0!
0%
#705375000000
1!
1%
#705380000000
0!
0%
#705385000000
1!
1%
#705390000000
0!
0%
#705395000000
1!
1%
#705400000000
0!
0%
#705405000000
1!
1%
#705410000000
0!
0%
#705415000000
1!
1%
#705420000000
0!
0%
#705425000000
1!
1%
#705430000000
0!
0%
#705435000000
1!
1%
#705440000000
0!
0%
#705445000000
1!
1%
#705450000000
0!
0%
#705455000000
1!
1%
#705460000000
0!
0%
#705465000000
1!
1%
#705470000000
0!
0%
#705475000000
1!
1%
#705480000000
0!
0%
#705485000000
1!
1%
#705490000000
0!
0%
#705495000000
1!
1%
#705500000000
0!
0%
#705505000000
1!
1%
#705510000000
0!
0%
#705515000000
1!
1%
#705520000000
0!
0%
#705525000000
1!
1%
#705530000000
0!
0%
#705535000000
1!
1%
#705540000000
0!
0%
#705545000000
1!
1%
#705550000000
0!
0%
#705555000000
1!
1%
#705560000000
0!
0%
#705565000000
1!
1%
#705570000000
0!
0%
#705575000000
1!
1%
#705580000000
0!
0%
#705585000000
1!
1%
#705590000000
0!
0%
#705595000000
1!
1%
#705600000000
0!
0%
#705605000000
1!
1%
#705610000000
0!
0%
#705615000000
1!
1%
#705620000000
0!
0%
#705625000000
1!
1%
#705630000000
0!
0%
#705635000000
1!
1%
#705640000000
0!
0%
#705645000000
1!
1%
#705650000000
0!
0%
#705655000000
1!
1%
#705660000000
0!
0%
#705665000000
1!
1%
#705670000000
0!
0%
#705675000000
1!
1%
#705680000000
0!
0%
#705685000000
1!
1%
#705690000000
0!
0%
#705695000000
1!
1%
#705700000000
0!
0%
#705705000000
1!
1%
#705710000000
0!
0%
#705715000000
1!
1%
#705720000000
0!
0%
#705725000000
1!
1%
#705730000000
0!
0%
#705735000000
1!
1%
#705740000000
0!
0%
#705745000000
1!
1%
#705750000000
0!
0%
#705755000000
1!
1%
#705760000000
0!
0%
#705765000000
1!
1%
#705770000000
0!
0%
#705775000000
1!
1%
#705780000000
0!
0%
#705785000000
1!
1%
#705790000000
0!
0%
#705795000000
1!
1%
#705800000000
0!
0%
#705805000000
1!
1%
#705810000000
0!
0%
#705815000000
1!
1%
#705820000000
0!
0%
#705825000000
1!
1%
#705830000000
0!
0%
#705835000000
1!
1%
#705840000000
0!
0%
#705845000000
1!
1%
#705850000000
0!
0%
#705855000000
1!
1%
#705860000000
0!
0%
#705865000000
1!
1%
#705870000000
0!
0%
#705875000000
1!
1%
#705880000000
0!
0%
#705885000000
1!
1%
#705890000000
0!
0%
#705895000000
1!
1%
#705900000000
0!
0%
#705905000000
1!
1%
#705910000000
0!
0%
#705915000000
1!
1%
#705920000000
0!
0%
#705925000000
1!
1%
#705930000000
0!
0%
#705935000000
1!
1%
#705940000000
0!
0%
#705945000000
1!
1%
#705950000000
0!
0%
#705955000000
1!
1%
#705960000000
0!
0%
#705965000000
1!
1%
#705970000000
0!
0%
#705975000000
1!
1%
#705980000000
0!
0%
#705985000000
1!
1%
#705990000000
0!
0%
#705995000000
1!
1%
#706000000000
0!
0%
#706005000000
1!
1%
#706010000000
0!
0%
#706015000000
1!
1%
#706020000000
0!
0%
#706025000000
1!
1%
#706030000000
0!
0%
#706035000000
1!
1%
#706040000000
0!
0%
#706045000000
1!
1%
#706050000000
0!
0%
#706055000000
1!
1%
#706060000000
0!
0%
#706065000000
1!
1%
#706070000000
0!
0%
#706075000000
1!
1%
#706080000000
0!
0%
#706085000000
1!
1%
#706090000000
0!
0%
#706095000000
1!
1%
#706100000000
0!
0%
#706105000000
1!
1%
#706110000000
0!
0%
#706115000000
1!
1%
#706120000000
0!
0%
#706125000000
1!
1%
#706130000000
0!
0%
#706135000000
1!
1%
#706140000000
0!
0%
#706145000000
1!
1%
#706150000000
0!
0%
#706155000000
1!
1%
#706160000000
0!
0%
#706165000000
1!
1%
#706170000000
0!
0%
#706175000000
1!
1%
#706180000000
0!
0%
#706185000000
1!
1%
#706190000000
0!
0%
#706195000000
1!
1%
#706200000000
0!
0%
#706205000000
1!
1%
#706210000000
0!
0%
#706215000000
1!
1%
#706220000000
0!
0%
#706225000000
1!
1%
#706230000000
0!
0%
#706235000000
1!
1%
#706240000000
0!
0%
#706245000000
1!
1%
#706250000000
0!
0%
#706255000000
1!
1%
#706260000000
0!
0%
#706265000000
1!
1%
#706270000000
0!
0%
#706275000000
1!
1%
#706280000000
0!
0%
#706285000000
1!
1%
#706290000000
0!
0%
#706295000000
1!
1%
#706300000000
0!
0%
#706305000000
1!
1%
#706310000000
0!
0%
#706315000000
1!
1%
#706320000000
0!
0%
#706325000000
1!
1%
#706330000000
0!
0%
#706335000000
1!
1%
#706340000000
0!
0%
#706345000000
1!
1%
#706350000000
0!
0%
#706355000000
1!
1%
#706360000000
0!
0%
#706365000000
1!
1%
#706370000000
0!
0%
#706375000000
1!
1%
#706380000000
0!
0%
#706385000000
1!
1%
#706390000000
0!
0%
#706395000000
1!
1%
#706400000000
0!
0%
#706405000000
1!
1%
#706410000000
0!
0%
#706415000000
1!
1%
#706420000000
0!
0%
#706425000000
1!
1%
#706430000000
0!
0%
#706435000000
1!
1%
#706440000000
0!
0%
#706445000000
1!
1%
#706450000000
0!
0%
#706455000000
1!
1%
#706460000000
0!
0%
#706465000000
1!
1%
#706470000000
0!
0%
#706475000000
1!
1%
#706480000000
0!
0%
#706485000000
1!
1%
#706490000000
0!
0%
#706495000000
1!
1%
#706500000000
0!
0%
#706505000000
1!
1%
#706510000000
0!
0%
#706515000000
1!
1%
#706520000000
0!
0%
#706525000000
1!
1%
#706530000000
0!
0%
#706535000000
1!
1%
#706540000000
0!
0%
#706545000000
1!
1%
#706550000000
0!
0%
#706555000000
1!
1%
#706560000000
0!
0%
#706565000000
1!
1%
#706570000000
0!
0%
#706575000000
1!
1%
#706580000000
0!
0%
#706585000000
1!
1%
#706590000000
0!
0%
#706595000000
1!
1%
#706600000000
0!
0%
#706605000000
1!
1%
#706610000000
0!
0%
#706615000000
1!
1%
#706620000000
0!
0%
#706625000000
1!
1%
#706630000000
0!
0%
#706635000000
1!
1%
#706640000000
0!
0%
#706645000000
1!
1%
#706650000000
0!
0%
#706655000000
1!
1%
#706660000000
0!
0%
#706665000000
1!
1%
#706670000000
0!
0%
#706675000000
1!
1%
#706680000000
0!
0%
#706685000000
1!
1%
#706690000000
0!
0%
#706695000000
1!
1%
#706700000000
0!
0%
#706705000000
1!
1%
#706710000000
0!
0%
#706715000000
1!
1%
#706720000000
0!
0%
#706725000000
1!
1%
#706730000000
0!
0%
#706735000000
1!
1%
#706740000000
0!
0%
#706745000000
1!
1%
#706750000000
0!
0%
#706755000000
1!
1%
#706760000000
0!
0%
#706765000000
1!
1%
#706770000000
0!
0%
#706775000000
1!
1%
#706780000000
0!
0%
#706785000000
1!
1%
#706790000000
0!
0%
#706795000000
1!
1%
#706800000000
0!
0%
#706805000000
1!
1%
#706810000000
0!
0%
#706815000000
1!
1%
#706820000000
0!
0%
#706825000000
1!
1%
#706830000000
0!
0%
#706835000000
1!
1%
#706840000000
0!
0%
#706845000000
1!
1%
#706850000000
0!
0%
#706855000000
1!
1%
#706860000000
0!
0%
#706865000000
1!
1%
#706870000000
0!
0%
#706875000000
1!
1%
#706880000000
0!
0%
#706885000000
1!
1%
#706890000000
0!
0%
#706895000000
1!
1%
#706900000000
0!
0%
#706905000000
1!
1%
#706910000000
0!
0%
#706915000000
1!
1%
#706920000000
0!
0%
#706925000000
1!
1%
#706930000000
0!
0%
#706935000000
1!
1%
#706940000000
0!
0%
#706945000000
1!
1%
#706950000000
0!
0%
#706955000000
1!
1%
#706960000000
0!
0%
#706965000000
1!
1%
#706970000000
0!
0%
#706975000000
1!
1%
#706980000000
0!
0%
#706985000000
1!
1%
#706990000000
0!
0%
#706995000000
1!
1%
#707000000000
0!
0%
#707005000000
1!
1%
#707010000000
0!
0%
#707015000000
1!
1%
#707020000000
0!
0%
#707025000000
1!
1%
#707030000000
0!
0%
#707035000000
1!
1%
#707040000000
0!
0%
#707045000000
1!
1%
#707050000000
0!
0%
#707055000000
1!
1%
#707060000000
0!
0%
#707065000000
1!
1%
#707070000000
0!
0%
#707075000000
1!
1%
#707080000000
0!
0%
#707085000000
1!
1%
#707090000000
0!
0%
#707095000000
1!
1%
#707100000000
0!
0%
#707105000000
1!
1%
#707110000000
0!
0%
#707115000000
1!
1%
#707120000000
0!
0%
#707125000000
1!
1%
#707130000000
0!
0%
#707135000000
1!
1%
#707140000000
0!
0%
#707145000000
1!
1%
#707150000000
0!
0%
#707155000000
1!
1%
#707160000000
0!
0%
#707165000000
1!
1%
#707170000000
0!
0%
#707175000000
1!
1%
#707180000000
0!
0%
#707185000000
1!
1%
#707190000000
0!
0%
#707195000000
1!
1%
#707200000000
0!
0%
#707205000000
1!
1%
#707210000000
0!
0%
#707215000000
1!
1%
#707220000000
0!
0%
#707225000000
1!
1%
#707230000000
0!
0%
#707235000000
1!
1%
#707240000000
0!
0%
#707245000000
1!
1%
#707250000000
0!
0%
#707255000000
1!
1%
#707260000000
0!
0%
#707265000000
1!
1%
#707270000000
0!
0%
#707275000000
1!
1%
#707280000000
0!
0%
#707285000000
1!
1%
#707290000000
0!
0%
#707295000000
1!
1%
#707300000000
0!
0%
#707305000000
1!
1%
#707310000000
0!
0%
#707315000000
1!
1%
#707320000000
0!
0%
#707325000000
1!
1%
#707330000000
0!
0%
#707335000000
1!
1%
#707340000000
0!
0%
#707345000000
1!
1%
#707350000000
0!
0%
#707355000000
1!
1%
#707360000000
0!
0%
#707365000000
1!
1%
#707370000000
0!
0%
#707375000000
1!
1%
#707380000000
0!
0%
#707385000000
1!
1%
#707390000000
0!
0%
#707395000000
1!
1%
#707400000000
0!
0%
#707405000000
1!
1%
#707410000000
0!
0%
#707415000000
1!
1%
#707420000000
0!
0%
#707425000000
1!
1%
#707430000000
0!
0%
#707435000000
1!
1%
#707440000000
0!
0%
#707445000000
1!
1%
#707450000000
0!
0%
#707455000000
1!
1%
#707460000000
0!
0%
#707465000000
1!
1%
#707470000000
0!
0%
#707475000000
1!
1%
#707480000000
0!
0%
#707485000000
1!
1%
#707490000000
0!
0%
#707495000000
1!
1%
#707500000000
0!
0%
#707505000000
1!
1%
#707510000000
0!
0%
#707515000000
1!
1%
#707520000000
0!
0%
#707525000000
1!
1%
#707530000000
0!
0%
#707535000000
1!
1%
#707540000000
0!
0%
#707545000000
1!
1%
#707550000000
0!
0%
#707555000000
1!
1%
#707560000000
0!
0%
#707565000000
1!
1%
#707570000000
0!
0%
#707575000000
1!
1%
#707580000000
0!
0%
#707585000000
1!
1%
#707590000000
0!
0%
#707595000000
1!
1%
#707600000000
0!
0%
#707605000000
1!
1%
#707610000000
0!
0%
#707615000000
1!
1%
#707620000000
0!
0%
#707625000000
1!
1%
#707630000000
0!
0%
#707635000000
1!
1%
#707640000000
0!
0%
#707645000000
1!
1%
#707650000000
0!
0%
#707655000000
1!
1%
#707660000000
0!
0%
#707665000000
1!
1%
#707670000000
0!
0%
#707675000000
1!
1%
#707680000000
0!
0%
#707685000000
1!
1%
#707690000000
0!
0%
#707695000000
1!
1%
#707700000000
0!
0%
#707705000000
1!
1%
#707710000000
0!
0%
#707715000000
1!
1%
#707720000000
0!
0%
#707725000000
1!
1%
#707730000000
0!
0%
#707735000000
1!
1%
#707740000000
0!
0%
#707745000000
1!
1%
#707750000000
0!
0%
#707755000000
1!
1%
#707760000000
0!
0%
#707765000000
1!
1%
#707770000000
0!
0%
#707775000000
1!
1%
#707780000000
0!
0%
#707785000000
1!
1%
#707790000000
0!
0%
#707795000000
1!
1%
#707800000000
0!
0%
#707805000000
1!
1%
#707810000000
0!
0%
#707815000000
1!
1%
#707820000000
0!
0%
#707825000000
1!
1%
#707830000000
0!
0%
#707835000000
1!
1%
#707840000000
0!
0%
#707845000000
1!
1%
#707850000000
0!
0%
#707855000000
1!
1%
#707860000000
0!
0%
#707865000000
1!
1%
#707870000000
0!
0%
#707875000000
1!
1%
#707880000000
0!
0%
#707885000000
1!
1%
#707890000000
0!
0%
#707895000000
1!
1%
#707900000000
0!
0%
#707905000000
1!
1%
#707910000000
0!
0%
#707915000000
1!
1%
#707920000000
0!
0%
#707925000000
1!
1%
#707930000000
0!
0%
#707935000000
1!
1%
#707940000000
0!
0%
#707945000000
1!
1%
#707950000000
0!
0%
#707955000000
1!
1%
#707960000000
0!
0%
#707965000000
1!
1%
#707970000000
0!
0%
#707975000000
1!
1%
#707980000000
0!
0%
#707985000000
1!
1%
#707990000000
0!
0%
#707995000000
1!
1%
#708000000000
0!
0%
#708005000000
1!
1%
#708010000000
0!
0%
#708015000000
1!
1%
#708020000000
0!
0%
#708025000000
1!
1%
#708030000000
0!
0%
#708035000000
1!
1%
#708040000000
0!
0%
#708045000000
1!
1%
#708050000000
0!
0%
#708055000000
1!
1%
#708060000000
0!
0%
#708065000000
1!
1%
#708070000000
0!
0%
#708075000000
1!
1%
#708080000000
0!
0%
#708085000000
1!
1%
#708090000000
0!
0%
#708095000000
1!
1%
#708100000000
0!
0%
#708105000000
1!
1%
#708110000000
0!
0%
#708115000000
1!
1%
#708120000000
0!
0%
#708125000000
1!
1%
#708130000000
0!
0%
#708135000000
1!
1%
#708140000000
0!
0%
#708145000000
1!
1%
#708150000000
0!
0%
#708155000000
1!
1%
#708160000000
0!
0%
#708165000000
1!
1%
#708170000000
0!
0%
#708175000000
1!
1%
#708180000000
0!
0%
#708185000000
1!
1%
#708190000000
0!
0%
#708195000000
1!
1%
#708200000000
0!
0%
#708205000000
1!
1%
#708210000000
0!
0%
#708215000000
1!
1%
#708220000000
0!
0%
#708225000000
1!
1%
#708230000000
0!
0%
#708235000000
1!
1%
#708240000000
0!
0%
#708245000000
1!
1%
#708250000000
0!
0%
#708255000000
1!
1%
#708260000000
0!
0%
#708265000000
1!
1%
#708270000000
0!
0%
#708275000000
1!
1%
#708280000000
0!
0%
#708285000000
1!
1%
#708290000000
0!
0%
#708295000000
1!
1%
#708300000000
0!
0%
#708305000000
1!
1%
#708310000000
0!
0%
#708315000000
1!
1%
#708320000000
0!
0%
#708325000000
1!
1%
#708330000000
0!
0%
#708335000000
1!
1%
#708340000000
0!
0%
#708345000000
1!
1%
#708350000000
0!
0%
#708355000000
1!
1%
#708360000000
0!
0%
#708365000000
1!
1%
#708370000000
0!
0%
#708375000000
1!
1%
#708380000000
0!
0%
#708385000000
1!
1%
#708390000000
0!
0%
#708395000000
1!
1%
#708400000000
0!
0%
#708405000000
1!
1%
#708410000000
0!
0%
#708415000000
1!
1%
#708420000000
0!
0%
#708425000000
1!
1%
#708430000000
0!
0%
#708435000000
1!
1%
#708440000000
0!
0%
#708445000000
1!
1%
#708450000000
0!
0%
#708455000000
1!
1%
#708460000000
0!
0%
#708465000000
1!
1%
#708470000000
0!
0%
#708475000000
1!
1%
#708480000000
0!
0%
#708485000000
1!
1%
#708490000000
0!
0%
#708495000000
1!
1%
#708500000000
0!
0%
#708505000000
1!
1%
#708510000000
0!
0%
#708515000000
1!
1%
#708520000000
0!
0%
#708525000000
1!
1%
#708530000000
0!
0%
#708535000000
1!
1%
#708540000000
0!
0%
#708545000000
1!
1%
#708550000000
0!
0%
#708555000000
1!
1%
#708560000000
0!
0%
#708565000000
1!
1%
#708570000000
0!
0%
#708575000000
1!
1%
#708580000000
0!
0%
#708585000000
1!
1%
#708590000000
0!
0%
#708595000000
1!
1%
#708600000000
0!
0%
#708605000000
1!
1%
#708610000000
0!
0%
#708615000000
1!
1%
#708620000000
0!
0%
#708625000000
1!
1%
#708630000000
0!
0%
#708635000000
1!
1%
#708640000000
0!
0%
#708645000000
1!
1%
#708650000000
0!
0%
#708655000000
1!
1%
#708660000000
0!
0%
#708665000000
1!
1%
#708670000000
0!
0%
#708675000000
1!
1%
#708680000000
0!
0%
#708685000000
1!
1%
#708690000000
0!
0%
#708695000000
1!
1%
#708700000000
0!
0%
#708705000000
1!
1%
#708710000000
0!
0%
#708715000000
1!
1%
#708720000000
0!
0%
#708725000000
1!
1%
#708730000000
0!
0%
#708735000000
1!
1%
#708740000000
0!
0%
#708745000000
1!
1%
#708750000000
0!
0%
#708755000000
1!
1%
#708760000000
0!
0%
#708765000000
1!
1%
#708770000000
0!
0%
#708775000000
1!
1%
#708780000000
0!
0%
#708785000000
1!
1%
#708790000000
0!
0%
#708795000000
1!
1%
#708800000000
0!
0%
#708805000000
1!
1%
#708810000000
0!
0%
#708815000000
1!
1%
#708820000000
0!
0%
#708825000000
1!
1%
#708830000000
0!
0%
#708835000000
1!
1%
#708840000000
0!
0%
#708845000000
1!
1%
#708850000000
0!
0%
#708855000000
1!
1%
#708860000000
0!
0%
#708865000000
1!
1%
#708870000000
0!
0%
#708875000000
1!
1%
#708880000000
0!
0%
#708885000000
1!
1%
#708890000000
0!
0%
#708895000000
1!
1%
#708900000000
0!
0%
#708905000000
1!
1%
#708910000000
0!
0%
#708915000000
1!
1%
#708920000000
0!
0%
#708925000000
1!
1%
#708930000000
0!
0%
#708935000000
1!
1%
#708940000000
0!
0%
#708945000000
1!
1%
#708950000000
0!
0%
#708955000000
1!
1%
#708960000000
0!
0%
#708965000000
1!
1%
#708970000000
0!
0%
#708975000000
1!
1%
#708980000000
0!
0%
#708985000000
1!
1%
#708990000000
0!
0%
#708995000000
1!
1%
#709000000000
0!
0%
#709005000000
1!
1%
#709010000000
0!
0%
#709015000000
1!
1%
#709020000000
0!
0%
#709025000000
1!
1%
#709030000000
0!
0%
#709035000000
1!
1%
#709040000000
0!
0%
#709045000000
1!
1%
#709050000000
0!
0%
#709055000000
1!
1%
#709060000000
0!
0%
#709065000000
1!
1%
#709070000000
0!
0%
#709075000000
1!
1%
#709080000000
0!
0%
#709085000000
1!
1%
#709090000000
0!
0%
#709095000000
1!
1%
#709100000000
0!
0%
#709105000000
1!
1%
#709110000000
0!
0%
#709115000000
1!
1%
#709120000000
0!
0%
#709125000000
1!
1%
#709130000000
0!
0%
#709135000000
1!
1%
#709140000000
0!
0%
#709145000000
1!
1%
#709150000000
0!
0%
#709155000000
1!
1%
#709160000000
0!
0%
#709165000000
1!
1%
#709170000000
0!
0%
#709175000000
1!
1%
#709180000000
0!
0%
#709185000000
1!
1%
#709190000000
0!
0%
#709195000000
1!
1%
#709200000000
0!
0%
#709205000000
1!
1%
#709210000000
0!
0%
#709215000000
1!
1%
#709220000000
0!
0%
#709225000000
1!
1%
#709230000000
0!
0%
#709235000000
1!
1%
#709240000000
0!
0%
#709245000000
1!
1%
#709250000000
0!
0%
#709255000000
1!
1%
#709260000000
0!
0%
#709265000000
1!
1%
#709270000000
0!
0%
#709275000000
1!
1%
#709280000000
0!
0%
#709285000000
1!
1%
#709290000000
0!
0%
#709295000000
1!
1%
#709300000000
0!
0%
#709305000000
1!
1%
#709310000000
0!
0%
#709315000000
1!
1%
#709320000000
0!
0%
#709325000000
1!
1%
#709330000000
0!
0%
#709335000000
1!
1%
#709340000000
0!
0%
#709345000000
1!
1%
#709350000000
0!
0%
#709355000000
1!
1%
#709360000000
0!
0%
#709365000000
1!
1%
#709370000000
0!
0%
#709375000000
1!
1%
#709380000000
0!
0%
#709385000000
1!
1%
#709390000000
0!
0%
#709395000000
1!
1%
#709400000000
0!
0%
#709405000000
1!
1%
#709410000000
0!
0%
#709415000000
1!
1%
#709420000000
0!
0%
#709425000000
1!
1%
#709430000000
0!
0%
#709435000000
1!
1%
#709440000000
0!
0%
#709445000000
1!
1%
#709450000000
0!
0%
#709455000000
1!
1%
#709460000000
0!
0%
#709465000000
1!
1%
#709470000000
0!
0%
#709475000000
1!
1%
#709480000000
0!
0%
#709485000000
1!
1%
#709490000000
0!
0%
#709495000000
1!
1%
#709500000000
0!
0%
#709505000000
1!
1%
#709510000000
0!
0%
#709515000000
1!
1%
#709520000000
0!
0%
#709525000000
1!
1%
#709530000000
0!
0%
#709535000000
1!
1%
#709540000000
0!
0%
#709545000000
1!
1%
#709550000000
0!
0%
#709555000000
1!
1%
#709560000000
0!
0%
#709565000000
1!
1%
#709570000000
0!
0%
#709575000000
1!
1%
#709580000000
0!
0%
#709585000000
1!
1%
#709590000000
0!
0%
#709595000000
1!
1%
#709600000000
0!
0%
#709605000000
1!
1%
#709610000000
0!
0%
#709615000000
1!
1%
#709620000000
0!
0%
#709625000000
1!
1%
#709630000000
0!
0%
#709635000000
1!
1%
#709640000000
0!
0%
#709645000000
1!
1%
#709650000000
0!
0%
#709655000000
1!
1%
#709660000000
0!
0%
#709665000000
1!
1%
#709670000000
0!
0%
#709675000000
1!
1%
#709680000000
0!
0%
#709685000000
1!
1%
#709690000000
0!
0%
#709695000000
1!
1%
#709700000000
0!
0%
#709705000000
1!
1%
#709710000000
0!
0%
#709715000000
1!
1%
#709720000000
0!
0%
#709725000000
1!
1%
#709730000000
0!
0%
#709735000000
1!
1%
#709740000000
0!
0%
#709745000000
1!
1%
#709750000000
0!
0%
#709755000000
1!
1%
#709760000000
0!
0%
#709765000000
1!
1%
#709770000000
0!
0%
#709775000000
1!
1%
#709780000000
0!
0%
#709785000000
1!
1%
#709790000000
0!
0%
#709795000000
1!
1%
#709800000000
0!
0%
#709805000000
1!
1%
#709810000000
0!
0%
#709815000000
1!
1%
#709820000000
0!
0%
#709825000000
1!
1%
#709830000000
0!
0%
#709835000000
1!
1%
#709840000000
0!
0%
#709845000000
1!
1%
#709850000000
0!
0%
#709855000000
1!
1%
#709860000000
0!
0%
#709865000000
1!
1%
#709870000000
0!
0%
#709875000000
1!
1%
#709880000000
0!
0%
#709885000000
1!
1%
#709890000000
0!
0%
#709895000000
1!
1%
#709900000000
0!
0%
#709905000000
1!
1%
#709910000000
0!
0%
#709915000000
1!
1%
#709920000000
0!
0%
#709925000000
1!
1%
#709930000000
0!
0%
#709935000000
1!
1%
#709940000000
0!
0%
#709945000000
1!
1%
#709950000000
0!
0%
#709955000000
1!
1%
#709960000000
0!
0%
#709965000000
1!
1%
#709970000000
0!
0%
#709975000000
1!
1%
#709980000000
0!
0%
#709985000000
1!
1%
#709990000000
0!
0%
#709995000000
1!
1%
#710000000000
0!
0%
#710005000000
1!
1%
#710010000000
0!
0%
#710015000000
1!
1%
#710020000000
0!
0%
#710025000000
1!
1%
#710030000000
0!
0%
#710035000000
1!
1%
#710040000000
0!
0%
#710045000000
1!
1%
#710050000000
0!
0%
#710055000000
1!
1%
#710060000000
0!
0%
#710065000000
1!
1%
#710070000000
0!
0%
#710075000000
1!
1%
#710080000000
0!
0%
#710085000000
1!
1%
#710090000000
0!
0%
#710095000000
1!
1%
#710100000000
0!
0%
#710105000000
1!
1%
#710110000000
0!
0%
#710115000000
1!
1%
#710120000000
0!
0%
#710125000000
1!
1%
#710130000000
0!
0%
#710135000000
1!
1%
#710140000000
0!
0%
#710145000000
1!
1%
#710150000000
0!
0%
#710155000000
1!
1%
#710160000000
0!
0%
#710165000000
1!
1%
#710170000000
0!
0%
#710175000000
1!
1%
#710180000000
0!
0%
#710185000000
1!
1%
#710190000000
0!
0%
#710195000000
1!
1%
#710200000000
0!
0%
#710205000000
1!
1%
#710210000000
0!
0%
#710215000000
1!
1%
#710220000000
0!
0%
#710225000000
1!
1%
#710230000000
0!
0%
#710235000000
1!
1%
#710240000000
0!
0%
#710245000000
1!
1%
#710250000000
0!
0%
#710255000000
1!
1%
#710260000000
0!
0%
#710265000000
1!
1%
#710270000000
0!
0%
#710275000000
1!
1%
#710280000000
0!
0%
#710285000000
1!
1%
#710290000000
0!
0%
#710295000000
1!
1%
#710300000000
0!
0%
#710305000000
1!
1%
#710310000000
0!
0%
#710315000000
1!
1%
#710320000000
0!
0%
#710325000000
1!
1%
#710330000000
0!
0%
#710335000000
1!
1%
#710340000000
0!
0%
#710345000000
1!
1%
#710350000000
0!
0%
#710355000000
1!
1%
#710360000000
0!
0%
#710365000000
1!
1%
#710370000000
0!
0%
#710375000000
1!
1%
#710380000000
0!
0%
#710385000000
1!
1%
#710390000000
0!
0%
#710395000000
1!
1%
#710400000000
0!
0%
#710405000000
1!
1%
#710410000000
0!
0%
#710415000000
1!
1%
#710420000000
0!
0%
#710425000000
1!
1%
#710430000000
0!
0%
#710435000000
1!
1%
#710440000000
0!
0%
#710445000000
1!
1%
#710450000000
0!
0%
#710455000000
1!
1%
#710460000000
0!
0%
#710465000000
1!
1%
#710470000000
0!
0%
#710475000000
1!
1%
#710480000000
0!
0%
#710485000000
1!
1%
#710490000000
0!
0%
#710495000000
1!
1%
#710500000000
0!
0%
#710505000000
1!
1%
#710510000000
0!
0%
#710515000000
1!
1%
#710520000000
0!
0%
#710525000000
1!
1%
#710530000000
0!
0%
#710535000000
1!
1%
#710540000000
0!
0%
#710545000000
1!
1%
#710550000000
0!
0%
#710555000000
1!
1%
#710560000000
0!
0%
#710565000000
1!
1%
#710570000000
0!
0%
#710575000000
1!
1%
#710580000000
0!
0%
#710585000000
1!
1%
#710590000000
0!
0%
#710595000000
1!
1%
#710600000000
0!
0%
#710605000000
1!
1%
#710610000000
0!
0%
#710615000000
1!
1%
#710620000000
0!
0%
#710625000000
1!
1%
#710630000000
0!
0%
#710635000000
1!
1%
#710640000000
0!
0%
#710645000000
1!
1%
#710650000000
0!
0%
#710655000000
1!
1%
#710660000000
0!
0%
#710665000000
1!
1%
#710670000000
0!
0%
#710675000000
1!
1%
#710680000000
0!
0%
#710685000000
1!
1%
#710690000000
0!
0%
#710695000000
1!
1%
#710700000000
0!
0%
#710705000000
1!
1%
#710710000000
0!
0%
#710715000000
1!
1%
#710720000000
0!
0%
#710725000000
1!
1%
#710730000000
0!
0%
#710735000000
1!
1%
#710740000000
0!
0%
#710745000000
1!
1%
#710750000000
0!
0%
#710755000000
1!
1%
#710760000000
0!
0%
#710765000000
1!
1%
#710770000000
0!
0%
#710775000000
1!
1%
#710780000000
0!
0%
#710785000000
1!
1%
#710790000000
0!
0%
#710795000000
1!
1%
#710800000000
0!
0%
#710805000000
1!
1%
#710810000000
0!
0%
#710815000000
1!
1%
#710820000000
0!
0%
#710825000000
1!
1%
#710830000000
0!
0%
#710835000000
1!
1%
#710840000000
0!
0%
#710845000000
1!
1%
#710850000000
0!
0%
#710855000000
1!
1%
#710860000000
0!
0%
#710865000000
1!
1%
#710870000000
0!
0%
#710875000000
1!
1%
#710880000000
0!
0%
#710885000000
1!
1%
#710890000000
0!
0%
#710895000000
1!
1%
#710900000000
0!
0%
#710905000000
1!
1%
#710910000000
0!
0%
#710915000000
1!
1%
#710920000000
0!
0%
#710925000000
1!
1%
#710930000000
0!
0%
#710935000000
1!
1%
#710940000000
0!
0%
#710945000000
1!
1%
#710950000000
0!
0%
#710955000000
1!
1%
#710960000000
0!
0%
#710965000000
1!
1%
#710970000000
0!
0%
#710975000000
1!
1%
#710980000000
0!
0%
#710985000000
1!
1%
#710990000000
0!
0%
#710995000000
1!
1%
#711000000000
0!
0%
#711005000000
1!
1%
#711010000000
0!
0%
#711015000000
1!
1%
#711020000000
0!
0%
#711025000000
1!
1%
#711030000000
0!
0%
#711035000000
1!
1%
#711040000000
0!
0%
#711045000000
1!
1%
#711050000000
0!
0%
#711055000000
1!
1%
#711060000000
0!
0%
#711065000000
1!
1%
#711070000000
0!
0%
#711075000000
1!
1%
#711080000000
0!
0%
#711085000000
1!
1%
#711090000000
0!
0%
#711095000000
1!
1%
#711100000000
0!
0%
#711105000000
1!
1%
#711110000000
0!
0%
#711115000000
1!
1%
#711120000000
0!
0%
#711125000000
1!
1%
#711130000000
0!
0%
#711135000000
1!
1%
#711140000000
0!
0%
#711145000000
1!
1%
#711150000000
0!
0%
#711155000000
1!
1%
#711160000000
0!
0%
#711165000000
1!
1%
#711170000000
0!
0%
#711175000000
1!
1%
#711180000000
0!
0%
#711185000000
1!
1%
#711190000000
0!
0%
#711195000000
1!
1%
#711200000000
0!
0%
#711205000000
1!
1%
#711210000000
0!
0%
#711215000000
1!
1%
#711220000000
0!
0%
#711225000000
1!
1%
#711230000000
0!
0%
#711235000000
1!
1%
#711240000000
0!
0%
#711245000000
1!
1%
#711250000000
0!
0%
#711255000000
1!
1%
#711260000000
0!
0%
#711265000000
1!
1%
#711270000000
0!
0%
#711275000000
1!
1%
#711280000000
0!
0%
#711285000000
1!
1%
#711290000000
0!
0%
#711295000000
1!
1%
#711300000000
0!
0%
#711305000000
1!
1%
#711310000000
0!
0%
#711315000000
1!
1%
#711320000000
0!
0%
#711325000000
1!
1%
#711330000000
0!
0%
#711335000000
1!
1%
#711340000000
0!
0%
#711345000000
1!
1%
#711350000000
0!
0%
#711355000000
1!
1%
#711360000000
0!
0%
#711365000000
1!
1%
#711370000000
0!
0%
#711375000000
1!
1%
#711380000000
0!
0%
#711385000000
1!
1%
#711390000000
0!
0%
#711395000000
1!
1%
#711400000000
0!
0%
#711405000000
1!
1%
#711410000000
0!
0%
#711415000000
1!
1%
#711420000000
0!
0%
#711425000000
1!
1%
#711430000000
0!
0%
#711435000000
1!
1%
#711440000000
0!
0%
#711445000000
1!
1%
#711450000000
0!
0%
#711455000000
1!
1%
#711460000000
0!
0%
#711465000000
1!
1%
#711470000000
0!
0%
#711475000000
1!
1%
#711480000000
0!
0%
#711485000000
1!
1%
#711490000000
0!
0%
#711495000000
1!
1%
#711500000000
0!
0%
#711505000000
1!
1%
#711510000000
0!
0%
#711515000000
1!
1%
#711520000000
0!
0%
#711525000000
1!
1%
#711530000000
0!
0%
#711535000000
1!
1%
#711540000000
0!
0%
#711545000000
1!
1%
#711550000000
0!
0%
#711555000000
1!
1%
#711560000000
0!
0%
#711565000000
1!
1%
#711570000000
0!
0%
#711575000000
1!
1%
#711580000000
0!
0%
#711585000000
1!
1%
#711590000000
0!
0%
#711595000000
1!
1%
#711600000000
0!
0%
#711605000000
1!
1%
#711610000000
0!
0%
#711615000000
1!
1%
#711620000000
0!
0%
#711625000000
1!
1%
#711630000000
0!
0%
#711635000000
1!
1%
#711640000000
0!
0%
#711645000000
1!
1%
#711650000000
0!
0%
#711655000000
1!
1%
#711660000000
0!
0%
#711665000000
1!
1%
#711670000000
0!
0%
#711675000000
1!
1%
#711680000000
0!
0%
#711685000000
1!
1%
#711690000000
0!
0%
#711695000000
1!
1%
#711700000000
0!
0%
#711705000000
1!
1%
#711710000000
0!
0%
#711715000000
1!
1%
#711720000000
0!
0%
#711725000000
1!
1%
#711730000000
0!
0%
#711735000000
1!
1%
#711740000000
0!
0%
#711745000000
1!
1%
#711750000000
0!
0%
#711755000000
1!
1%
#711760000000
0!
0%
#711765000000
1!
1%
#711770000000
0!
0%
#711775000000
1!
1%
#711780000000
0!
0%
#711785000000
1!
1%
#711790000000
0!
0%
#711795000000
1!
1%
#711800000000
0!
0%
#711805000000
1!
1%
#711810000000
0!
0%
#711815000000
1!
1%
#711820000000
0!
0%
#711825000000
1!
1%
#711830000000
0!
0%
#711835000000
1!
1%
#711840000000
0!
0%
#711845000000
1!
1%
#711850000000
0!
0%
#711855000000
1!
1%
#711860000000
0!
0%
#711865000000
1!
1%
#711870000000
0!
0%
#711875000000
1!
1%
#711880000000
0!
0%
#711885000000
1!
1%
#711890000000
0!
0%
#711895000000
1!
1%
#711900000000
0!
0%
#711905000000
1!
1%
#711910000000
0!
0%
#711915000000
1!
1%
#711920000000
0!
0%
#711925000000
1!
1%
#711930000000
0!
0%
#711935000000
1!
1%
#711940000000
0!
0%
#711945000000
1!
1%
#711950000000
0!
0%
#711955000000
1!
1%
#711960000000
0!
0%
#711965000000
1!
1%
#711970000000
0!
0%
#711975000000
1!
1%
#711980000000
0!
0%
#711985000000
1!
1%
#711990000000
0!
0%
#711995000000
1!
1%
#712000000000
0!
0%
#712005000000
1!
1%
#712010000000
0!
0%
#712015000000
1!
1%
#712020000000
0!
0%
#712025000000
1!
1%
#712030000000
0!
0%
#712035000000
1!
1%
#712040000000
0!
0%
#712045000000
1!
1%
#712050000000
0!
0%
#712055000000
1!
1%
#712060000000
0!
0%
#712065000000
1!
1%
#712070000000
0!
0%
#712075000000
1!
1%
#712080000000
0!
0%
#712085000000
1!
1%
#712090000000
0!
0%
#712095000000
1!
1%
#712100000000
0!
0%
#712105000000
1!
1%
#712110000000
0!
0%
#712115000000
1!
1%
#712120000000
0!
0%
#712125000000
1!
1%
#712130000000
0!
0%
#712135000000
1!
1%
#712140000000
0!
0%
#712145000000
1!
1%
#712150000000
0!
0%
#712155000000
1!
1%
#712160000000
0!
0%
#712165000000
1!
1%
#712170000000
0!
0%
#712175000000
1!
1%
#712180000000
0!
0%
#712185000000
1!
1%
#712190000000
0!
0%
#712195000000
1!
1%
#712200000000
0!
0%
#712205000000
1!
1%
#712210000000
0!
0%
#712215000000
1!
1%
#712220000000
0!
0%
#712225000000
1!
1%
#712230000000
0!
0%
#712235000000
1!
1%
#712240000000
0!
0%
#712245000000
1!
1%
#712250000000
0!
0%
#712255000000
1!
1%
#712260000000
0!
0%
#712265000000
1!
1%
#712270000000
0!
0%
#712275000000
1!
1%
#712280000000
0!
0%
#712285000000
1!
1%
#712290000000
0!
0%
#712295000000
1!
1%
#712300000000
0!
0%
#712305000000
1!
1%
#712310000000
0!
0%
#712315000000
1!
1%
#712320000000
0!
0%
#712325000000
1!
1%
#712330000000
0!
0%
#712335000000
1!
1%
#712340000000
0!
0%
#712345000000
1!
1%
#712350000000
0!
0%
#712355000000
1!
1%
#712360000000
0!
0%
#712365000000
1!
1%
#712370000000
0!
0%
#712375000000
1!
1%
#712380000000
0!
0%
#712385000000
1!
1%
#712390000000
0!
0%
#712395000000
1!
1%
#712400000000
0!
0%
#712405000000
1!
1%
#712410000000
0!
0%
#712415000000
1!
1%
#712420000000
0!
0%
#712425000000
1!
1%
#712430000000
0!
0%
#712435000000
1!
1%
#712440000000
0!
0%
#712445000000
1!
1%
#712450000000
0!
0%
#712455000000
1!
1%
#712460000000
0!
0%
#712465000000
1!
1%
#712470000000
0!
0%
#712475000000
1!
1%
#712480000000
0!
0%
#712485000000
1!
1%
#712490000000
0!
0%
#712495000000
1!
1%
#712500000000
0!
0%
#712505000000
1!
1%
#712510000000
0!
0%
#712515000000
1!
1%
#712520000000
0!
0%
#712525000000
1!
1%
#712530000000
0!
0%
#712535000000
1!
1%
#712540000000
0!
0%
#712545000000
1!
1%
#712550000000
0!
0%
#712555000000
1!
1%
#712560000000
0!
0%
#712565000000
1!
1%
#712570000000
0!
0%
#712575000000
1!
1%
#712580000000
0!
0%
#712585000000
1!
1%
#712590000000
0!
0%
#712595000000
1!
1%
#712600000000
0!
0%
#712605000000
1!
1%
#712610000000
0!
0%
#712615000000
1!
1%
#712620000000
0!
0%
#712625000000
1!
1%
#712630000000
0!
0%
#712635000000
1!
1%
#712640000000
0!
0%
#712645000000
1!
1%
#712650000000
0!
0%
#712655000000
1!
1%
#712660000000
0!
0%
#712665000000
1!
1%
#712670000000
0!
0%
#712675000000
1!
1%
#712680000000
0!
0%
#712685000000
1!
1%
#712690000000
0!
0%
#712695000000
1!
1%
#712700000000
0!
0%
#712705000000
1!
1%
#712710000000
0!
0%
#712715000000
1!
1%
#712720000000
0!
0%
#712725000000
1!
1%
#712730000000
0!
0%
#712735000000
1!
1%
#712740000000
0!
0%
#712745000000
1!
1%
#712750000000
0!
0%
#712755000000
1!
1%
#712760000000
0!
0%
#712765000000
1!
1%
#712770000000
0!
0%
#712775000000
1!
1%
#712780000000
0!
0%
#712785000000
1!
1%
#712790000000
0!
0%
#712795000000
1!
1%
#712800000000
0!
0%
#712805000000
1!
1%
#712810000000
0!
0%
#712815000000
1!
1%
#712820000000
0!
0%
#712825000000
1!
1%
#712830000000
0!
0%
#712835000000
1!
1%
#712840000000
0!
0%
#712845000000
1!
1%
#712850000000
0!
0%
#712855000000
1!
1%
#712860000000
0!
0%
#712865000000
1!
1%
#712870000000
0!
0%
#712875000000
1!
1%
#712880000000
0!
0%
#712885000000
1!
1%
#712890000000
0!
0%
#712895000000
1!
1%
#712900000000
0!
0%
#712905000000
1!
1%
#712910000000
0!
0%
#712915000000
1!
1%
#712920000000
0!
0%
#712925000000
1!
1%
#712930000000
0!
0%
#712935000000
1!
1%
#712940000000
0!
0%
#712945000000
1!
1%
#712950000000
0!
0%
#712955000000
1!
1%
#712960000000
0!
0%
#712965000000
1!
1%
#712970000000
0!
0%
#712975000000
1!
1%
#712980000000
0!
0%
#712985000000
1!
1%
#712990000000
0!
0%
#712995000000
1!
1%
#713000000000
0!
0%
#713005000000
1!
1%
#713010000000
0!
0%
#713015000000
1!
1%
#713020000000
0!
0%
#713025000000
1!
1%
#713030000000
0!
0%
#713035000000
1!
1%
#713040000000
0!
0%
#713045000000
1!
1%
#713050000000
0!
0%
#713055000000
1!
1%
#713060000000
0!
0%
#713065000000
1!
1%
#713070000000
0!
0%
#713075000000
1!
1%
#713080000000
0!
0%
#713085000000
1!
1%
#713090000000
0!
0%
#713095000000
1!
1%
#713100000000
0!
0%
#713105000000
1!
1%
#713110000000
0!
0%
#713115000000
1!
1%
#713120000000
0!
0%
#713125000000
1!
1%
#713130000000
0!
0%
#713135000000
1!
1%
#713140000000
0!
0%
#713145000000
1!
1%
#713150000000
0!
0%
#713155000000
1!
1%
#713160000000
0!
0%
#713165000000
1!
1%
#713170000000
0!
0%
#713175000000
1!
1%
#713180000000
0!
0%
#713185000000
1!
1%
#713190000000
0!
0%
#713195000000
1!
1%
#713200000000
0!
0%
#713205000000
1!
1%
#713210000000
0!
0%
#713215000000
1!
1%
#713220000000
0!
0%
#713225000000
1!
1%
#713230000000
0!
0%
#713235000000
1!
1%
#713240000000
0!
0%
#713245000000
1!
1%
#713250000000
0!
0%
#713255000000
1!
1%
#713260000000
0!
0%
#713265000000
1!
1%
#713270000000
0!
0%
#713275000000
1!
1%
#713280000000
0!
0%
#713285000000
1!
1%
#713290000000
0!
0%
#713295000000
1!
1%
#713300000000
0!
0%
#713305000000
1!
1%
#713310000000
0!
0%
#713315000000
1!
1%
#713320000000
0!
0%
#713325000000
1!
1%
#713330000000
0!
0%
#713335000000
1!
1%
#713340000000
0!
0%
#713345000000
1!
1%
#713350000000
0!
0%
#713355000000
1!
1%
#713360000000
0!
0%
#713365000000
1!
1%
#713370000000
0!
0%
#713375000000
1!
1%
#713380000000
0!
0%
#713385000000
1!
1%
#713390000000
0!
0%
#713395000000
1!
1%
#713400000000
0!
0%
#713405000000
1!
1%
#713410000000
0!
0%
#713415000000
1!
1%
#713420000000
0!
0%
#713425000000
1!
1%
#713430000000
0!
0%
#713435000000
1!
1%
#713440000000
0!
0%
#713445000000
1!
1%
#713450000000
0!
0%
#713455000000
1!
1%
#713460000000
0!
0%
#713465000000
1!
1%
#713470000000
0!
0%
#713475000000
1!
1%
#713480000000
0!
0%
#713485000000
1!
1%
#713490000000
0!
0%
#713495000000
1!
1%
#713500000000
0!
0%
#713505000000
1!
1%
#713510000000
0!
0%
#713515000000
1!
1%
#713520000000
0!
0%
#713525000000
1!
1%
#713530000000
0!
0%
#713535000000
1!
1%
#713540000000
0!
0%
#713545000000
1!
1%
#713550000000
0!
0%
#713555000000
1!
1%
#713560000000
0!
0%
#713565000000
1!
1%
#713570000000
0!
0%
#713575000000
1!
1%
#713580000000
0!
0%
#713585000000
1!
1%
#713590000000
0!
0%
#713595000000
1!
1%
#713600000000
0!
0%
#713605000000
1!
1%
#713610000000
0!
0%
#713615000000
1!
1%
#713620000000
0!
0%
#713625000000
1!
1%
#713630000000
0!
0%
#713635000000
1!
1%
#713640000000
0!
0%
#713645000000
1!
1%
#713650000000
0!
0%
#713655000000
1!
1%
#713660000000
0!
0%
#713665000000
1!
1%
#713670000000
0!
0%
#713675000000
1!
1%
#713680000000
0!
0%
#713685000000
1!
1%
#713690000000
0!
0%
#713695000000
1!
1%
#713700000000
0!
0%
#713705000000
1!
1%
#713710000000
0!
0%
#713715000000
1!
1%
#713720000000
0!
0%
#713725000000
1!
1%
#713730000000
0!
0%
#713735000000
1!
1%
#713740000000
0!
0%
#713745000000
1!
1%
#713750000000
0!
0%
#713755000000
1!
1%
#713760000000
0!
0%
#713765000000
1!
1%
#713770000000
0!
0%
#713775000000
1!
1%
#713780000000
0!
0%
#713785000000
1!
1%
#713790000000
0!
0%
#713795000000
1!
1%
#713800000000
0!
0%
#713805000000
1!
1%
#713810000000
0!
0%
#713815000000
1!
1%
#713820000000
0!
0%
#713825000000
1!
1%
#713830000000
0!
0%
#713835000000
1!
1%
#713840000000
0!
0%
#713845000000
1!
1%
#713850000000
0!
0%
#713855000000
1!
1%
#713860000000
0!
0%
#713865000000
1!
1%
#713870000000
0!
0%
#713875000000
1!
1%
#713880000000
0!
0%
#713885000000
1!
1%
#713890000000
0!
0%
#713895000000
1!
1%
#713900000000
0!
0%
#713905000000
1!
1%
#713910000000
0!
0%
#713915000000
1!
1%
#713920000000
0!
0%
#713925000000
1!
1%
#713930000000
0!
0%
#713935000000
1!
1%
#713940000000
0!
0%
#713945000000
1!
1%
#713950000000
0!
0%
#713955000000
1!
1%
#713960000000
0!
0%
#713965000000
1!
1%
#713970000000
0!
0%
#713975000000
1!
1%
#713980000000
0!
0%
#713985000000
1!
1%
#713990000000
0!
0%
#713995000000
1!
1%
#714000000000
0!
0%
#714005000000
1!
1%
#714010000000
0!
0%
#714015000000
1!
1%
#714020000000
0!
0%
#714025000000
1!
1%
#714030000000
0!
0%
#714035000000
1!
1%
#714040000000
0!
0%
#714045000000
1!
1%
#714050000000
0!
0%
#714055000000
1!
1%
#714060000000
0!
0%
#714065000000
1!
1%
#714070000000
0!
0%
#714075000000
1!
1%
#714080000000
0!
0%
#714085000000
1!
1%
#714090000000
0!
0%
#714095000000
1!
1%
#714100000000
0!
0%
#714105000000
1!
1%
#714110000000
0!
0%
#714115000000
1!
1%
#714120000000
0!
0%
#714125000000
1!
1%
#714130000000
0!
0%
#714135000000
1!
1%
#714140000000
0!
0%
#714145000000
1!
1%
#714150000000
0!
0%
#714155000000
1!
1%
#714160000000
0!
0%
#714165000000
1!
1%
#714170000000
0!
0%
#714175000000
1!
1%
#714180000000
0!
0%
#714185000000
1!
1%
#714190000000
0!
0%
#714195000000
1!
1%
#714200000000
0!
0%
#714205000000
1!
1%
#714210000000
0!
0%
#714215000000
1!
1%
#714220000000
0!
0%
#714225000000
1!
1%
#714230000000
0!
0%
#714235000000
1!
1%
#714240000000
0!
0%
#714245000000
1!
1%
#714250000000
0!
0%
#714255000000
1!
1%
#714260000000
0!
0%
#714265000000
1!
1%
#714270000000
0!
0%
#714275000000
1!
1%
#714280000000
0!
0%
#714285000000
1!
1%
#714290000000
0!
0%
#714295000000
1!
1%
#714300000000
0!
0%
#714305000000
1!
1%
#714310000000
0!
0%
#714315000000
1!
1%
#714320000000
0!
0%
#714325000000
1!
1%
#714330000000
0!
0%
#714335000000
1!
1%
#714340000000
0!
0%
#714345000000
1!
1%
#714350000000
0!
0%
#714355000000
1!
1%
#714360000000
0!
0%
#714365000000
1!
1%
#714370000000
0!
0%
#714375000000
1!
1%
#714380000000
0!
0%
#714385000000
1!
1%
#714390000000
0!
0%
#714395000000
1!
1%
#714400000000
0!
0%
#714405000000
1!
1%
#714410000000
0!
0%
#714415000000
1!
1%
#714420000000
0!
0%
#714425000000
1!
1%
#714430000000
0!
0%
#714435000000
1!
1%
#714440000000
0!
0%
#714445000000
1!
1%
#714450000000
0!
0%
#714455000000
1!
1%
#714460000000
0!
0%
#714465000000
1!
1%
#714470000000
0!
0%
#714475000000
1!
1%
#714480000000
0!
0%
#714485000000
1!
1%
#714490000000
0!
0%
#714495000000
1!
1%
#714500000000
0!
0%
#714505000000
1!
1%
#714510000000
0!
0%
#714515000000
1!
1%
#714520000000
0!
0%
#714525000000
1!
1%
#714530000000
0!
0%
#714535000000
1!
1%
#714540000000
0!
0%
#714545000000
1!
1%
#714550000000
0!
0%
#714555000000
1!
1%
#714560000000
0!
0%
#714565000000
1!
1%
#714570000000
0!
0%
#714575000000
1!
1%
#714580000000
0!
0%
#714585000000
1!
1%
#714590000000
0!
0%
#714595000000
1!
1%
#714600000000
0!
0%
#714605000000
1!
1%
#714610000000
0!
0%
#714615000000
1!
1%
#714620000000
0!
0%
#714625000000
1!
1%
#714630000000
0!
0%
#714635000000
1!
1%
#714640000000
0!
0%
#714645000000
1!
1%
#714650000000
0!
0%
#714655000000
1!
1%
#714660000000
0!
0%
#714665000000
1!
1%
#714670000000
0!
0%
#714675000000
1!
1%
#714680000000
0!
0%
#714685000000
1!
1%
#714690000000
0!
0%
#714695000000
1!
1%
#714700000000
0!
0%
#714705000000
1!
1%
#714710000000
0!
0%
#714715000000
1!
1%
#714720000000
0!
0%
#714725000000
1!
1%
#714730000000
0!
0%
#714735000000
1!
1%
#714740000000
0!
0%
#714745000000
1!
1%
#714750000000
0!
0%
#714755000000
1!
1%
#714760000000
0!
0%
#714765000000
1!
1%
#714770000000
0!
0%
#714775000000
1!
1%
#714780000000
0!
0%
#714785000000
1!
1%
#714790000000
0!
0%
#714795000000
1!
1%
#714800000000
0!
0%
#714805000000
1!
1%
#714810000000
0!
0%
#714815000000
1!
1%
#714820000000
0!
0%
#714825000000
1!
1%
#714830000000
0!
0%
#714835000000
1!
1%
#714840000000
0!
0%
#714845000000
1!
1%
#714850000000
0!
0%
#714855000000
1!
1%
#714860000000
0!
0%
#714865000000
1!
1%
#714870000000
0!
0%
#714875000000
1!
1%
#714880000000
0!
0%
#714885000000
1!
1%
#714890000000
0!
0%
#714895000000
1!
1%
#714900000000
0!
0%
#714905000000
1!
1%
#714910000000
0!
0%
#714915000000
1!
1%
#714920000000
0!
0%
#714925000000
1!
1%
#714930000000
0!
0%
#714935000000
1!
1%
#714940000000
0!
0%
#714945000000
1!
1%
#714950000000
0!
0%
#714955000000
1!
1%
#714960000000
0!
0%
#714965000000
1!
1%
#714970000000
0!
0%
#714975000000
1!
1%
#714980000000
0!
0%
#714985000000
1!
1%
#714990000000
0!
0%
#714995000000
1!
1%
#715000000000
0!
0%
#715005000000
1!
1%
#715010000000
0!
0%
#715015000000
1!
1%
#715020000000
0!
0%
#715025000000
1!
1%
#715030000000
0!
0%
#715035000000
1!
1%
#715040000000
0!
0%
#715045000000
1!
1%
#715050000000
0!
0%
#715055000000
1!
1%
#715060000000
0!
0%
#715065000000
1!
1%
#715070000000
0!
0%
#715075000000
1!
1%
#715080000000
0!
0%
#715085000000
1!
1%
#715090000000
0!
0%
#715095000000
1!
1%
#715100000000
0!
0%
#715105000000
1!
1%
#715110000000
0!
0%
#715115000000
1!
1%
#715120000000
0!
0%
#715125000000
1!
1%
#715130000000
0!
0%
#715135000000
1!
1%
#715140000000
0!
0%
#715145000000
1!
1%
#715150000000
0!
0%
#715155000000
1!
1%
#715160000000
0!
0%
#715165000000
1!
1%
#715170000000
0!
0%
#715175000000
1!
1%
#715180000000
0!
0%
#715185000000
1!
1%
#715190000000
0!
0%
#715195000000
1!
1%
#715200000000
0!
0%
#715205000000
1!
1%
#715210000000
0!
0%
#715215000000
1!
1%
#715220000000
0!
0%
#715225000000
1!
1%
#715230000000
0!
0%
#715235000000
1!
1%
#715240000000
0!
0%
#715245000000
1!
1%
#715250000000
0!
0%
#715255000000
1!
1%
#715260000000
0!
0%
#715265000000
1!
1%
#715270000000
0!
0%
#715275000000
1!
1%
#715280000000
0!
0%
#715285000000
1!
1%
#715290000000
0!
0%
#715295000000
1!
1%
#715300000000
0!
0%
#715305000000
1!
1%
#715310000000
0!
0%
#715315000000
1!
1%
#715320000000
0!
0%
#715325000000
1!
1%
#715330000000
0!
0%
#715335000000
1!
1%
#715340000000
0!
0%
#715345000000
1!
1%
#715350000000
0!
0%
#715355000000
1!
1%
#715360000000
0!
0%
#715365000000
1!
1%
#715370000000
0!
0%
#715375000000
1!
1%
#715380000000
0!
0%
#715385000000
1!
1%
#715390000000
0!
0%
#715395000000
1!
1%
#715400000000
0!
0%
#715405000000
1!
1%
#715410000000
0!
0%
#715415000000
1!
1%
#715420000000
0!
0%
#715425000000
1!
1%
#715430000000
0!
0%
#715435000000
1!
1%
#715440000000
0!
0%
#715445000000
1!
1%
#715450000000
0!
0%
#715455000000
1!
1%
#715460000000
0!
0%
#715465000000
1!
1%
#715470000000
0!
0%
#715475000000
1!
1%
#715480000000
0!
0%
#715485000000
1!
1%
#715490000000
0!
0%
#715495000000
1!
1%
#715500000000
0!
0%
#715505000000
1!
1%
#715510000000
0!
0%
#715515000000
1!
1%
#715520000000
0!
0%
#715525000000
1!
1%
#715530000000
0!
0%
#715535000000
1!
1%
#715540000000
0!
0%
#715545000000
1!
1%
#715550000000
0!
0%
#715555000000
1!
1%
#715560000000
0!
0%
#715565000000
1!
1%
#715570000000
0!
0%
#715575000000
1!
1%
#715580000000
0!
0%
#715585000000
1!
1%
#715590000000
0!
0%
#715595000000
1!
1%
#715600000000
0!
0%
#715605000000
1!
1%
#715610000000
0!
0%
#715615000000
1!
1%
#715620000000
0!
0%
#715625000000
1!
1%
#715630000000
0!
0%
#715635000000
1!
1%
#715640000000
0!
0%
#715645000000
1!
1%
#715650000000
0!
0%
#715655000000
1!
1%
#715660000000
0!
0%
#715665000000
1!
1%
#715670000000
0!
0%
#715675000000
1!
1%
#715680000000
0!
0%
#715685000000
1!
1%
#715690000000
0!
0%
#715695000000
1!
1%
#715700000000
0!
0%
#715705000000
1!
1%
#715710000000
0!
0%
#715715000000
1!
1%
#715720000000
0!
0%
#715725000000
1!
1%
#715730000000
0!
0%
#715735000000
1!
1%
#715740000000
0!
0%
#715745000000
1!
1%
#715750000000
0!
0%
#715755000000
1!
1%
#715760000000
0!
0%
#715765000000
1!
1%
#715770000000
0!
0%
#715775000000
1!
1%
#715780000000
0!
0%
#715785000000
1!
1%
#715790000000
0!
0%
#715795000000
1!
1%
#715800000000
0!
0%
#715805000000
1!
1%
#715810000000
0!
0%
#715815000000
1!
1%
#715820000000
0!
0%
#715825000000
1!
1%
#715830000000
0!
0%
#715835000000
1!
1%
#715840000000
0!
0%
#715845000000
1!
1%
#715850000000
0!
0%
#715855000000
1!
1%
#715860000000
0!
0%
#715865000000
1!
1%
#715870000000
0!
0%
#715875000000
1!
1%
#715880000000
0!
0%
#715885000000
1!
1%
#715890000000
0!
0%
#715895000000
1!
1%
#715900000000
0!
0%
#715905000000
1!
1%
#715910000000
0!
0%
#715915000000
1!
1%
#715920000000
0!
0%
#715925000000
1!
1%
#715930000000
0!
0%
#715935000000
1!
1%
#715940000000
0!
0%
#715945000000
1!
1%
#715950000000
0!
0%
#715955000000
1!
1%
#715960000000
0!
0%
#715965000000
1!
1%
#715970000000
0!
0%
#715975000000
1!
1%
#715980000000
0!
0%
#715985000000
1!
1%
#715990000000
0!
0%
#715995000000
1!
1%
#716000000000
0!
0%
#716005000000
1!
1%
#716010000000
0!
0%
#716015000000
1!
1%
#716020000000
0!
0%
#716025000000
1!
1%
#716030000000
0!
0%
#716035000000
1!
1%
#716040000000
0!
0%
#716045000000
1!
1%
#716050000000
0!
0%
#716055000000
1!
1%
#716060000000
0!
0%
#716065000000
1!
1%
#716070000000
0!
0%
#716075000000
1!
1%
#716080000000
0!
0%
#716085000000
1!
1%
#716090000000
0!
0%
#716095000000
1!
1%
#716100000000
0!
0%
#716105000000
1!
1%
#716110000000
0!
0%
#716115000000
1!
1%
#716120000000
0!
0%
#716125000000
1!
1%
#716130000000
0!
0%
#716135000000
1!
1%
#716140000000
0!
0%
#716145000000
1!
1%
#716150000000
0!
0%
#716155000000
1!
1%
#716160000000
0!
0%
#716165000000
1!
1%
#716170000000
0!
0%
#716175000000
1!
1%
#716180000000
0!
0%
#716185000000
1!
1%
#716190000000
0!
0%
#716195000000
1!
1%
#716200000000
0!
0%
#716205000000
1!
1%
#716210000000
0!
0%
#716215000000
1!
1%
#716220000000
0!
0%
#716225000000
1!
1%
#716230000000
0!
0%
#716235000000
1!
1%
#716240000000
0!
0%
#716245000000
1!
1%
#716250000000
0!
0%
#716255000000
1!
1%
#716260000000
0!
0%
#716265000000
1!
1%
#716270000000
0!
0%
#716275000000
1!
1%
#716280000000
0!
0%
#716285000000
1!
1%
#716290000000
0!
0%
#716295000000
1!
1%
#716300000000
0!
0%
#716305000000
1!
1%
#716310000000
0!
0%
#716315000000
1!
1%
#716320000000
0!
0%
#716325000000
1!
1%
#716330000000
0!
0%
#716335000000
1!
1%
#716340000000
0!
0%
#716345000000
1!
1%
#716350000000
0!
0%
#716355000000
1!
1%
#716360000000
0!
0%
#716365000000
1!
1%
#716370000000
0!
0%
#716375000000
1!
1%
#716380000000
0!
0%
#716385000000
1!
1%
#716390000000
0!
0%
#716395000000
1!
1%
#716400000000
0!
0%
#716405000000
1!
1%
#716410000000
0!
0%
#716415000000
1!
1%
#716420000000
0!
0%
#716425000000
1!
1%
#716430000000
0!
0%
#716435000000
1!
1%
#716440000000
0!
0%
#716445000000
1!
1%
#716450000000
0!
0%
#716455000000
1!
1%
#716460000000
0!
0%
#716465000000
1!
1%
#716470000000
0!
0%
#716475000000
1!
1%
#716480000000
0!
0%
#716485000000
1!
1%
#716490000000
0!
0%
#716495000000
1!
1%
#716500000000
0!
0%
#716505000000
1!
1%
#716510000000
0!
0%
#716515000000
1!
1%
#716520000000
0!
0%
#716525000000
1!
1%
#716530000000
0!
0%
#716535000000
1!
1%
#716540000000
0!
0%
#716545000000
1!
1%
#716550000000
0!
0%
#716555000000
1!
1%
#716560000000
0!
0%
#716565000000
1!
1%
#716570000000
0!
0%
#716575000000
1!
1%
#716580000000
0!
0%
#716585000000
1!
1%
#716590000000
0!
0%
#716595000000
1!
1%
#716600000000
0!
0%
#716605000000
1!
1%
#716610000000
0!
0%
#716615000000
1!
1%
#716620000000
0!
0%
#716625000000
1!
1%
#716630000000
0!
0%
#716635000000
1!
1%
#716640000000
0!
0%
#716645000000
1!
1%
#716650000000
0!
0%
#716655000000
1!
1%
#716660000000
0!
0%
#716665000000
1!
1%
#716670000000
0!
0%
#716675000000
1!
1%
#716680000000
0!
0%
#716685000000
1!
1%
#716690000000
0!
0%
#716695000000
1!
1%
#716700000000
0!
0%
#716705000000
1!
1%
#716710000000
0!
0%
#716715000000
1!
1%
#716720000000
0!
0%
#716725000000
1!
1%
#716730000000
0!
0%
#716735000000
1!
1%
#716740000000
0!
0%
#716745000000
1!
1%
#716750000000
0!
0%
#716755000000
1!
1%
#716760000000
0!
0%
#716765000000
1!
1%
#716770000000
0!
0%
#716775000000
1!
1%
#716780000000
0!
0%
#716785000000
1!
1%
#716790000000
0!
0%
#716795000000
1!
1%
#716800000000
0!
0%
#716805000000
1!
1%
#716810000000
0!
0%
#716815000000
1!
1%
#716820000000
0!
0%
#716825000000
1!
1%
#716830000000
0!
0%
#716835000000
1!
1%
#716840000000
0!
0%
#716845000000
1!
1%
#716850000000
0!
0%
#716855000000
1!
1%
#716860000000
0!
0%
#716865000000
1!
1%
#716870000000
0!
0%
#716875000000
1!
1%
#716880000000
0!
0%
#716885000000
1!
1%
#716890000000
0!
0%
#716895000000
1!
1%
#716900000000
0!
0%
#716905000000
1!
1%
#716910000000
0!
0%
#716915000000
1!
1%
#716920000000
0!
0%
#716925000000
1!
1%
#716930000000
0!
0%
#716935000000
1!
1%
#716940000000
0!
0%
#716945000000
1!
1%
#716950000000
0!
0%
#716955000000
1!
1%
#716960000000
0!
0%
#716965000000
1!
1%
#716970000000
0!
0%
#716975000000
1!
1%
#716980000000
0!
0%
#716985000000
1!
1%
#716990000000
0!
0%
#716995000000
1!
1%
#717000000000
0!
0%
#717005000000
1!
1%
#717010000000
0!
0%
#717015000000
1!
1%
#717020000000
0!
0%
#717025000000
1!
1%
#717030000000
0!
0%
#717035000000
1!
1%
#717040000000
0!
0%
#717045000000
1!
1%
#717050000000
0!
0%
#717055000000
1!
1%
#717060000000
0!
0%
#717065000000
1!
1%
#717070000000
0!
0%
#717075000000
1!
1%
#717080000000
0!
0%
#717085000000
1!
1%
#717090000000
0!
0%
#717095000000
1!
1%
#717100000000
0!
0%
#717105000000
1!
1%
#717110000000
0!
0%
#717115000000
1!
1%
#717120000000
0!
0%
#717125000000
1!
1%
#717130000000
0!
0%
#717135000000
1!
1%
#717140000000
0!
0%
#717145000000
1!
1%
#717150000000
0!
0%
#717155000000
1!
1%
#717160000000
0!
0%
#717165000000
1!
1%
#717170000000
0!
0%
#717175000000
1!
1%
#717180000000
0!
0%
#717185000000
1!
1%
#717190000000
0!
0%
#717195000000
1!
1%
#717200000000
0!
0%
#717205000000
1!
1%
#717210000000
0!
0%
#717215000000
1!
1%
#717220000000
0!
0%
#717225000000
1!
1%
#717230000000
0!
0%
#717235000000
1!
1%
#717240000000
0!
0%
#717245000000
1!
1%
#717250000000
0!
0%
#717255000000
1!
1%
#717260000000
0!
0%
#717265000000
1!
1%
#717270000000
0!
0%
#717275000000
1!
1%
#717280000000
0!
0%
#717285000000
1!
1%
#717290000000
0!
0%
#717295000000
1!
1%
#717300000000
0!
0%
#717305000000
1!
1%
#717310000000
0!
0%
#717315000000
1!
1%
#717320000000
0!
0%
#717325000000
1!
1%
#717330000000
0!
0%
#717335000000
1!
1%
#717340000000
0!
0%
#717345000000
1!
1%
#717350000000
0!
0%
#717355000000
1!
1%
#717360000000
0!
0%
#717365000000
1!
1%
#717370000000
0!
0%
#717375000000
1!
1%
#717380000000
0!
0%
#717385000000
1!
1%
#717390000000
0!
0%
#717395000000
1!
1%
#717400000000
0!
0%
#717405000000
1!
1%
#717410000000
0!
0%
#717415000000
1!
1%
#717420000000
0!
0%
#717425000000
1!
1%
#717430000000
0!
0%
#717435000000
1!
1%
#717440000000
0!
0%
#717445000000
1!
1%
#717450000000
0!
0%
#717455000000
1!
1%
#717460000000
0!
0%
#717465000000
1!
1%
#717470000000
0!
0%
#717475000000
1!
1%
#717480000000
0!
0%
#717485000000
1!
1%
#717490000000
0!
0%
#717495000000
1!
1%
#717500000000
0!
0%
#717505000000
1!
1%
#717510000000
0!
0%
#717515000000
1!
1%
#717520000000
0!
0%
#717525000000
1!
1%
#717530000000
0!
0%
#717535000000
1!
1%
#717540000000
0!
0%
#717545000000
1!
1%
#717550000000
0!
0%
#717555000000
1!
1%
#717560000000
0!
0%
#717565000000
1!
1%
#717570000000
0!
0%
#717575000000
1!
1%
#717580000000
0!
0%
#717585000000
1!
1%
#717590000000
0!
0%
#717595000000
1!
1%
#717600000000
0!
0%
#717605000000
1!
1%
#717610000000
0!
0%
#717615000000
1!
1%
#717620000000
0!
0%
#717625000000
1!
1%
#717630000000
0!
0%
#717635000000
1!
1%
#717640000000
0!
0%
#717645000000
1!
1%
#717650000000
0!
0%
#717655000000
1!
1%
#717660000000
0!
0%
#717665000000
1!
1%
#717670000000
0!
0%
#717675000000
1!
1%
#717680000000
0!
0%
#717685000000
1!
1%
#717690000000
0!
0%
#717695000000
1!
1%
#717700000000
0!
0%
#717705000000
1!
1%
#717710000000
0!
0%
#717715000000
1!
1%
#717720000000
0!
0%
#717725000000
1!
1%
#717730000000
0!
0%
#717735000000
1!
1%
#717740000000
0!
0%
#717745000000
1!
1%
#717750000000
0!
0%
#717755000000
1!
1%
#717760000000
0!
0%
#717765000000
1!
1%
#717770000000
0!
0%
#717775000000
1!
1%
#717780000000
0!
0%
#717785000000
1!
1%
#717790000000
0!
0%
#717795000000
1!
1%
#717800000000
0!
0%
#717805000000
1!
1%
#717810000000
0!
0%
#717815000000
1!
1%
#717820000000
0!
0%
#717825000000
1!
1%
#717830000000
0!
0%
#717835000000
1!
1%
#717840000000
0!
0%
#717845000000
1!
1%
#717850000000
0!
0%
#717855000000
1!
1%
#717860000000
0!
0%
#717865000000
1!
1%
#717870000000
0!
0%
#717875000000
1!
1%
#717880000000
0!
0%
#717885000000
1!
1%
#717890000000
0!
0%
#717895000000
1!
1%
#717900000000
0!
0%
#717905000000
1!
1%
#717910000000
0!
0%
#717915000000
1!
1%
#717920000000
0!
0%
#717925000000
1!
1%
#717930000000
0!
0%
#717935000000
1!
1%
#717940000000
0!
0%
#717945000000
1!
1%
#717950000000
0!
0%
#717955000000
1!
1%
#717960000000
0!
0%
#717965000000
1!
1%
#717970000000
0!
0%
#717975000000
1!
1%
#717980000000
0!
0%
#717985000000
1!
1%
#717990000000
0!
0%
#717995000000
1!
1%
#718000000000
0!
0%
#718005000000
1!
1%
#718010000000
0!
0%
#718015000000
1!
1%
#718020000000
0!
0%
#718025000000
1!
1%
#718030000000
0!
0%
#718035000000
1!
1%
#718040000000
0!
0%
#718045000000
1!
1%
#718050000000
0!
0%
#718055000000
1!
1%
#718060000000
0!
0%
#718065000000
1!
1%
#718070000000
0!
0%
#718075000000
1!
1%
#718080000000
0!
0%
#718085000000
1!
1%
#718090000000
0!
0%
#718095000000
1!
1%
#718100000000
0!
0%
#718105000000
1!
1%
#718110000000
0!
0%
#718115000000
1!
1%
#718120000000
0!
0%
#718125000000
1!
1%
#718130000000
0!
0%
#718135000000
1!
1%
#718140000000
0!
0%
#718145000000
1!
1%
#718150000000
0!
0%
#718155000000
1!
1%
#718160000000
0!
0%
#718165000000
1!
1%
#718170000000
0!
0%
#718175000000
1!
1%
#718180000000
0!
0%
#718185000000
1!
1%
#718190000000
0!
0%
#718195000000
1!
1%
#718200000000
0!
0%
#718205000000
1!
1%
#718210000000
0!
0%
#718215000000
1!
1%
#718220000000
0!
0%
#718225000000
1!
1%
#718230000000
0!
0%
#718235000000
1!
1%
#718240000000
0!
0%
#718245000000
1!
1%
#718250000000
0!
0%
#718255000000
1!
1%
#718260000000
0!
0%
#718265000000
1!
1%
#718270000000
0!
0%
#718275000000
1!
1%
#718280000000
0!
0%
#718285000000
1!
1%
#718290000000
0!
0%
#718295000000
1!
1%
#718300000000
0!
0%
#718305000000
1!
1%
#718310000000
0!
0%
#718315000000
1!
1%
#718320000000
0!
0%
#718325000000
1!
1%
#718330000000
0!
0%
#718335000000
1!
1%
#718340000000
0!
0%
#718345000000
1!
1%
#718350000000
0!
0%
#718355000000
1!
1%
#718360000000
0!
0%
#718365000000
1!
1%
#718370000000
0!
0%
#718375000000
1!
1%
#718380000000
0!
0%
#718385000000
1!
1%
#718390000000
0!
0%
#718395000000
1!
1%
#718400000000
0!
0%
#718405000000
1!
1%
#718410000000
0!
0%
#718415000000
1!
1%
#718420000000
0!
0%
#718425000000
1!
1%
#718430000000
0!
0%
#718435000000
1!
1%
#718440000000
0!
0%
#718445000000
1!
1%
#718450000000
0!
0%
#718455000000
1!
1%
#718460000000
0!
0%
#718465000000
1!
1%
#718470000000
0!
0%
#718475000000
1!
1%
#718480000000
0!
0%
#718485000000
1!
1%
#718490000000
0!
0%
#718495000000
1!
1%
#718500000000
0!
0%
#718505000000
1!
1%
#718510000000
0!
0%
#718515000000
1!
1%
#718520000000
0!
0%
#718525000000
1!
1%
#718530000000
0!
0%
#718535000000
1!
1%
#718540000000
0!
0%
#718545000000
1!
1%
#718550000000
0!
0%
#718555000000
1!
1%
#718560000000
0!
0%
#718565000000
1!
1%
#718570000000
0!
0%
#718575000000
1!
1%
#718580000000
0!
0%
#718585000000
1!
1%
#718590000000
0!
0%
#718595000000
1!
1%
#718600000000
0!
0%
#718605000000
1!
1%
#718610000000
0!
0%
#718615000000
1!
1%
#718620000000
0!
0%
#718625000000
1!
1%
#718630000000
0!
0%
#718635000000
1!
1%
#718640000000
0!
0%
#718645000000
1!
1%
#718650000000
0!
0%
#718655000000
1!
1%
#718660000000
0!
0%
#718665000000
1!
1%
#718670000000
0!
0%
#718675000000
1!
1%
#718680000000
0!
0%
#718685000000
1!
1%
#718690000000
0!
0%
#718695000000
1!
1%
#718700000000
0!
0%
#718705000000
1!
1%
#718710000000
0!
0%
#718715000000
1!
1%
#718720000000
0!
0%
#718725000000
1!
1%
#718730000000
0!
0%
#718735000000
1!
1%
#718740000000
0!
0%
#718745000000
1!
1%
#718750000000
0!
0%
#718755000000
1!
1%
#718760000000
0!
0%
#718765000000
1!
1%
#718770000000
0!
0%
#718775000000
1!
1%
#718780000000
0!
0%
#718785000000
1!
1%
#718790000000
0!
0%
#718795000000
1!
1%
#718800000000
0!
0%
#718805000000
1!
1%
#718810000000
0!
0%
#718815000000
1!
1%
#718820000000
0!
0%
#718825000000
1!
1%
#718830000000
0!
0%
#718835000000
1!
1%
#718840000000
0!
0%
#718845000000
1!
1%
#718850000000
0!
0%
#718855000000
1!
1%
#718860000000
0!
0%
#718865000000
1!
1%
#718870000000
0!
0%
#718875000000
1!
1%
#718880000000
0!
0%
#718885000000
1!
1%
#718890000000
0!
0%
#718895000000
1!
1%
#718900000000
0!
0%
#718905000000
1!
1%
#718910000000
0!
0%
#718915000000
1!
1%
#718920000000
0!
0%
#718925000000
1!
1%
#718930000000
0!
0%
#718935000000
1!
1%
#718940000000
0!
0%
#718945000000
1!
1%
#718950000000
0!
0%
#718955000000
1!
1%
#718960000000
0!
0%
#718965000000
1!
1%
#718970000000
0!
0%
#718975000000
1!
1%
#718980000000
0!
0%
#718985000000
1!
1%
#718990000000
0!
0%
#718995000000
1!
1%
#719000000000
0!
0%
#719005000000
1!
1%
#719010000000
0!
0%
#719015000000
1!
1%
#719020000000
0!
0%
#719025000000
1!
1%
#719030000000
0!
0%
#719035000000
1!
1%
#719040000000
0!
0%
#719045000000
1!
1%
#719050000000
0!
0%
#719055000000
1!
1%
#719060000000
0!
0%
#719065000000
1!
1%
#719070000000
0!
0%
#719075000000
1!
1%
#719080000000
0!
0%
#719085000000
1!
1%
#719090000000
0!
0%
#719095000000
1!
1%
#719100000000
0!
0%
#719105000000
1!
1%
#719110000000
0!
0%
#719115000000
1!
1%
#719120000000
0!
0%
#719125000000
1!
1%
#719130000000
0!
0%
#719135000000
1!
1%
#719140000000
0!
0%
#719145000000
1!
1%
#719150000000
0!
0%
#719155000000
1!
1%
#719160000000
0!
0%
#719165000000
1!
1%
#719170000000
0!
0%
#719175000000
1!
1%
#719180000000
0!
0%
#719185000000
1!
1%
#719190000000
0!
0%
#719195000000
1!
1%
#719200000000
0!
0%
#719205000000
1!
1%
#719210000000
0!
0%
#719215000000
1!
1%
#719220000000
0!
0%
#719225000000
1!
1%
#719230000000
0!
0%
#719235000000
1!
1%
#719240000000
0!
0%
#719245000000
1!
1%
#719250000000
0!
0%
#719255000000
1!
1%
#719260000000
0!
0%
#719265000000
1!
1%
#719270000000
0!
0%
#719275000000
1!
1%
#719280000000
0!
0%
#719285000000
1!
1%
#719290000000
0!
0%
#719295000000
1!
1%
#719300000000
0!
0%
#719305000000
1!
1%
#719310000000
0!
0%
#719315000000
1!
1%
#719320000000
0!
0%
#719325000000
1!
1%
#719330000000
0!
0%
#719335000000
1!
1%
#719340000000
0!
0%
#719345000000
1!
1%
#719350000000
0!
0%
#719355000000
1!
1%
#719360000000
0!
0%
#719365000000
1!
1%
#719370000000
0!
0%
#719375000000
1!
1%
#719380000000
0!
0%
#719385000000
1!
1%
#719390000000
0!
0%
#719395000000
1!
1%
#719400000000
0!
0%
#719405000000
1!
1%
#719410000000
0!
0%
#719415000000
1!
1%
#719420000000
0!
0%
#719425000000
1!
1%
#719430000000
0!
0%
#719435000000
1!
1%
#719440000000
0!
0%
#719445000000
1!
1%
#719450000000
0!
0%
#719455000000
1!
1%
#719460000000
0!
0%
#719465000000
1!
1%
#719470000000
0!
0%
#719475000000
1!
1%
#719480000000
0!
0%
#719485000000
1!
1%
#719490000000
0!
0%
#719495000000
1!
1%
#719500000000
0!
0%
#719505000000
1!
1%
#719510000000
0!
0%
#719515000000
1!
1%
#719520000000
0!
0%
#719525000000
1!
1%
#719530000000
0!
0%
#719535000000
1!
1%
#719540000000
0!
0%
#719545000000
1!
1%
#719550000000
0!
0%
#719555000000
1!
1%
#719560000000
0!
0%
#719565000000
1!
1%
#719570000000
0!
0%
#719575000000
1!
1%
#719580000000
0!
0%
#719585000000
1!
1%
#719590000000
0!
0%
#719595000000
1!
1%
#719600000000
0!
0%
#719605000000
1!
1%
#719610000000
0!
0%
#719615000000
1!
1%
#719620000000
0!
0%
#719625000000
1!
1%
#719630000000
0!
0%
#719635000000
1!
1%
#719640000000
0!
0%
#719645000000
1!
1%
#719650000000
0!
0%
#719655000000
1!
1%
#719660000000
0!
0%
#719665000000
1!
1%
#719670000000
0!
0%
#719675000000
1!
1%
#719680000000
0!
0%
#719685000000
1!
1%
#719690000000
0!
0%
#719695000000
1!
1%
#719700000000
0!
0%
#719705000000
1!
1%
#719710000000
0!
0%
#719715000000
1!
1%
#719720000000
0!
0%
#719725000000
1!
1%
#719730000000
0!
0%
#719735000000
1!
1%
#719740000000
0!
0%
#719745000000
1!
1%
#719750000000
0!
0%
#719755000000
1!
1%
#719760000000
0!
0%
#719765000000
1!
1%
#719770000000
0!
0%
#719775000000
1!
1%
#719780000000
0!
0%
#719785000000
1!
1%
#719790000000
0!
0%
#719795000000
1!
1%
#719800000000
0!
0%
#719805000000
1!
1%
#719810000000
0!
0%
#719815000000
1!
1%
#719820000000
0!
0%
#719825000000
1!
1%
#719830000000
0!
0%
#719835000000
1!
1%
#719840000000
0!
0%
#719845000000
1!
1%
#719850000000
0!
0%
#719855000000
1!
1%
#719860000000
0!
0%
#719865000000
1!
1%
#719870000000
0!
0%
#719875000000
1!
1%
#719880000000
0!
0%
#719885000000
1!
1%
#719890000000
0!
0%
#719895000000
1!
1%
#719900000000
0!
0%
#719905000000
1!
1%
#719910000000
0!
0%
#719915000000
1!
1%
#719920000000
0!
0%
#719925000000
1!
1%
#719930000000
0!
0%
#719935000000
1!
1%
#719940000000
0!
0%
#719945000000
1!
1%
#719950000000
0!
0%
#719955000000
1!
1%
#719960000000
0!
0%
#719965000000
1!
1%
#719970000000
0!
0%
#719975000000
1!
1%
#719980000000
0!
0%
#719985000000
1!
1%
#719990000000
0!
0%
#719995000000
1!
1%
#720000000000
0!
0%
#720005000000
1!
1%
#720010000000
0!
0%
#720015000000
1!
1%
#720020000000
0!
0%
#720025000000
1!
1%
#720030000000
0!
0%
#720035000000
1!
1%
#720040000000
0!
0%
#720045000000
1!
1%
#720050000000
0!
0%
#720055000000
1!
1%
#720060000000
0!
0%
#720065000000
1!
1%
#720070000000
0!
0%
#720075000000
1!
1%
#720080000000
0!
0%
#720085000000
1!
1%
#720090000000
0!
0%
#720095000000
1!
1%
#720100000000
0!
0%
#720105000000
1!
1%
#720110000000
0!
0%
#720115000000
1!
1%
#720120000000
0!
0%
#720125000000
1!
1%
#720130000000
0!
0%
#720135000000
1!
1%
#720140000000
0!
0%
#720145000000
1!
1%
#720150000000
0!
0%
#720155000000
1!
1%
#720160000000
0!
0%
#720165000000
1!
1%
#720170000000
0!
0%
#720175000000
1!
1%
#720180000000
0!
0%
#720185000000
1!
1%
#720190000000
0!
0%
#720195000000
1!
1%
#720200000000
0!
0%
#720205000000
1!
1%
#720210000000
0!
0%
#720215000000
1!
1%
#720220000000
0!
0%
#720225000000
1!
1%
#720230000000
0!
0%
#720235000000
1!
1%
#720240000000
0!
0%
#720245000000
1!
1%
#720250000000
0!
0%
#720255000000
1!
1%
#720260000000
0!
0%
#720265000000
1!
1%
#720270000000
0!
0%
#720275000000
1!
1%
#720280000000
0!
0%
#720285000000
1!
1%
#720290000000
0!
0%
#720295000000
1!
1%
#720300000000
0!
0%
#720305000000
1!
1%
#720310000000
0!
0%
#720315000000
1!
1%
#720320000000
0!
0%
#720325000000
1!
1%
#720330000000
0!
0%
#720335000000
1!
1%
#720340000000
0!
0%
#720345000000
1!
1%
#720350000000
0!
0%
#720355000000
1!
1%
#720360000000
0!
0%
#720365000000
1!
1%
#720370000000
0!
0%
#720375000000
1!
1%
#720380000000
0!
0%
#720385000000
1!
1%
#720390000000
0!
0%
#720395000000
1!
1%
#720400000000
0!
0%
#720405000000
1!
1%
#720410000000
0!
0%
#720415000000
1!
1%
#720420000000
0!
0%
#720425000000
1!
1%
#720430000000
0!
0%
#720435000000
1!
1%
#720440000000
0!
0%
#720445000000
1!
1%
#720450000000
0!
0%
#720455000000
1!
1%
#720460000000
0!
0%
#720465000000
1!
1%
#720470000000
0!
0%
#720475000000
1!
1%
#720480000000
0!
0%
#720485000000
1!
1%
#720490000000
0!
0%
#720495000000
1!
1%
#720500000000
0!
0%
#720505000000
1!
1%
#720510000000
0!
0%
#720515000000
1!
1%
#720520000000
0!
0%
#720525000000
1!
1%
#720530000000
0!
0%
#720535000000
1!
1%
#720540000000
0!
0%
#720545000000
1!
1%
#720550000000
0!
0%
#720555000000
1!
1%
#720560000000
0!
0%
#720565000000
1!
1%
#720570000000
0!
0%
#720575000000
1!
1%
#720580000000
0!
0%
#720585000000
1!
1%
#720590000000
0!
0%
#720595000000
1!
1%
#720600000000
0!
0%
#720605000000
1!
1%
#720610000000
0!
0%
#720615000000
1!
1%
#720620000000
0!
0%
#720625000000
1!
1%
#720630000000
0!
0%
#720635000000
1!
1%
#720640000000
0!
0%
#720645000000
1!
1%
#720650000000
0!
0%
#720655000000
1!
1%
#720660000000
0!
0%
#720665000000
1!
1%
#720670000000
0!
0%
#720675000000
1!
1%
#720680000000
0!
0%
#720685000000
1!
1%
#720690000000
0!
0%
#720695000000
1!
1%
#720700000000
0!
0%
#720705000000
1!
1%
#720710000000
0!
0%
#720715000000
1!
1%
#720720000000
0!
0%
#720725000000
1!
1%
#720730000000
0!
0%
#720735000000
1!
1%
#720740000000
0!
0%
#720745000000
1!
1%
#720750000000
0!
0%
#720755000000
1!
1%
#720760000000
0!
0%
#720765000000
1!
1%
#720770000000
0!
0%
#720775000000
1!
1%
#720780000000
0!
0%
#720785000000
1!
1%
#720790000000
0!
0%
#720795000000
1!
1%
#720800000000
0!
0%
#720805000000
1!
1%
#720810000000
0!
0%
#720815000000
1!
1%
#720820000000
0!
0%
#720825000000
1!
1%
#720830000000
0!
0%
#720835000000
1!
1%
#720840000000
0!
0%
#720845000000
1!
1%
#720850000000
0!
0%
#720855000000
1!
1%
#720860000000
0!
0%
#720865000000
1!
1%
#720870000000
0!
0%
#720875000000
1!
1%
#720880000000
0!
0%
#720885000000
1!
1%
#720890000000
0!
0%
#720895000000
1!
1%
#720900000000
0!
0%
#720905000000
1!
1%
#720910000000
0!
0%
#720915000000
1!
1%
#720920000000
0!
0%
#720925000000
1!
1%
#720930000000
0!
0%
#720935000000
1!
1%
#720940000000
0!
0%
#720945000000
1!
1%
#720950000000
0!
0%
#720955000000
1!
1%
#720960000000
0!
0%
#720965000000
1!
1%
#720970000000
0!
0%
#720975000000
1!
1%
#720980000000
0!
0%
#720985000000
1!
1%
#720990000000
0!
0%
#720995000000
1!
1%
#721000000000
0!
0%
#721005000000
1!
1%
#721010000000
0!
0%
#721015000000
1!
1%
#721020000000
0!
0%
#721025000000
1!
1%
#721030000000
0!
0%
#721035000000
1!
1%
#721040000000
0!
0%
#721045000000
1!
1%
#721050000000
0!
0%
#721055000000
1!
1%
#721060000000
0!
0%
#721065000000
1!
1%
#721070000000
0!
0%
#721075000000
1!
1%
#721080000000
0!
0%
#721085000000
1!
1%
#721090000000
0!
0%
#721095000000
1!
1%
#721100000000
0!
0%
#721105000000
1!
1%
#721110000000
0!
0%
#721115000000
1!
1%
#721120000000
0!
0%
#721125000000
1!
1%
#721130000000
0!
0%
#721135000000
1!
1%
#721140000000
0!
0%
#721145000000
1!
1%
#721150000000
0!
0%
#721155000000
1!
1%
#721160000000
0!
0%
#721165000000
1!
1%
#721170000000
0!
0%
#721175000000
1!
1%
#721180000000
0!
0%
#721185000000
1!
1%
#721190000000
0!
0%
#721195000000
1!
1%
#721200000000
0!
0%
#721205000000
1!
1%
#721210000000
0!
0%
#721215000000
1!
1%
#721220000000
0!
0%
#721225000000
1!
1%
#721230000000
0!
0%
#721235000000
1!
1%
#721240000000
0!
0%
#721245000000
1!
1%
#721250000000
0!
0%
#721255000000
1!
1%
#721260000000
0!
0%
#721265000000
1!
1%
#721270000000
0!
0%
#721275000000
1!
1%
#721280000000
0!
0%
#721285000000
1!
1%
#721290000000
0!
0%
#721295000000
1!
1%
#721300000000
0!
0%
#721305000000
1!
1%
#721310000000
0!
0%
#721315000000
1!
1%
#721320000000
0!
0%
#721325000000
1!
1%
#721330000000
0!
0%
#721335000000
1!
1%
#721340000000
0!
0%
#721345000000
1!
1%
#721350000000
0!
0%
#721355000000
1!
1%
#721360000000
0!
0%
#721365000000
1!
1%
#721370000000
0!
0%
#721375000000
1!
1%
#721380000000
0!
0%
#721385000000
1!
1%
#721390000000
0!
0%
#721395000000
1!
1%
#721400000000
0!
0%
#721405000000
1!
1%
#721410000000
0!
0%
#721415000000
1!
1%
#721420000000
0!
0%
#721425000000
1!
1%
#721430000000
0!
0%
#721435000000
1!
1%
#721440000000
0!
0%
#721445000000
1!
1%
#721450000000
0!
0%
#721455000000
1!
1%
#721460000000
0!
0%
#721465000000
1!
1%
#721470000000
0!
0%
#721475000000
1!
1%
#721480000000
0!
0%
#721485000000
1!
1%
#721490000000
0!
0%
#721495000000
1!
1%
#721500000000
0!
0%
#721505000000
1!
1%
#721510000000
0!
0%
#721515000000
1!
1%
#721520000000
0!
0%
#721525000000
1!
1%
#721530000000
0!
0%
#721535000000
1!
1%
#721540000000
0!
0%
#721545000000
1!
1%
#721550000000
0!
0%
#721555000000
1!
1%
#721560000000
0!
0%
#721565000000
1!
1%
#721570000000
0!
0%
#721575000000
1!
1%
#721580000000
0!
0%
#721585000000
1!
1%
#721590000000
0!
0%
#721595000000
1!
1%
#721600000000
0!
0%
#721605000000
1!
1%
#721610000000
0!
0%
#721615000000
1!
1%
#721620000000
0!
0%
#721625000000
1!
1%
#721630000000
0!
0%
#721635000000
1!
1%
#721640000000
0!
0%
#721645000000
1!
1%
#721650000000
0!
0%
#721655000000
1!
1%
#721660000000
0!
0%
#721665000000
1!
1%
#721670000000
0!
0%
#721675000000
1!
1%
#721680000000
0!
0%
#721685000000
1!
1%
#721690000000
0!
0%
#721695000000
1!
1%
#721700000000
0!
0%
#721705000000
1!
1%
#721710000000
0!
0%
#721715000000
1!
1%
#721720000000
0!
0%
#721725000000
1!
1%
#721730000000
0!
0%
#721735000000
1!
1%
#721740000000
0!
0%
#721745000000
1!
1%
#721750000000
0!
0%
#721755000000
1!
1%
#721760000000
0!
0%
#721765000000
1!
1%
#721770000000
0!
0%
#721775000000
1!
1%
#721780000000
0!
0%
#721785000000
1!
1%
#721790000000
0!
0%
#721795000000
1!
1%
#721800000000
0!
0%
#721805000000
1!
1%
#721810000000
0!
0%
#721815000000
1!
1%
#721820000000
0!
0%
#721825000000
1!
1%
#721830000000
0!
0%
#721835000000
1!
1%
#721840000000
0!
0%
#721845000000
1!
1%
#721850000000
0!
0%
#721855000000
1!
1%
#721860000000
0!
0%
#721865000000
1!
1%
#721870000000
0!
0%
#721875000000
1!
1%
#721880000000
0!
0%
#721885000000
1!
1%
#721890000000
0!
0%
#721895000000
1!
1%
#721900000000
0!
0%
#721905000000
1!
1%
#721910000000
0!
0%
#721915000000
1!
1%
#721920000000
0!
0%
#721925000000
1!
1%
#721930000000
0!
0%
#721935000000
1!
1%
#721940000000
0!
0%
#721945000000
1!
1%
#721950000000
0!
0%
#721955000000
1!
1%
#721960000000
0!
0%
#721965000000
1!
1%
#721970000000
0!
0%
#721975000000
1!
1%
#721980000000
0!
0%
#721985000000
1!
1%
#721990000000
0!
0%
#721995000000
1!
1%
#722000000000
0!
0%
#722005000000
1!
1%
#722010000000
0!
0%
#722015000000
1!
1%
#722020000000
0!
0%
#722025000000
1!
1%
#722030000000
0!
0%
#722035000000
1!
1%
#722040000000
0!
0%
#722045000000
1!
1%
#722050000000
0!
0%
#722055000000
1!
1%
#722060000000
0!
0%
#722065000000
1!
1%
#722070000000
0!
0%
#722075000000
1!
1%
#722080000000
0!
0%
#722085000000
1!
1%
#722090000000
0!
0%
#722095000000
1!
1%
#722100000000
0!
0%
#722105000000
1!
1%
#722110000000
0!
0%
#722115000000
1!
1%
#722120000000
0!
0%
#722125000000
1!
1%
#722130000000
0!
0%
#722135000000
1!
1%
#722140000000
0!
0%
#722145000000
1!
1%
#722150000000
0!
0%
#722155000000
1!
1%
#722160000000
0!
0%
#722165000000
1!
1%
#722170000000
0!
0%
#722175000000
1!
1%
#722180000000
0!
0%
#722185000000
1!
1%
#722190000000
0!
0%
#722195000000
1!
1%
#722200000000
0!
0%
#722205000000
1!
1%
#722210000000
0!
0%
#722215000000
1!
1%
#722220000000
0!
0%
#722225000000
1!
1%
#722230000000
0!
0%
#722235000000
1!
1%
#722240000000
0!
0%
#722245000000
1!
1%
#722250000000
0!
0%
#722255000000
1!
1%
#722260000000
0!
0%
#722265000000
1!
1%
#722270000000
0!
0%
#722275000000
1!
1%
#722280000000
0!
0%
#722285000000
1!
1%
#722290000000
0!
0%
#722295000000
1!
1%
#722300000000
0!
0%
#722305000000
1!
1%
#722310000000
0!
0%
#722315000000
1!
1%
#722320000000
0!
0%
#722325000000
1!
1%
#722330000000
0!
0%
#722335000000
1!
1%
#722340000000
0!
0%
#722345000000
1!
1%
#722350000000
0!
0%
#722355000000
1!
1%
#722360000000
0!
0%
#722365000000
1!
1%
#722370000000
0!
0%
#722375000000
1!
1%
#722380000000
0!
0%
#722385000000
1!
1%
#722390000000
0!
0%
#722395000000
1!
1%
#722400000000
0!
0%
#722405000000
1!
1%
#722410000000
0!
0%
#722415000000
1!
1%
#722420000000
0!
0%
#722425000000
1!
1%
#722430000000
0!
0%
#722435000000
1!
1%
#722440000000
0!
0%
#722445000000
1!
1%
#722450000000
0!
0%
#722455000000
1!
1%
#722460000000
0!
0%
#722465000000
1!
1%
#722470000000
0!
0%
#722475000000
1!
1%
#722480000000
0!
0%
#722485000000
1!
1%
#722490000000
0!
0%
#722495000000
1!
1%
#722500000000
0!
0%
#722505000000
1!
1%
#722510000000
0!
0%
#722515000000
1!
1%
#722520000000
0!
0%
#722525000000
1!
1%
#722530000000
0!
0%
#722535000000
1!
1%
#722540000000
0!
0%
#722545000000
1!
1%
#722550000000
0!
0%
#722555000000
1!
1%
#722560000000
0!
0%
#722565000000
1!
1%
#722570000000
0!
0%
#722575000000
1!
1%
#722580000000
0!
0%
#722585000000
1!
1%
#722590000000
0!
0%
#722595000000
1!
1%
#722600000000
0!
0%
#722605000000
1!
1%
#722610000000
0!
0%
#722615000000
1!
1%
#722620000000
0!
0%
#722625000000
1!
1%
#722630000000
0!
0%
#722635000000
1!
1%
#722640000000
0!
0%
#722645000000
1!
1%
#722650000000
0!
0%
#722655000000
1!
1%
#722660000000
0!
0%
#722665000000
1!
1%
#722670000000
0!
0%
#722675000000
1!
1%
#722680000000
0!
0%
#722685000000
1!
1%
#722690000000
0!
0%
#722695000000
1!
1%
#722700000000
0!
0%
#722705000000
1!
1%
#722710000000
0!
0%
#722715000000
1!
1%
#722720000000
0!
0%
#722725000000
1!
1%
#722730000000
0!
0%
#722735000000
1!
1%
#722740000000
0!
0%
#722745000000
1!
1%
#722750000000
0!
0%
#722755000000
1!
1%
#722760000000
0!
0%
#722765000000
1!
1%
#722770000000
0!
0%
#722775000000
1!
1%
#722780000000
0!
0%
#722785000000
1!
1%
#722790000000
0!
0%
#722795000000
1!
1%
#722800000000
0!
0%
#722805000000
1!
1%
#722810000000
0!
0%
#722815000000
1!
1%
#722820000000
0!
0%
#722825000000
1!
1%
#722830000000
0!
0%
#722835000000
1!
1%
#722840000000
0!
0%
#722845000000
1!
1%
#722850000000
0!
0%
#722855000000
1!
1%
#722860000000
0!
0%
#722865000000
1!
1%
#722870000000
0!
0%
#722875000000
1!
1%
#722880000000
0!
0%
#722885000000
1!
1%
#722890000000
0!
0%
#722895000000
1!
1%
#722900000000
0!
0%
#722905000000
1!
1%
#722910000000
0!
0%
#722915000000
1!
1%
#722920000000
0!
0%
#722925000000
1!
1%
#722930000000
0!
0%
#722935000000
1!
1%
#722940000000
0!
0%
#722945000000
1!
1%
#722950000000
0!
0%
#722955000000
1!
1%
#722960000000
0!
0%
#722965000000
1!
1%
#722970000000
0!
0%
#722975000000
1!
1%
#722980000000
0!
0%
#722985000000
1!
1%
#722990000000
0!
0%
#722995000000
1!
1%
#723000000000
0!
0%
#723005000000
1!
1%
#723010000000
0!
0%
#723015000000
1!
1%
#723020000000
0!
0%
#723025000000
1!
1%
#723030000000
0!
0%
#723035000000
1!
1%
#723040000000
0!
0%
#723045000000
1!
1%
#723050000000
0!
0%
#723055000000
1!
1%
#723060000000
0!
0%
#723065000000
1!
1%
#723070000000
0!
0%
#723075000000
1!
1%
#723080000000
0!
0%
#723085000000
1!
1%
#723090000000
0!
0%
#723095000000
1!
1%
#723100000000
0!
0%
#723105000000
1!
1%
#723110000000
0!
0%
#723115000000
1!
1%
#723120000000
0!
0%
#723125000000
1!
1%
#723130000000
0!
0%
#723135000000
1!
1%
#723140000000
0!
0%
#723145000000
1!
1%
#723150000000
0!
0%
#723155000000
1!
1%
#723160000000
0!
0%
#723165000000
1!
1%
#723170000000
0!
0%
#723175000000
1!
1%
#723180000000
0!
0%
#723185000000
1!
1%
#723190000000
0!
0%
#723195000000
1!
1%
#723200000000
0!
0%
#723205000000
1!
1%
#723210000000
0!
0%
#723215000000
1!
1%
#723220000000
0!
0%
#723225000000
1!
1%
#723230000000
0!
0%
#723235000000
1!
1%
#723240000000
0!
0%
#723245000000
1!
1%
#723250000000
0!
0%
#723255000000
1!
1%
#723260000000
0!
0%
#723265000000
1!
1%
#723270000000
0!
0%
#723275000000
1!
1%
#723280000000
0!
0%
#723285000000
1!
1%
#723290000000
0!
0%
#723295000000
1!
1%
#723300000000
0!
0%
#723305000000
1!
1%
#723310000000
0!
0%
#723315000000
1!
1%
#723320000000
0!
0%
#723325000000
1!
1%
#723330000000
0!
0%
#723335000000
1!
1%
#723340000000
0!
0%
#723345000000
1!
1%
#723350000000
0!
0%
#723355000000
1!
1%
#723360000000
0!
0%
#723365000000
1!
1%
#723370000000
0!
0%
#723375000000
1!
1%
#723380000000
0!
0%
#723385000000
1!
1%
#723390000000
0!
0%
#723395000000
1!
1%
#723400000000
0!
0%
#723405000000
1!
1%
#723410000000
0!
0%
#723415000000
1!
1%
#723420000000
0!
0%
#723425000000
1!
1%
#723430000000
0!
0%
#723435000000
1!
1%
#723440000000
0!
0%
#723445000000
1!
1%
#723450000000
0!
0%
#723455000000
1!
1%
#723460000000
0!
0%
#723465000000
1!
1%
#723470000000
0!
0%
#723475000000
1!
1%
#723480000000
0!
0%
#723485000000
1!
1%
#723490000000
0!
0%
#723495000000
1!
1%
#723500000000
0!
0%
#723505000000
1!
1%
#723510000000
0!
0%
#723515000000
1!
1%
#723520000000
0!
0%
#723525000000
1!
1%
#723530000000
0!
0%
#723535000000
1!
1%
#723540000000
0!
0%
#723545000000
1!
1%
#723550000000
0!
0%
#723555000000
1!
1%
#723560000000
0!
0%
#723565000000
1!
1%
#723570000000
0!
0%
#723575000000
1!
1%
#723580000000
0!
0%
#723585000000
1!
1%
#723590000000
0!
0%
#723595000000
1!
1%
#723600000000
0!
0%
#723605000000
1!
1%
#723610000000
0!
0%
#723615000000
1!
1%
#723620000000
0!
0%
#723625000000
1!
1%
#723630000000
0!
0%
#723635000000
1!
1%
#723640000000
0!
0%
#723645000000
1!
1%
#723650000000
0!
0%
#723655000000
1!
1%
#723660000000
0!
0%
#723665000000
1!
1%
#723670000000
0!
0%
#723675000000
1!
1%
#723680000000
0!
0%
#723685000000
1!
1%
#723690000000
0!
0%
#723695000000
1!
1%
#723700000000
0!
0%
#723705000000
1!
1%
#723710000000
0!
0%
#723715000000
1!
1%
#723720000000
0!
0%
#723725000000
1!
1%
#723730000000
0!
0%
#723735000000
1!
1%
#723740000000
0!
0%
#723745000000
1!
1%
#723750000000
0!
0%
#723755000000
1!
1%
#723760000000
0!
0%
#723765000000
1!
1%
#723770000000
0!
0%
#723775000000
1!
1%
#723780000000
0!
0%
#723785000000
1!
1%
#723790000000
0!
0%
#723795000000
1!
1%
#723800000000
0!
0%
#723805000000
1!
1%
#723810000000
0!
0%
#723815000000
1!
1%
#723820000000
0!
0%
#723825000000
1!
1%
#723830000000
0!
0%
#723835000000
1!
1%
#723840000000
0!
0%
#723845000000
1!
1%
#723850000000
0!
0%
#723855000000
1!
1%
#723860000000
0!
0%
#723865000000
1!
1%
#723870000000
0!
0%
#723875000000
1!
1%
#723880000000
0!
0%
#723885000000
1!
1%
#723890000000
0!
0%
#723895000000
1!
1%
#723900000000
0!
0%
#723905000000
1!
1%
#723910000000
0!
0%
#723915000000
1!
1%
#723920000000
0!
0%
#723925000000
1!
1%
#723930000000
0!
0%
#723935000000
1!
1%
#723940000000
0!
0%
#723945000000
1!
1%
#723950000000
0!
0%
#723955000000
1!
1%
#723960000000
0!
0%
#723965000000
1!
1%
#723970000000
0!
0%
#723975000000
1!
1%
#723980000000
0!
0%
#723985000000
1!
1%
#723990000000
0!
0%
#723995000000
1!
1%
#724000000000
0!
0%
#724005000000
1!
1%
#724010000000
0!
0%
#724015000000
1!
1%
#724020000000
0!
0%
#724025000000
1!
1%
#724030000000
0!
0%
#724035000000
1!
1%
#724040000000
0!
0%
#724045000000
1!
1%
#724050000000
0!
0%
#724055000000
1!
1%
#724060000000
0!
0%
#724065000000
1!
1%
#724070000000
0!
0%
#724075000000
1!
1%
#724080000000
0!
0%
#724085000000
1!
1%
#724090000000
0!
0%
#724095000000
1!
1%
#724100000000
0!
0%
#724105000000
1!
1%
#724110000000
0!
0%
#724115000000
1!
1%
#724120000000
0!
0%
#724125000000
1!
1%
#724130000000
0!
0%
#724135000000
1!
1%
#724140000000
0!
0%
#724145000000
1!
1%
#724150000000
0!
0%
#724155000000
1!
1%
#724160000000
0!
0%
#724165000000
1!
1%
#724170000000
0!
0%
#724175000000
1!
1%
#724180000000
0!
0%
#724185000000
1!
1%
#724190000000
0!
0%
#724195000000
1!
1%
#724200000000
0!
0%
#724205000000
1!
1%
#724210000000
0!
0%
#724215000000
1!
1%
#724220000000
0!
0%
#724225000000
1!
1%
#724230000000
0!
0%
#724235000000
1!
1%
#724240000000
0!
0%
#724245000000
1!
1%
#724250000000
0!
0%
#724255000000
1!
1%
#724260000000
0!
0%
#724265000000
1!
1%
#724270000000
0!
0%
#724275000000
1!
1%
#724280000000
0!
0%
#724285000000
1!
1%
#724290000000
0!
0%
#724295000000
1!
1%
#724300000000
0!
0%
#724305000000
1!
1%
#724310000000
0!
0%
#724315000000
1!
1%
#724320000000
0!
0%
#724325000000
1!
1%
#724330000000
0!
0%
#724335000000
1!
1%
#724340000000
0!
0%
#724345000000
1!
1%
#724350000000
0!
0%
#724355000000
1!
1%
#724360000000
0!
0%
#724365000000
1!
1%
#724370000000
0!
0%
#724375000000
1!
1%
#724380000000
0!
0%
#724385000000
1!
1%
#724390000000
0!
0%
#724395000000
1!
1%
#724400000000
0!
0%
#724405000000
1!
1%
#724410000000
0!
0%
#724415000000
1!
1%
#724420000000
0!
0%
#724425000000
1!
1%
#724430000000
0!
0%
#724435000000
1!
1%
#724440000000
0!
0%
#724445000000
1!
1%
#724450000000
0!
0%
#724455000000
1!
1%
#724460000000
0!
0%
#724465000000
1!
1%
#724470000000
0!
0%
#724475000000
1!
1%
#724480000000
0!
0%
#724485000000
1!
1%
#724490000000
0!
0%
#724495000000
1!
1%
#724500000000
0!
0%
#724505000000
1!
1%
#724510000000
0!
0%
#724515000000
1!
1%
#724520000000
0!
0%
#724525000000
1!
1%
#724530000000
0!
0%
#724535000000
1!
1%
#724540000000
0!
0%
#724545000000
1!
1%
#724550000000
0!
0%
#724555000000
1!
1%
#724560000000
0!
0%
#724565000000
1!
1%
#724570000000
0!
0%
#724575000000
1!
1%
#724580000000
0!
0%
#724585000000
1!
1%
#724590000000
0!
0%
#724595000000
1!
1%
#724600000000
0!
0%
#724605000000
1!
1%
#724610000000
0!
0%
#724615000000
1!
1%
#724620000000
0!
0%
#724625000000
1!
1%
#724630000000
0!
0%
#724635000000
1!
1%
#724640000000
0!
0%
#724645000000
1!
1%
#724650000000
0!
0%
#724655000000
1!
1%
#724660000000
0!
0%
#724665000000
1!
1%
#724670000000
0!
0%
#724675000000
1!
1%
#724680000000
0!
0%
#724685000000
1!
1%
#724690000000
0!
0%
#724695000000
1!
1%
#724700000000
0!
0%
#724705000000
1!
1%
#724710000000
0!
0%
#724715000000
1!
1%
#724720000000
0!
0%
#724725000000
1!
1%
#724730000000
0!
0%
#724735000000
1!
1%
#724740000000
0!
0%
#724745000000
1!
1%
#724750000000
0!
0%
#724755000000
1!
1%
#724760000000
0!
0%
#724765000000
1!
1%
#724770000000
0!
0%
#724775000000
1!
1%
#724780000000
0!
0%
#724785000000
1!
1%
#724790000000
0!
0%
#724795000000
1!
1%
#724800000000
0!
0%
#724805000000
1!
1%
#724810000000
0!
0%
#724815000000
1!
1%
#724820000000
0!
0%
#724825000000
1!
1%
#724830000000
0!
0%
#724835000000
1!
1%
#724840000000
0!
0%
#724845000000
1!
1%
#724850000000
0!
0%
#724855000000
1!
1%
#724860000000
0!
0%
#724865000000
1!
1%
#724870000000
0!
0%
#724875000000
1!
1%
#724880000000
0!
0%
#724885000000
1!
1%
#724890000000
0!
0%
#724895000000
1!
1%
#724900000000
0!
0%
#724905000000
1!
1%
#724910000000
0!
0%
#724915000000
1!
1%
#724920000000
0!
0%
#724925000000
1!
1%
#724930000000
0!
0%
#724935000000
1!
1%
#724940000000
0!
0%
#724945000000
1!
1%
#724950000000
0!
0%
#724955000000
1!
1%
#724960000000
0!
0%
#724965000000
1!
1%
#724970000000
0!
0%
#724975000000
1!
1%
#724980000000
0!
0%
#724985000000
1!
1%
#724990000000
0!
0%
#724995000000
1!
1%
#725000000000
0!
0%
#725005000000
1!
1%
#725010000000
0!
0%
#725015000000
1!
1%
#725020000000
0!
0%
#725025000000
1!
1%
#725030000000
0!
0%
#725035000000
1!
1%
#725040000000
0!
0%
#725045000000
1!
1%
#725050000000
0!
0%
#725055000000
1!
1%
#725060000000
0!
0%
#725065000000
1!
1%
#725070000000
0!
0%
#725075000000
1!
1%
#725080000000
0!
0%
#725085000000
1!
1%
#725090000000
0!
0%
#725095000000
1!
1%
#725100000000
0!
0%
#725105000000
1!
1%
#725110000000
0!
0%
#725115000000
1!
1%
#725120000000
0!
0%
#725125000000
1!
1%
#725130000000
0!
0%
#725135000000
1!
1%
#725140000000
0!
0%
#725145000000
1!
1%
#725150000000
0!
0%
#725155000000
1!
1%
#725160000000
0!
0%
#725165000000
1!
1%
#725170000000
0!
0%
#725175000000
1!
1%
#725180000000
0!
0%
#725185000000
1!
1%
#725190000000
0!
0%
#725195000000
1!
1%
#725200000000
0!
0%
#725205000000
1!
1%
#725210000000
0!
0%
#725215000000
1!
1%
#725220000000
0!
0%
#725225000000
1!
1%
#725230000000
0!
0%
#725235000000
1!
1%
#725240000000
0!
0%
#725245000000
1!
1%
#725250000000
0!
0%
#725255000000
1!
1%
#725260000000
0!
0%
#725265000000
1!
1%
#725270000000
0!
0%
#725275000000
1!
1%
#725280000000
0!
0%
#725285000000
1!
1%
#725290000000
0!
0%
#725295000000
1!
1%
#725300000000
0!
0%
#725305000000
1!
1%
#725310000000
0!
0%
#725315000000
1!
1%
#725320000000
0!
0%
#725325000000
1!
1%
#725330000000
0!
0%
#725335000000
1!
1%
#725340000000
0!
0%
#725345000000
1!
1%
#725350000000
0!
0%
#725355000000
1!
1%
#725360000000
0!
0%
#725365000000
1!
1%
#725370000000
0!
0%
#725375000000
1!
1%
#725380000000
0!
0%
#725385000000
1!
1%
#725390000000
0!
0%
#725395000000
1!
1%
#725400000000
0!
0%
#725405000000
1!
1%
#725410000000
0!
0%
#725415000000
1!
1%
#725420000000
0!
0%
#725425000000
1!
1%
#725430000000
0!
0%
#725435000000
1!
1%
#725440000000
0!
0%
#725445000000
1!
1%
#725450000000
0!
0%
#725455000000
1!
1%
#725460000000
0!
0%
#725465000000
1!
1%
#725470000000
0!
0%
#725475000000
1!
1%
#725480000000
0!
0%
#725485000000
1!
1%
#725490000000
0!
0%
#725495000000
1!
1%
#725500000000
0!
0%
#725505000000
1!
1%
#725510000000
0!
0%
#725515000000
1!
1%
#725520000000
0!
0%
#725525000000
1!
1%
#725530000000
0!
0%
#725535000000
1!
1%
#725540000000
0!
0%
#725545000000
1!
1%
#725550000000
0!
0%
#725555000000
1!
1%
#725560000000
0!
0%
#725565000000
1!
1%
#725570000000
0!
0%
#725575000000
1!
1%
#725580000000
0!
0%
#725585000000
1!
1%
#725590000000
0!
0%
#725595000000
1!
1%
#725600000000
0!
0%
#725605000000
1!
1%
#725610000000
0!
0%
#725615000000
1!
1%
#725620000000
0!
0%
#725625000000
1!
1%
#725630000000
0!
0%
#725635000000
1!
1%
#725640000000
0!
0%
#725645000000
1!
1%
#725650000000
0!
0%
#725655000000
1!
1%
#725660000000
0!
0%
#725665000000
1!
1%
#725670000000
0!
0%
#725675000000
1!
1%
#725680000000
0!
0%
#725685000000
1!
1%
#725690000000
0!
0%
#725695000000
1!
1%
#725700000000
0!
0%
#725705000000
1!
1%
#725710000000
0!
0%
#725715000000
1!
1%
#725720000000
0!
0%
#725725000000
1!
1%
#725730000000
0!
0%
#725735000000
1!
1%
#725740000000
0!
0%
#725745000000
1!
1%
#725750000000
0!
0%
#725755000000
1!
1%
#725760000000
0!
0%
#725765000000
1!
1%
#725770000000
0!
0%
#725775000000
1!
1%
#725780000000
0!
0%
#725785000000
1!
1%
#725790000000
0!
0%
#725795000000
1!
1%
#725800000000
0!
0%
#725805000000
1!
1%
#725810000000
0!
0%
#725815000000
1!
1%
#725820000000
0!
0%
#725825000000
1!
1%
#725830000000
0!
0%
#725835000000
1!
1%
#725840000000
0!
0%
#725845000000
1!
1%
#725850000000
0!
0%
#725855000000
1!
1%
#725860000000
0!
0%
#725865000000
1!
1%
#725870000000
0!
0%
#725875000000
1!
1%
#725880000000
0!
0%
#725885000000
1!
1%
#725890000000
0!
0%
#725895000000
1!
1%
#725900000000
0!
0%
#725905000000
1!
1%
#725910000000
0!
0%
#725915000000
1!
1%
#725920000000
0!
0%
#725925000000
1!
1%
#725930000000
0!
0%
#725935000000
1!
1%
#725940000000
0!
0%
#725945000000
1!
1%
#725950000000
0!
0%
#725955000000
1!
1%
#725960000000
0!
0%
#725965000000
1!
1%
#725970000000
0!
0%
#725975000000
1!
1%
#725980000000
0!
0%
#725985000000
1!
1%
#725990000000
0!
0%
#725995000000
1!
1%
#726000000000
0!
0%
#726005000000
1!
1%
#726010000000
0!
0%
#726015000000
1!
1%
#726020000000
0!
0%
#726025000000
1!
1%
#726030000000
0!
0%
#726035000000
1!
1%
#726040000000
0!
0%
#726045000000
1!
1%
#726050000000
0!
0%
#726055000000
1!
1%
#726060000000
0!
0%
#726065000000
1!
1%
#726070000000
0!
0%
#726075000000
1!
1%
#726080000000
0!
0%
#726085000000
1!
1%
#726090000000
0!
0%
#726095000000
1!
1%
#726100000000
0!
0%
#726105000000
1!
1%
#726110000000
0!
0%
#726115000000
1!
1%
#726120000000
0!
0%
#726125000000
1!
1%
#726130000000
0!
0%
#726135000000
1!
1%
#726140000000
0!
0%
#726145000000
1!
1%
#726150000000
0!
0%
#726155000000
1!
1%
#726160000000
0!
0%
#726165000000
1!
1%
#726170000000
0!
0%
#726175000000
1!
1%
#726180000000
0!
0%
#726185000000
1!
1%
#726190000000
0!
0%
#726195000000
1!
1%
#726200000000
0!
0%
#726205000000
1!
1%
#726210000000
0!
0%
#726215000000
1!
1%
#726220000000
0!
0%
#726225000000
1!
1%
#726230000000
0!
0%
#726235000000
1!
1%
#726240000000
0!
0%
#726245000000
1!
1%
#726250000000
0!
0%
#726255000000
1!
1%
#726260000000
0!
0%
#726265000000
1!
1%
#726270000000
0!
0%
#726275000000
1!
1%
#726280000000
0!
0%
#726285000000
1!
1%
#726290000000
0!
0%
#726295000000
1!
1%
#726300000000
0!
0%
#726305000000
1!
1%
#726310000000
0!
0%
#726315000000
1!
1%
#726320000000
0!
0%
#726325000000
1!
1%
#726330000000
0!
0%
#726335000000
1!
1%
#726340000000
0!
0%
#726345000000
1!
1%
#726350000000
0!
0%
#726355000000
1!
1%
#726360000000
0!
0%
#726365000000
1!
1%
#726370000000
0!
0%
#726375000000
1!
1%
#726380000000
0!
0%
#726385000000
1!
1%
#726390000000
0!
0%
#726395000000
1!
1%
#726400000000
0!
0%
#726405000000
1!
1%
#726410000000
0!
0%
#726415000000
1!
1%
#726420000000
0!
0%
#726425000000
1!
1%
#726430000000
0!
0%
#726435000000
1!
1%
#726440000000
0!
0%
#726445000000
1!
1%
#726450000000
0!
0%
#726455000000
1!
1%
#726460000000
0!
0%
#726465000000
1!
1%
#726470000000
0!
0%
#726475000000
1!
1%
#726480000000
0!
0%
#726485000000
1!
1%
#726490000000
0!
0%
#726495000000
1!
1%
#726500000000
0!
0%
#726505000000
1!
1%
#726510000000
0!
0%
#726515000000
1!
1%
#726520000000
0!
0%
#726525000000
1!
1%
#726530000000
0!
0%
#726535000000
1!
1%
#726540000000
0!
0%
#726545000000
1!
1%
#726550000000
0!
0%
#726555000000
1!
1%
#726560000000
0!
0%
#726565000000
1!
1%
#726570000000
0!
0%
#726575000000
1!
1%
#726580000000
0!
0%
#726585000000
1!
1%
#726590000000
0!
0%
#726595000000
1!
1%
#726600000000
0!
0%
#726605000000
1!
1%
#726610000000
0!
0%
#726615000000
1!
1%
#726620000000
0!
0%
#726625000000
1!
1%
#726630000000
0!
0%
#726635000000
1!
1%
#726640000000
0!
0%
#726645000000
1!
1%
#726650000000
0!
0%
#726655000000
1!
1%
#726660000000
0!
0%
#726665000000
1!
1%
#726670000000
0!
0%
#726675000000
1!
1%
#726680000000
0!
0%
#726685000000
1!
1%
#726690000000
0!
0%
#726695000000
1!
1%
#726700000000
0!
0%
#726705000000
1!
1%
#726710000000
0!
0%
#726715000000
1!
1%
#726720000000
0!
0%
#726725000000
1!
1%
#726730000000
0!
0%
#726735000000
1!
1%
#726740000000
0!
0%
#726745000000
1!
1%
#726750000000
0!
0%
#726755000000
1!
1%
#726760000000
0!
0%
#726765000000
1!
1%
#726770000000
0!
0%
#726775000000
1!
1%
#726780000000
0!
0%
#726785000000
1!
1%
#726790000000
0!
0%
#726795000000
1!
1%
#726800000000
0!
0%
#726805000000
1!
1%
#726810000000
0!
0%
#726815000000
1!
1%
#726820000000
0!
0%
#726825000000
1!
1%
#726830000000
0!
0%
#726835000000
1!
1%
#726840000000
0!
0%
#726845000000
1!
1%
#726850000000
0!
0%
#726855000000
1!
1%
#726860000000
0!
0%
#726865000000
1!
1%
#726870000000
0!
0%
#726875000000
1!
1%
#726880000000
0!
0%
#726885000000
1!
1%
#726890000000
0!
0%
#726895000000
1!
1%
#726900000000
0!
0%
#726905000000
1!
1%
#726910000000
0!
0%
#726915000000
1!
1%
#726920000000
0!
0%
#726925000000
1!
1%
#726930000000
0!
0%
#726935000000
1!
1%
#726940000000
0!
0%
#726945000000
1!
1%
#726950000000
0!
0%
#726955000000
1!
1%
#726960000000
0!
0%
#726965000000
1!
1%
#726970000000
0!
0%
#726975000000
1!
1%
#726980000000
0!
0%
#726985000000
1!
1%
#726990000000
0!
0%
#726995000000
1!
1%
#727000000000
0!
0%
#727005000000
1!
1%
#727010000000
0!
0%
#727015000000
1!
1%
#727020000000
0!
0%
#727025000000
1!
1%
#727030000000
0!
0%
#727035000000
1!
1%
#727040000000
0!
0%
#727045000000
1!
1%
#727050000000
0!
0%
#727055000000
1!
1%
#727060000000
0!
0%
#727065000000
1!
1%
#727070000000
0!
0%
#727075000000
1!
1%
#727080000000
0!
0%
#727085000000
1!
1%
#727090000000
0!
0%
#727095000000
1!
1%
#727100000000
0!
0%
#727105000000
1!
1%
#727110000000
0!
0%
#727115000000
1!
1%
#727120000000
0!
0%
#727125000000
1!
1%
#727130000000
0!
0%
#727135000000
1!
1%
#727140000000
0!
0%
#727145000000
1!
1%
#727150000000
0!
0%
#727155000000
1!
1%
#727160000000
0!
0%
#727165000000
1!
1%
#727170000000
0!
0%
#727175000000
1!
1%
#727180000000
0!
0%
#727185000000
1!
1%
#727190000000
0!
0%
#727195000000
1!
1%
#727200000000
0!
0%
#727205000000
1!
1%
#727210000000
0!
0%
#727215000000
1!
1%
#727220000000
0!
0%
#727225000000
1!
1%
#727230000000
0!
0%
#727235000000
1!
1%
#727240000000
0!
0%
#727245000000
1!
1%
#727250000000
0!
0%
#727255000000
1!
1%
#727260000000
0!
0%
#727265000000
1!
1%
#727270000000
0!
0%
#727275000000
1!
1%
#727280000000
0!
0%
#727285000000
1!
1%
#727290000000
0!
0%
#727295000000
1!
1%
#727300000000
0!
0%
#727305000000
1!
1%
#727310000000
0!
0%
#727315000000
1!
1%
#727320000000
0!
0%
#727325000000
1!
1%
#727330000000
0!
0%
#727335000000
1!
1%
#727340000000
0!
0%
#727345000000
1!
1%
#727350000000
0!
0%
#727355000000
1!
1%
#727360000000
0!
0%
#727365000000
1!
1%
#727370000000
0!
0%
#727375000000
1!
1%
#727380000000
0!
0%
#727385000000
1!
1%
#727390000000
0!
0%
#727395000000
1!
1%
#727400000000
0!
0%
#727405000000
1!
1%
#727410000000
0!
0%
#727415000000
1!
1%
#727420000000
0!
0%
#727425000000
1!
1%
#727430000000
0!
0%
#727435000000
1!
1%
#727440000000
0!
0%
#727445000000
1!
1%
#727450000000
0!
0%
#727455000000
1!
1%
#727460000000
0!
0%
#727465000000
1!
1%
#727470000000
0!
0%
#727475000000
1!
1%
#727480000000
0!
0%
#727485000000
1!
1%
#727490000000
0!
0%
#727495000000
1!
1%
#727500000000
0!
0%
#727505000000
1!
1%
#727510000000
0!
0%
#727515000000
1!
1%
#727520000000
0!
0%
#727525000000
1!
1%
#727530000000
0!
0%
#727535000000
1!
1%
#727540000000
0!
0%
#727545000000
1!
1%
#727550000000
0!
0%
#727555000000
1!
1%
#727560000000
0!
0%
#727565000000
1!
1%
#727570000000
0!
0%
#727575000000
1!
1%
#727580000000
0!
0%
#727585000000
1!
1%
#727590000000
0!
0%
#727595000000
1!
1%
#727600000000
0!
0%
#727605000000
1!
1%
#727610000000
0!
0%
#727615000000
1!
1%
#727620000000
0!
0%
#727625000000
1!
1%
#727630000000
0!
0%
#727635000000
1!
1%
#727640000000
0!
0%
#727645000000
1!
1%
#727650000000
0!
0%
#727655000000
1!
1%
#727660000000
0!
0%
#727665000000
1!
1%
#727670000000
0!
0%
#727675000000
1!
1%
#727680000000
0!
0%
#727685000000
1!
1%
#727690000000
0!
0%
#727695000000
1!
1%
#727700000000
0!
0%
#727705000000
1!
1%
#727710000000
0!
0%
#727715000000
1!
1%
#727720000000
0!
0%
#727725000000
1!
1%
#727730000000
0!
0%
#727735000000
1!
1%
#727740000000
0!
0%
#727745000000
1!
1%
#727750000000
0!
0%
#727755000000
1!
1%
#727760000000
0!
0%
#727765000000
1!
1%
#727770000000
0!
0%
#727775000000
1!
1%
#727780000000
0!
0%
#727785000000
1!
1%
#727790000000
0!
0%
#727795000000
1!
1%
#727800000000
0!
0%
#727805000000
1!
1%
#727810000000
0!
0%
#727815000000
1!
1%
#727820000000
0!
0%
#727825000000
1!
1%
#727830000000
0!
0%
#727835000000
1!
1%
#727840000000
0!
0%
#727845000000
1!
1%
#727850000000
0!
0%
#727855000000
1!
1%
#727860000000
0!
0%
#727865000000
1!
1%
#727870000000
0!
0%
#727875000000
1!
1%
#727880000000
0!
0%
#727885000000
1!
1%
#727890000000
0!
0%
#727895000000
1!
1%
#727900000000
0!
0%
#727905000000
1!
1%
#727910000000
0!
0%
#727915000000
1!
1%
#727920000000
0!
0%
#727925000000
1!
1%
#727930000000
0!
0%
#727935000000
1!
1%
#727940000000
0!
0%
#727945000000
1!
1%
#727950000000
0!
0%
#727955000000
1!
1%
#727960000000
0!
0%
#727965000000
1!
1%
#727970000000
0!
0%
#727975000000
1!
1%
#727980000000
0!
0%
#727985000000
1!
1%
#727990000000
0!
0%
#727995000000
1!
1%
#728000000000
0!
0%
#728005000000
1!
1%
#728010000000
0!
0%
#728015000000
1!
1%
#728020000000
0!
0%
#728025000000
1!
1%
#728030000000
0!
0%
#728035000000
1!
1%
#728040000000
0!
0%
#728045000000
1!
1%
#728050000000
0!
0%
#728055000000
1!
1%
#728060000000
0!
0%
#728065000000
1!
1%
#728070000000
0!
0%
#728075000000
1!
1%
#728080000000
0!
0%
#728085000000
1!
1%
#728090000000
0!
0%
#728095000000
1!
1%
#728100000000
0!
0%
#728105000000
1!
1%
#728110000000
0!
0%
#728115000000
1!
1%
#728120000000
0!
0%
#728125000000
1!
1%
#728130000000
0!
0%
#728135000000
1!
1%
#728140000000
0!
0%
#728145000000
1!
1%
#728150000000
0!
0%
#728155000000
1!
1%
#728160000000
0!
0%
#728165000000
1!
1%
#728170000000
0!
0%
#728175000000
1!
1%
#728180000000
0!
0%
#728185000000
1!
1%
#728190000000
0!
0%
#728195000000
1!
1%
#728200000000
0!
0%
#728205000000
1!
1%
#728210000000
0!
0%
#728215000000
1!
1%
#728220000000
0!
0%
#728225000000
1!
1%
#728230000000
0!
0%
#728235000000
1!
1%
#728240000000
0!
0%
#728245000000
1!
1%
#728250000000
0!
0%
#728255000000
1!
1%
#728260000000
0!
0%
#728265000000
1!
1%
#728270000000
0!
0%
#728275000000
1!
1%
#728280000000
0!
0%
#728285000000
1!
1%
#728290000000
0!
0%
#728295000000
1!
1%
#728300000000
0!
0%
#728305000000
1!
1%
#728310000000
0!
0%
#728315000000
1!
1%
#728320000000
0!
0%
#728325000000
1!
1%
#728330000000
0!
0%
#728335000000
1!
1%
#728340000000
0!
0%
#728345000000
1!
1%
#728350000000
0!
0%
#728355000000
1!
1%
#728360000000
0!
0%
#728365000000
1!
1%
#728370000000
0!
0%
#728375000000
1!
1%
#728380000000
0!
0%
#728385000000
1!
1%
#728390000000
0!
0%
#728395000000
1!
1%
#728400000000
0!
0%
#728405000000
1!
1%
#728410000000
0!
0%
#728415000000
1!
1%
#728420000000
0!
0%
#728425000000
1!
1%
#728430000000
0!
0%
#728435000000
1!
1%
#728440000000
0!
0%
#728445000000
1!
1%
#728450000000
0!
0%
#728455000000
1!
1%
#728460000000
0!
0%
#728465000000
1!
1%
#728470000000
0!
0%
#728475000000
1!
1%
#728480000000
0!
0%
#728485000000
1!
1%
#728490000000
0!
0%
#728495000000
1!
1%
#728500000000
0!
0%
#728505000000
1!
1%
#728510000000
0!
0%
#728515000000
1!
1%
#728520000000
0!
0%
#728525000000
1!
1%
#728530000000
0!
0%
#728535000000
1!
1%
#728540000000
0!
0%
#728545000000
1!
1%
#728550000000
0!
0%
#728555000000
1!
1%
#728560000000
0!
0%
#728565000000
1!
1%
#728570000000
0!
0%
#728575000000
1!
1%
#728580000000
0!
0%
#728585000000
1!
1%
#728590000000
0!
0%
#728595000000
1!
1%
#728600000000
0!
0%
#728605000000
1!
1%
#728610000000
0!
0%
#728615000000
1!
1%
#728620000000
0!
0%
#728625000000
1!
1%
#728630000000
0!
0%
#728635000000
1!
1%
#728640000000
0!
0%
#728645000000
1!
1%
#728650000000
0!
0%
#728655000000
1!
1%
#728660000000
0!
0%
#728665000000
1!
1%
#728670000000
0!
0%
#728675000000
1!
1%
#728680000000
0!
0%
#728685000000
1!
1%
#728690000000
0!
0%
#728695000000
1!
1%
#728700000000
0!
0%
#728705000000
1!
1%
#728710000000
0!
0%
#728715000000
1!
1%
#728720000000
0!
0%
#728725000000
1!
1%
#728730000000
0!
0%
#728735000000
1!
1%
#728740000000
0!
0%
#728745000000
1!
1%
#728750000000
0!
0%
#728755000000
1!
1%
#728760000000
0!
0%
#728765000000
1!
1%
#728770000000
0!
0%
#728775000000
1!
1%
#728780000000
0!
0%
#728785000000
1!
1%
#728790000000
0!
0%
#728795000000
1!
1%
#728800000000
0!
0%
#728805000000
1!
1%
#728810000000
0!
0%
#728815000000
1!
1%
#728820000000
0!
0%
#728825000000
1!
1%
#728830000000
0!
0%
#728835000000
1!
1%
#728840000000
0!
0%
#728845000000
1!
1%
#728850000000
0!
0%
#728855000000
1!
1%
#728860000000
0!
0%
#728865000000
1!
1%
#728870000000
0!
0%
#728875000000
1!
1%
#728880000000
0!
0%
#728885000000
1!
1%
#728890000000
0!
0%
#728895000000
1!
1%
#728900000000
0!
0%
#728905000000
1!
1%
#728910000000
0!
0%
#728915000000
1!
1%
#728920000000
0!
0%
#728925000000
1!
1%
#728930000000
0!
0%
#728935000000
1!
1%
#728940000000
0!
0%
#728945000000
1!
1%
#728950000000
0!
0%
#728955000000
1!
1%
#728960000000
0!
0%
#728965000000
1!
1%
#728970000000
0!
0%
#728975000000
1!
1%
#728980000000
0!
0%
#728985000000
1!
1%
#728990000000
0!
0%
#728995000000
1!
1%
#729000000000
0!
0%
#729005000000
1!
1%
#729010000000
0!
0%
#729015000000
1!
1%
#729020000000
0!
0%
#729025000000
1!
1%
#729030000000
0!
0%
#729035000000
1!
1%
#729040000000
0!
0%
#729045000000
1!
1%
#729050000000
0!
0%
#729055000000
1!
1%
#729060000000
0!
0%
#729065000000
1!
1%
#729070000000
0!
0%
#729075000000
1!
1%
#729080000000
0!
0%
#729085000000
1!
1%
#729090000000
0!
0%
#729095000000
1!
1%
#729100000000
0!
0%
#729105000000
1!
1%
#729110000000
0!
0%
#729115000000
1!
1%
#729120000000
0!
0%
#729125000000
1!
1%
#729130000000
0!
0%
#729135000000
1!
1%
#729140000000
0!
0%
#729145000000
1!
1%
#729150000000
0!
0%
#729155000000
1!
1%
#729160000000
0!
0%
#729165000000
1!
1%
#729170000000
0!
0%
#729175000000
1!
1%
#729180000000
0!
0%
#729185000000
1!
1%
#729190000000
0!
0%
#729195000000
1!
1%
#729200000000
0!
0%
#729205000000
1!
1%
#729210000000
0!
0%
#729215000000
1!
1%
#729220000000
0!
0%
#729225000000
1!
1%
#729230000000
0!
0%
#729235000000
1!
1%
#729240000000
0!
0%
#729245000000
1!
1%
#729250000000
0!
0%
#729255000000
1!
1%
#729260000000
0!
0%
#729265000000
1!
1%
#729270000000
0!
0%
#729275000000
1!
1%
#729280000000
0!
0%
#729285000000
1!
1%
#729290000000
0!
0%
#729295000000
1!
1%
#729300000000
0!
0%
#729305000000
1!
1%
#729310000000
0!
0%
#729315000000
1!
1%
#729320000000
0!
0%
#729325000000
1!
1%
#729330000000
0!
0%
#729335000000
1!
1%
#729340000000
0!
0%
#729345000000
1!
1%
#729350000000
0!
0%
#729355000000
1!
1%
#729360000000
0!
0%
#729365000000
1!
1%
#729370000000
0!
0%
#729375000000
1!
1%
#729380000000
0!
0%
#729385000000
1!
1%
#729390000000
0!
0%
#729395000000
1!
1%
#729400000000
0!
0%
#729405000000
1!
1%
#729410000000
0!
0%
#729415000000
1!
1%
#729420000000
0!
0%
#729425000000
1!
1%
#729430000000
0!
0%
#729435000000
1!
1%
#729440000000
0!
0%
#729445000000
1!
1%
#729450000000
0!
0%
#729455000000
1!
1%
#729460000000
0!
0%
#729465000000
1!
1%
#729470000000
0!
0%
#729475000000
1!
1%
#729480000000
0!
0%
#729485000000
1!
1%
#729490000000
0!
0%
#729495000000
1!
1%
#729500000000
0!
0%
#729505000000
1!
1%
#729510000000
0!
0%
#729515000000
1!
1%
#729520000000
0!
0%
#729525000000
1!
1%
#729530000000
0!
0%
#729535000000
1!
1%
#729540000000
0!
0%
#729545000000
1!
1%
#729550000000
0!
0%
#729555000000
1!
1%
#729560000000
0!
0%
#729565000000
1!
1%
#729570000000
0!
0%
#729575000000
1!
1%
#729580000000
0!
0%
#729585000000
1!
1%
#729590000000
0!
0%
#729595000000
1!
1%
#729600000000
0!
0%
#729605000000
1!
1%
#729610000000
0!
0%
#729615000000
1!
1%
#729620000000
0!
0%
#729625000000
1!
1%
#729630000000
0!
0%
#729635000000
1!
1%
#729640000000
0!
0%
#729645000000
1!
1%
#729650000000
0!
0%
#729655000000
1!
1%
#729660000000
0!
0%
#729665000000
1!
1%
#729670000000
0!
0%
#729675000000
1!
1%
#729680000000
0!
0%
#729685000000
1!
1%
#729690000000
0!
0%
#729695000000
1!
1%
#729700000000
0!
0%
#729705000000
1!
1%
#729710000000
0!
0%
#729715000000
1!
1%
#729720000000
0!
0%
#729725000000
1!
1%
#729730000000
0!
0%
#729735000000
1!
1%
#729740000000
0!
0%
#729745000000
1!
1%
#729750000000
0!
0%
#729755000000
1!
1%
#729760000000
0!
0%
#729765000000
1!
1%
#729770000000
0!
0%
#729775000000
1!
1%
#729780000000
0!
0%
#729785000000
1!
1%
#729790000000
0!
0%
#729795000000
1!
1%
#729800000000
0!
0%
#729805000000
1!
1%
#729810000000
0!
0%
#729815000000
1!
1%
#729820000000
0!
0%
#729825000000
1!
1%
#729830000000
0!
0%
#729835000000
1!
1%
#729840000000
0!
0%
#729845000000
1!
1%
#729850000000
0!
0%
#729855000000
1!
1%
#729860000000
0!
0%
#729865000000
1!
1%
#729870000000
0!
0%
#729875000000
1!
1%
#729880000000
0!
0%
#729885000000
1!
1%
#729890000000
0!
0%
#729895000000
1!
1%
#729900000000
0!
0%
#729905000000
1!
1%
#729910000000
0!
0%
#729915000000
1!
1%
#729920000000
0!
0%
#729925000000
1!
1%
#729930000000
0!
0%
#729935000000
1!
1%
#729940000000
0!
0%
#729945000000
1!
1%
#729950000000
0!
0%
#729955000000
1!
1%
#729960000000
0!
0%
#729965000000
1!
1%
#729970000000
0!
0%
#729975000000
1!
1%
#729980000000
0!
0%
#729985000000
1!
1%
#729990000000
0!
0%
#729995000000
1!
1%
#730000000000
0!
0%
#730005000000
1!
1%
#730010000000
0!
0%
#730015000000
1!
1%
#730020000000
0!
0%
#730025000000
1!
1%
#730030000000
0!
0%
#730035000000
1!
1%
#730040000000
0!
0%
#730045000000
1!
1%
#730050000000
0!
0%
#730055000000
1!
1%
#730060000000
0!
0%
#730065000000
1!
1%
#730070000000
0!
0%
#730075000000
1!
1%
#730080000000
0!
0%
#730085000000
1!
1%
#730090000000
0!
0%
#730095000000
1!
1%
#730100000000
0!
0%
#730105000000
1!
1%
#730110000000
0!
0%
#730115000000
1!
1%
#730120000000
0!
0%
#730125000000
1!
1%
#730130000000
0!
0%
#730135000000
1!
1%
#730140000000
0!
0%
#730145000000
1!
1%
#730150000000
0!
0%
#730155000000
1!
1%
#730160000000
0!
0%
#730165000000
1!
1%
#730170000000
0!
0%
#730175000000
1!
1%
#730180000000
0!
0%
#730185000000
1!
1%
#730190000000
0!
0%
#730195000000
1!
1%
#730200000000
0!
0%
#730205000000
1!
1%
#730210000000
0!
0%
#730215000000
1!
1%
#730220000000
0!
0%
#730225000000
1!
1%
#730230000000
0!
0%
#730235000000
1!
1%
#730240000000
0!
0%
#730245000000
1!
1%
#730250000000
0!
0%
#730255000000
1!
1%
#730260000000
0!
0%
#730265000000
1!
1%
#730270000000
0!
0%
#730275000000
1!
1%
#730280000000
0!
0%
#730285000000
1!
1%
#730290000000
0!
0%
#730295000000
1!
1%
#730300000000
0!
0%
#730305000000
1!
1%
#730310000000
0!
0%
#730315000000
1!
1%
#730320000000
0!
0%
#730325000000
1!
1%
#730330000000
0!
0%
#730335000000
1!
1%
#730340000000
0!
0%
#730345000000
1!
1%
#730350000000
0!
0%
#730355000000
1!
1%
#730360000000
0!
0%
#730365000000
1!
1%
#730370000000
0!
0%
#730375000000
1!
1%
#730380000000
0!
0%
#730385000000
1!
1%
#730390000000
0!
0%
#730395000000
1!
1%
#730400000000
0!
0%
#730405000000
1!
1%
#730410000000
0!
0%
#730415000000
1!
1%
#730420000000
0!
0%
#730425000000
1!
1%
#730430000000
0!
0%
#730435000000
1!
1%
#730440000000
0!
0%
#730445000000
1!
1%
#730450000000
0!
0%
#730455000000
1!
1%
#730460000000
0!
0%
#730465000000
1!
1%
#730470000000
0!
0%
#730475000000
1!
1%
#730480000000
0!
0%
#730485000000
1!
1%
#730490000000
0!
0%
#730495000000
1!
1%
#730500000000
0!
0%
#730505000000
1!
1%
#730510000000
0!
0%
#730515000000
1!
1%
#730520000000
0!
0%
#730525000000
1!
1%
#730530000000
0!
0%
#730535000000
1!
1%
#730540000000
0!
0%
#730545000000
1!
1%
#730550000000
0!
0%
#730555000000
1!
1%
#730560000000
0!
0%
#730565000000
1!
1%
#730570000000
0!
0%
#730575000000
1!
1%
#730580000000
0!
0%
#730585000000
1!
1%
#730590000000
0!
0%
#730595000000
1!
1%
#730600000000
0!
0%
#730605000000
1!
1%
#730610000000
0!
0%
#730615000000
1!
1%
#730620000000
0!
0%
#730625000000
1!
1%
#730630000000
0!
0%
#730635000000
1!
1%
#730640000000
0!
0%
#730645000000
1!
1%
#730650000000
0!
0%
#730655000000
1!
1%
#730660000000
0!
0%
#730665000000
1!
1%
#730670000000
0!
0%
#730675000000
1!
1%
#730680000000
0!
0%
#730685000000
1!
1%
#730690000000
0!
0%
#730695000000
1!
1%
#730700000000
0!
0%
#730705000000
1!
1%
#730710000000
0!
0%
#730715000000
1!
1%
#730720000000
0!
0%
#730725000000
1!
1%
#730730000000
0!
0%
#730735000000
1!
1%
#730740000000
0!
0%
#730745000000
1!
1%
#730750000000
0!
0%
#730755000000
1!
1%
#730760000000
0!
0%
#730765000000
1!
1%
#730770000000
0!
0%
#730775000000
1!
1%
#730780000000
0!
0%
#730785000000
1!
1%
#730790000000
0!
0%
#730795000000
1!
1%
#730800000000
0!
0%
#730805000000
1!
1%
#730810000000
0!
0%
#730815000000
1!
1%
#730820000000
0!
0%
#730825000000
1!
1%
#730830000000
0!
0%
#730835000000
1!
1%
#730840000000
0!
0%
#730845000000
1!
1%
#730850000000
0!
0%
#730855000000
1!
1%
#730860000000
0!
0%
#730865000000
1!
1%
#730870000000
0!
0%
#730875000000
1!
1%
#730880000000
0!
0%
#730885000000
1!
1%
#730890000000
0!
0%
#730895000000
1!
1%
#730900000000
0!
0%
#730905000000
1!
1%
#730910000000
0!
0%
#730915000000
1!
1%
#730920000000
0!
0%
#730925000000
1!
1%
#730930000000
0!
0%
#730935000000
1!
1%
#730940000000
0!
0%
#730945000000
1!
1%
#730950000000
0!
0%
#730955000000
1!
1%
#730960000000
0!
0%
#730965000000
1!
1%
#730970000000
0!
0%
#730975000000
1!
1%
#730980000000
0!
0%
#730985000000
1!
1%
#730990000000
0!
0%
#730995000000
1!
1%
#731000000000
0!
0%
#731005000000
1!
1%
#731010000000
0!
0%
#731015000000
1!
1%
#731020000000
0!
0%
#731025000000
1!
1%
#731030000000
0!
0%
#731035000000
1!
1%
#731040000000
0!
0%
#731045000000
1!
1%
#731050000000
0!
0%
#731055000000
1!
1%
#731060000000
0!
0%
#731065000000
1!
1%
#731070000000
0!
0%
#731075000000
1!
1%
#731080000000
0!
0%
#731085000000
1!
1%
#731090000000
0!
0%
#731095000000
1!
1%
#731100000000
0!
0%
#731105000000
1!
1%
#731110000000
0!
0%
#731115000000
1!
1%
#731120000000
0!
0%
#731125000000
1!
1%
#731130000000
0!
0%
#731135000000
1!
1%
#731140000000
0!
0%
#731145000000
1!
1%
#731150000000
0!
0%
#731155000000
1!
1%
#731160000000
0!
0%
#731165000000
1!
1%
#731170000000
0!
0%
#731175000000
1!
1%
#731180000000
0!
0%
#731185000000
1!
1%
#731190000000
0!
0%
#731195000000
1!
1%
#731200000000
0!
0%
#731205000000
1!
1%
#731210000000
0!
0%
#731215000000
1!
1%
#731220000000
0!
0%
#731225000000
1!
1%
#731230000000
0!
0%
#731235000000
1!
1%
#731240000000
0!
0%
#731245000000
1!
1%
#731250000000
0!
0%
#731255000000
1!
1%
#731260000000
0!
0%
#731265000000
1!
1%
#731270000000
0!
0%
#731275000000
1!
1%
#731280000000
0!
0%
#731285000000
1!
1%
#731290000000
0!
0%
#731295000000
1!
1%
#731300000000
0!
0%
#731305000000
1!
1%
#731310000000
0!
0%
#731315000000
1!
1%
#731320000000
0!
0%
#731325000000
1!
1%
#731330000000
0!
0%
#731335000000
1!
1%
#731340000000
0!
0%
#731345000000
1!
1%
#731350000000
0!
0%
#731355000000
1!
1%
#731360000000
0!
0%
#731365000000
1!
1%
#731370000000
0!
0%
#731375000000
1!
1%
#731380000000
0!
0%
#731385000000
1!
1%
#731390000000
0!
0%
#731395000000
1!
1%
#731400000000
0!
0%
#731405000000
1!
1%
#731410000000
0!
0%
#731415000000
1!
1%
#731420000000
0!
0%
#731425000000
1!
1%
#731430000000
0!
0%
#731435000000
1!
1%
#731440000000
0!
0%
#731445000000
1!
1%
#731450000000
0!
0%
#731455000000
1!
1%
#731460000000
0!
0%
#731465000000
1!
1%
#731470000000
0!
0%
#731475000000
1!
1%
#731480000000
0!
0%
#731485000000
1!
1%
#731490000000
0!
0%
#731495000000
1!
1%
#731500000000
0!
0%
#731505000000
1!
1%
#731510000000
0!
0%
#731515000000
1!
1%
#731520000000
0!
0%
#731525000000
1!
1%
#731530000000
0!
0%
#731535000000
1!
1%
#731540000000
0!
0%
#731545000000
1!
1%
#731550000000
0!
0%
#731555000000
1!
1%
#731560000000
0!
0%
#731565000000
1!
1%
#731570000000
0!
0%
#731575000000
1!
1%
#731580000000
0!
0%
#731585000000
1!
1%
#731590000000
0!
0%
#731595000000
1!
1%
#731600000000
0!
0%
#731605000000
1!
1%
#731610000000
0!
0%
#731615000000
1!
1%
#731620000000
0!
0%
#731625000000
1!
1%
#731630000000
0!
0%
#731635000000
1!
1%
#731640000000
0!
0%
#731645000000
1!
1%
#731650000000
0!
0%
#731655000000
1!
1%
#731660000000
0!
0%
#731665000000
1!
1%
#731670000000
0!
0%
#731675000000
1!
1%
#731680000000
0!
0%
#731685000000
1!
1%
#731690000000
0!
0%
#731695000000
1!
1%
#731700000000
0!
0%
#731705000000
1!
1%
#731710000000
0!
0%
#731715000000
1!
1%
#731720000000
0!
0%
#731725000000
1!
1%
#731730000000
0!
0%
#731735000000
1!
1%
#731740000000
0!
0%
#731745000000
1!
1%
#731750000000
0!
0%
#731755000000
1!
1%
#731760000000
0!
0%
#731765000000
1!
1%
#731770000000
0!
0%
#731775000000
1!
1%
#731780000000
0!
0%
#731785000000
1!
1%
#731790000000
0!
0%
#731795000000
1!
1%
#731800000000
0!
0%
#731805000000
1!
1%
#731810000000
0!
0%
#731815000000
1!
1%
#731820000000
0!
0%
#731825000000
1!
1%
#731830000000
0!
0%
#731835000000
1!
1%
#731840000000
0!
0%
#731845000000
1!
1%
#731850000000
0!
0%
#731855000000
1!
1%
#731860000000
0!
0%
#731865000000
1!
1%
#731870000000
0!
0%
#731875000000
1!
1%
#731880000000
0!
0%
#731885000000
1!
1%
#731890000000
0!
0%
#731895000000
1!
1%
#731900000000
0!
0%
#731905000000
1!
1%
#731910000000
0!
0%
#731915000000
1!
1%
#731920000000
0!
0%
#731925000000
1!
1%
#731930000000
0!
0%
#731935000000
1!
1%
#731940000000
0!
0%
#731945000000
1!
1%
#731950000000
0!
0%
#731955000000
1!
1%
#731960000000
0!
0%
#731965000000
1!
1%
#731970000000
0!
0%
#731975000000
1!
1%
#731980000000
0!
0%
#731985000000
1!
1%
#731990000000
0!
0%
#731995000000
1!
1%
#732000000000
0!
0%
#732005000000
1!
1%
#732010000000
0!
0%
#732015000000
1!
1%
#732020000000
0!
0%
#732025000000
1!
1%
#732030000000
0!
0%
#732035000000
1!
1%
#732040000000
0!
0%
#732045000000
1!
1%
#732050000000
0!
0%
#732055000000
1!
1%
#732060000000
0!
0%
#732065000000
1!
1%
#732070000000
0!
0%
#732075000000
1!
1%
#732080000000
0!
0%
#732085000000
1!
1%
#732090000000
0!
0%
#732095000000
1!
1%
#732100000000
0!
0%
#732105000000
1!
1%
#732110000000
0!
0%
#732115000000
1!
1%
#732120000000
0!
0%
#732125000000
1!
1%
#732130000000
0!
0%
#732135000000
1!
1%
#732140000000
0!
0%
#732145000000
1!
1%
#732150000000
0!
0%
#732155000000
1!
1%
#732160000000
0!
0%
#732165000000
1!
1%
#732170000000
0!
0%
#732175000000
1!
1%
#732180000000
0!
0%
#732185000000
1!
1%
#732190000000
0!
0%
#732195000000
1!
1%
#732200000000
0!
0%
#732205000000
1!
1%
#732210000000
0!
0%
#732215000000
1!
1%
#732220000000
0!
0%
#732225000000
1!
1%
#732230000000
0!
0%
#732235000000
1!
1%
#732240000000
0!
0%
#732245000000
1!
1%
#732250000000
0!
0%
#732255000000
1!
1%
#732260000000
0!
0%
#732265000000
1!
1%
#732270000000
0!
0%
#732275000000
1!
1%
#732280000000
0!
0%
#732285000000
1!
1%
#732290000000
0!
0%
#732295000000
1!
1%
#732300000000
0!
0%
#732305000000
1!
1%
#732310000000
0!
0%
#732315000000
1!
1%
#732320000000
0!
0%
#732325000000
1!
1%
#732330000000
0!
0%
#732335000000
1!
1%
#732340000000
0!
0%
#732345000000
1!
1%
#732350000000
0!
0%
#732355000000
1!
1%
#732360000000
0!
0%
#732365000000
1!
1%
#732370000000
0!
0%
#732375000000
1!
1%
#732380000000
0!
0%
#732385000000
1!
1%
#732390000000
0!
0%
#732395000000
1!
1%
#732400000000
0!
0%
#732405000000
1!
1%
#732410000000
0!
0%
#732415000000
1!
1%
#732420000000
0!
0%
#732425000000
1!
1%
#732430000000
0!
0%
#732435000000
1!
1%
#732440000000
0!
0%
#732445000000
1!
1%
#732450000000
0!
0%
#732455000000
1!
1%
#732460000000
0!
0%
#732465000000
1!
1%
#732470000000
0!
0%
#732475000000
1!
1%
#732480000000
0!
0%
#732485000000
1!
1%
#732490000000
0!
0%
#732495000000
1!
1%
#732500000000
0!
0%
#732505000000
1!
1%
#732510000000
0!
0%
#732515000000
1!
1%
#732520000000
0!
0%
#732525000000
1!
1%
#732530000000
0!
0%
#732535000000
1!
1%
#732540000000
0!
0%
#732545000000
1!
1%
#732550000000
0!
0%
#732555000000
1!
1%
#732560000000
0!
0%
#732565000000
1!
1%
#732570000000
0!
0%
#732575000000
1!
1%
#732580000000
0!
0%
#732585000000
1!
1%
#732590000000
0!
0%
#732595000000
1!
1%
#732600000000
0!
0%
#732605000000
1!
1%
#732610000000
0!
0%
#732615000000
1!
1%
#732620000000
0!
0%
#732625000000
1!
1%
#732630000000
0!
0%
#732635000000
1!
1%
#732640000000
0!
0%
#732645000000
1!
1%
#732650000000
0!
0%
#732655000000
1!
1%
#732660000000
0!
0%
#732665000000
1!
1%
#732670000000
0!
0%
#732675000000
1!
1%
#732680000000
0!
0%
#732685000000
1!
1%
#732690000000
0!
0%
#732695000000
1!
1%
#732700000000
0!
0%
#732705000000
1!
1%
#732710000000
0!
0%
#732715000000
1!
1%
#732720000000
0!
0%
#732725000000
1!
1%
#732730000000
0!
0%
#732735000000
1!
1%
#732740000000
0!
0%
#732745000000
1!
1%
#732750000000
0!
0%
#732755000000
1!
1%
#732760000000
0!
0%
#732765000000
1!
1%
#732770000000
0!
0%
#732775000000
1!
1%
#732780000000
0!
0%
#732785000000
1!
1%
#732790000000
0!
0%
#732795000000
1!
1%
#732800000000
0!
0%
#732805000000
1!
1%
#732810000000
0!
0%
#732815000000
1!
1%
#732820000000
0!
0%
#732825000000
1!
1%
#732830000000
0!
0%
#732835000000
1!
1%
#732840000000
0!
0%
#732845000000
1!
1%
#732850000000
0!
0%
#732855000000
1!
1%
#732860000000
0!
0%
#732865000000
1!
1%
#732870000000
0!
0%
#732875000000
1!
1%
#732880000000
0!
0%
#732885000000
1!
1%
#732890000000
0!
0%
#732895000000
1!
1%
#732900000000
0!
0%
#732905000000
1!
1%
#732910000000
0!
0%
#732915000000
1!
1%
#732920000000
0!
0%
#732925000000
1!
1%
#732930000000
0!
0%
#732935000000
1!
1%
#732940000000
0!
0%
#732945000000
1!
1%
#732950000000
0!
0%
#732955000000
1!
1%
#732960000000
0!
0%
#732965000000
1!
1%
#732970000000
0!
0%
#732975000000
1!
1%
#732980000000
0!
0%
#732985000000
1!
1%
#732990000000
0!
0%
#732995000000
1!
1%
#733000000000
0!
0%
#733005000000
1!
1%
#733010000000
0!
0%
#733015000000
1!
1%
#733020000000
0!
0%
#733025000000
1!
1%
#733030000000
0!
0%
#733035000000
1!
1%
#733040000000
0!
0%
#733045000000
1!
1%
#733050000000
0!
0%
#733055000000
1!
1%
#733060000000
0!
0%
#733065000000
1!
1%
#733070000000
0!
0%
#733075000000
1!
1%
#733080000000
0!
0%
#733085000000
1!
1%
#733090000000
0!
0%
#733095000000
1!
1%
#733100000000
0!
0%
#733105000000
1!
1%
#733110000000
0!
0%
#733115000000
1!
1%
#733120000000
0!
0%
#733125000000
1!
1%
#733130000000
0!
0%
#733135000000
1!
1%
#733140000000
0!
0%
#733145000000
1!
1%
#733150000000
0!
0%
#733155000000
1!
1%
#733160000000
0!
0%
#733165000000
1!
1%
#733170000000
0!
0%
#733175000000
1!
1%
#733180000000
0!
0%
#733185000000
1!
1%
#733190000000
0!
0%
#733195000000
1!
1%
#733200000000
0!
0%
#733205000000
1!
1%
#733210000000
0!
0%
#733215000000
1!
1%
#733220000000
0!
0%
#733225000000
1!
1%
#733230000000
0!
0%
#733235000000
1!
1%
#733240000000
0!
0%
#733245000000
1!
1%
#733250000000
0!
0%
#733255000000
1!
1%
#733260000000
0!
0%
#733265000000
1!
1%
#733270000000
0!
0%
#733275000000
1!
1%
#733280000000
0!
0%
#733285000000
1!
1%
#733290000000
0!
0%
#733295000000
1!
1%
#733300000000
0!
0%
#733305000000
1!
1%
#733310000000
0!
0%
#733315000000
1!
1%
#733320000000
0!
0%
#733325000000
1!
1%
#733330000000
0!
0%
#733335000000
1!
1%
#733340000000
0!
0%
#733345000000
1!
1%
#733350000000
0!
0%
#733355000000
1!
1%
#733360000000
0!
0%
#733365000000
1!
1%
#733370000000
0!
0%
#733375000000
1!
1%
#733380000000
0!
0%
#733385000000
1!
1%
#733390000000
0!
0%
#733395000000
1!
1%
#733400000000
0!
0%
#733405000000
1!
1%
#733410000000
0!
0%
#733415000000
1!
1%
#733420000000
0!
0%
#733425000000
1!
1%
#733430000000
0!
0%
#733435000000
1!
1%
#733440000000
0!
0%
#733445000000
1!
1%
#733450000000
0!
0%
#733455000000
1!
1%
#733460000000
0!
0%
#733465000000
1!
1%
#733470000000
0!
0%
#733475000000
1!
1%
#733480000000
0!
0%
#733485000000
1!
1%
#733490000000
0!
0%
#733495000000
1!
1%
#733500000000
0!
0%
#733505000000
1!
1%
#733510000000
0!
0%
#733515000000
1!
1%
#733520000000
0!
0%
#733525000000
1!
1%
#733530000000
0!
0%
#733535000000
1!
1%
#733540000000
0!
0%
#733545000000
1!
1%
#733550000000
0!
0%
#733555000000
1!
1%
#733560000000
0!
0%
#733565000000
1!
1%
#733570000000
0!
0%
#733575000000
1!
1%
#733580000000
0!
0%
#733585000000
1!
1%
#733590000000
0!
0%
#733595000000
1!
1%
#733600000000
0!
0%
#733605000000
1!
1%
#733610000000
0!
0%
#733615000000
1!
1%
#733620000000
0!
0%
#733625000000
1!
1%
#733630000000
0!
0%
#733635000000
1!
1%
#733640000000
0!
0%
#733645000000
1!
1%
#733650000000
0!
0%
#733655000000
1!
1%
#733660000000
0!
0%
#733665000000
1!
1%
#733670000000
0!
0%
#733675000000
1!
1%
#733680000000
0!
0%
#733685000000
1!
1%
#733690000000
0!
0%
#733695000000
1!
1%
#733700000000
0!
0%
#733705000000
1!
1%
#733710000000
0!
0%
#733715000000
1!
1%
#733720000000
0!
0%
#733725000000
1!
1%
#733730000000
0!
0%
#733735000000
1!
1%
#733740000000
0!
0%
#733745000000
1!
1%
#733750000000
0!
0%
#733755000000
1!
1%
#733760000000
0!
0%
#733765000000
1!
1%
#733770000000
0!
0%
#733775000000
1!
1%
#733780000000
0!
0%
#733785000000
1!
1%
#733790000000
0!
0%
#733795000000
1!
1%
#733800000000
0!
0%
#733805000000
1!
1%
#733810000000
0!
0%
#733815000000
1!
1%
#733820000000
0!
0%
#733825000000
1!
1%
#733830000000
0!
0%
#733835000000
1!
1%
#733840000000
0!
0%
#733845000000
1!
1%
#733850000000
0!
0%
#733855000000
1!
1%
#733860000000
0!
0%
#733865000000
1!
1%
#733870000000
0!
0%
#733875000000
1!
1%
#733880000000
0!
0%
#733885000000
1!
1%
#733890000000
0!
0%
#733895000000
1!
1%
#733900000000
0!
0%
#733905000000
1!
1%
#733910000000
0!
0%
#733915000000
1!
1%
#733920000000
0!
0%
#733925000000
1!
1%
#733930000000
0!
0%
#733935000000
1!
1%
#733940000000
0!
0%
#733945000000
1!
1%
#733950000000
0!
0%
#733955000000
1!
1%
#733960000000
0!
0%
#733965000000
1!
1%
#733970000000
0!
0%
#733975000000
1!
1%
#733980000000
0!
0%
#733985000000
1!
1%
#733990000000
0!
0%
#733995000000
1!
1%
#734000000000
0!
0%
#734005000000
1!
1%
#734010000000
0!
0%
#734015000000
1!
1%
#734020000000
0!
0%
#734025000000
1!
1%
#734030000000
0!
0%
#734035000000
1!
1%
#734040000000
0!
0%
#734045000000
1!
1%
#734050000000
0!
0%
#734055000000
1!
1%
#734060000000
0!
0%
#734065000000
1!
1%
#734070000000
0!
0%
#734075000000
1!
1%
#734080000000
0!
0%
#734085000000
1!
1%
#734090000000
0!
0%
#734095000000
1!
1%
#734100000000
0!
0%
#734105000000
1!
1%
#734110000000
0!
0%
#734115000000
1!
1%
#734120000000
0!
0%
#734125000000
1!
1%
#734130000000
0!
0%
#734135000000
1!
1%
#734140000000
0!
0%
#734145000000
1!
1%
#734150000000
0!
0%
#734155000000
1!
1%
#734160000000
0!
0%
#734165000000
1!
1%
#734170000000
0!
0%
#734175000000
1!
1%
#734180000000
0!
0%
#734185000000
1!
1%
#734190000000
0!
0%
#734195000000
1!
1%
#734200000000
0!
0%
#734205000000
1!
1%
#734210000000
0!
0%
#734215000000
1!
1%
#734220000000
0!
0%
#734225000000
1!
1%
#734230000000
0!
0%
#734235000000
1!
1%
#734240000000
0!
0%
#734245000000
1!
1%
#734250000000
0!
0%
#734255000000
1!
1%
#734260000000
0!
0%
#734265000000
1!
1%
#734270000000
0!
0%
#734275000000
1!
1%
#734280000000
0!
0%
#734285000000
1!
1%
#734290000000
0!
0%
#734295000000
1!
1%
#734300000000
0!
0%
#734305000000
1!
1%
#734310000000
0!
0%
#734315000000
1!
1%
#734320000000
0!
0%
#734325000000
1!
1%
#734330000000
0!
0%
#734335000000
1!
1%
#734340000000
0!
0%
#734345000000
1!
1%
#734350000000
0!
0%
#734355000000
1!
1%
#734360000000
0!
0%
#734365000000
1!
1%
#734370000000
0!
0%
#734375000000
1!
1%
#734380000000
0!
0%
#734385000000
1!
1%
#734390000000
0!
0%
#734395000000
1!
1%
#734400000000
0!
0%
#734405000000
1!
1%
#734410000000
0!
0%
#734415000000
1!
1%
#734420000000
0!
0%
#734425000000
1!
1%
#734430000000
0!
0%
#734435000000
1!
1%
#734440000000
0!
0%
#734445000000
1!
1%
#734450000000
0!
0%
#734455000000
1!
1%
#734460000000
0!
0%
#734465000000
1!
1%
#734470000000
0!
0%
#734475000000
1!
1%
#734480000000
0!
0%
#734485000000
1!
1%
#734490000000
0!
0%
#734495000000
1!
1%
#734500000000
0!
0%
#734505000000
1!
1%
#734510000000
0!
0%
#734515000000
1!
1%
#734520000000
0!
0%
#734525000000
1!
1%
#734530000000
0!
0%
#734535000000
1!
1%
#734540000000
0!
0%
#734545000000
1!
1%
#734550000000
0!
0%
#734555000000
1!
1%
#734560000000
0!
0%
#734565000000
1!
1%
#734570000000
0!
0%
#734575000000
1!
1%
#734580000000
0!
0%
#734585000000
1!
1%
#734590000000
0!
0%
#734595000000
1!
1%
#734600000000
0!
0%
#734605000000
1!
1%
#734610000000
0!
0%
#734615000000
1!
1%
#734620000000
0!
0%
#734625000000
1!
1%
#734630000000
0!
0%
#734635000000
1!
1%
#734640000000
0!
0%
#734645000000
1!
1%
#734650000000
0!
0%
#734655000000
1!
1%
#734660000000
0!
0%
#734665000000
1!
1%
#734670000000
0!
0%
#734675000000
1!
1%
#734680000000
0!
0%
#734685000000
1!
1%
#734690000000
0!
0%
#734695000000
1!
1%
#734700000000
0!
0%
#734705000000
1!
1%
#734710000000
0!
0%
#734715000000
1!
1%
#734720000000
0!
0%
#734725000000
1!
1%
#734730000000
0!
0%
#734735000000
1!
1%
#734740000000
0!
0%
#734745000000
1!
1%
#734750000000
0!
0%
#734755000000
1!
1%
#734760000000
0!
0%
#734765000000
1!
1%
#734770000000
0!
0%
#734775000000
1!
1%
#734780000000
0!
0%
#734785000000
1!
1%
#734790000000
0!
0%
#734795000000
1!
1%
#734800000000
0!
0%
#734805000000
1!
1%
#734810000000
0!
0%
#734815000000
1!
1%
#734820000000
0!
0%
#734825000000
1!
1%
#734830000000
0!
0%
#734835000000
1!
1%
#734840000000
0!
0%
#734845000000
1!
1%
#734850000000
0!
0%
#734855000000
1!
1%
#734860000000
0!
0%
#734865000000
1!
1%
#734870000000
0!
0%
#734875000000
1!
1%
#734880000000
0!
0%
#734885000000
1!
1%
#734890000000
0!
0%
#734895000000
1!
1%
#734900000000
0!
0%
#734905000000
1!
1%
#734910000000
0!
0%
#734915000000
1!
1%
#734920000000
0!
0%
#734925000000
1!
1%
#734930000000
0!
0%
#734935000000
1!
1%
#734940000000
0!
0%
#734945000000
1!
1%
#734950000000
0!
0%
#734955000000
1!
1%
#734960000000
0!
0%
#734965000000
1!
1%
#734970000000
0!
0%
#734975000000
1!
1%
#734980000000
0!
0%
#734985000000
1!
1%
#734990000000
0!
0%
#734995000000
1!
1%
#735000000000
0!
0%
#735005000000
1!
1%
#735010000000
0!
0%
#735015000000
1!
1%
#735020000000
0!
0%
#735025000000
1!
1%
#735030000000
0!
0%
#735035000000
1!
1%
#735040000000
0!
0%
#735045000000
1!
1%
#735050000000
0!
0%
#735055000000
1!
1%
#735060000000
0!
0%
#735065000000
1!
1%
#735070000000
0!
0%
#735075000000
1!
1%
#735080000000
0!
0%
#735085000000
1!
1%
#735090000000
0!
0%
#735095000000
1!
1%
#735100000000
0!
0%
#735105000000
1!
1%
#735110000000
0!
0%
#735115000000
1!
1%
#735120000000
0!
0%
#735125000000
1!
1%
#735130000000
0!
0%
#735135000000
1!
1%
#735140000000
0!
0%
#735145000000
1!
1%
#735150000000
0!
0%
#735155000000
1!
1%
#735160000000
0!
0%
#735165000000
1!
1%
#735170000000
0!
0%
#735175000000
1!
1%
#735180000000
0!
0%
#735185000000
1!
1%
#735190000000
0!
0%
#735195000000
1!
1%
#735200000000
0!
0%
#735205000000
1!
1%
#735210000000
0!
0%
#735215000000
1!
1%
#735220000000
0!
0%
#735225000000
1!
1%
#735230000000
0!
0%
#735235000000
1!
1%
#735240000000
0!
0%
#735245000000
1!
1%
#735250000000
0!
0%
#735255000000
1!
1%
#735260000000
0!
0%
#735265000000
1!
1%
#735270000000
0!
0%
#735275000000
1!
1%
#735280000000
0!
0%
#735285000000
1!
1%
#735290000000
0!
0%
#735295000000
1!
1%
#735300000000
0!
0%
#735305000000
1!
1%
#735310000000
0!
0%
#735315000000
1!
1%
#735320000000
0!
0%
#735325000000
1!
1%
#735330000000
0!
0%
#735335000000
1!
1%
#735340000000
0!
0%
#735345000000
1!
1%
#735350000000
0!
0%
#735355000000
1!
1%
#735360000000
0!
0%
#735365000000
1!
1%
#735370000000
0!
0%
#735375000000
1!
1%
#735380000000
0!
0%
#735385000000
1!
1%
#735390000000
0!
0%
#735395000000
1!
1%
#735400000000
0!
0%
#735405000000
1!
1%
#735410000000
0!
0%
#735415000000
1!
1%
#735420000000
0!
0%
#735425000000
1!
1%
#735430000000
0!
0%
#735435000000
1!
1%
#735440000000
0!
0%
#735445000000
1!
1%
#735450000000
0!
0%
#735455000000
1!
1%
#735460000000
0!
0%
#735465000000
1!
1%
#735470000000
0!
0%
#735475000000
1!
1%
#735480000000
0!
0%
#735485000000
1!
1%
#735490000000
0!
0%
#735495000000
1!
1%
#735500000000
0!
0%
#735505000000
1!
1%
#735510000000
0!
0%
#735515000000
1!
1%
#735520000000
0!
0%
#735525000000
1!
1%
#735530000000
0!
0%
#735535000000
1!
1%
#735540000000
0!
0%
#735545000000
1!
1%
#735550000000
0!
0%
#735555000000
1!
1%
#735560000000
0!
0%
#735565000000
1!
1%
#735570000000
0!
0%
#735575000000
1!
1%
#735580000000
0!
0%
#735585000000
1!
1%
#735590000000
0!
0%
#735595000000
1!
1%
#735600000000
0!
0%
#735605000000
1!
1%
#735610000000
0!
0%
#735615000000
1!
1%
#735620000000
0!
0%
#735625000000
1!
1%
#735630000000
0!
0%
#735635000000
1!
1%
#735640000000
0!
0%
#735645000000
1!
1%
#735650000000
0!
0%
#735655000000
1!
1%
#735660000000
0!
0%
#735665000000
1!
1%
#735670000000
0!
0%
#735675000000
1!
1%
#735680000000
0!
0%
#735685000000
1!
1%
#735690000000
0!
0%
#735695000000
1!
1%
#735700000000
0!
0%
#735705000000
1!
1%
#735710000000
0!
0%
#735715000000
1!
1%
#735720000000
0!
0%
#735725000000
1!
1%
#735730000000
0!
0%
#735735000000
1!
1%
#735740000000
0!
0%
#735745000000
1!
1%
#735750000000
0!
0%
#735755000000
1!
1%
#735760000000
0!
0%
#735765000000
1!
1%
#735770000000
0!
0%
#735775000000
1!
1%
#735780000000
0!
0%
#735785000000
1!
1%
#735790000000
0!
0%
#735795000000
1!
1%
#735800000000
0!
0%
#735805000000
1!
1%
#735810000000
0!
0%
#735815000000
1!
1%
#735820000000
0!
0%
#735825000000
1!
1%
#735830000000
0!
0%
#735835000000
1!
1%
#735840000000
0!
0%
#735845000000
1!
1%
#735850000000
0!
0%
#735855000000
1!
1%
#735860000000
0!
0%
#735865000000
1!
1%
#735870000000
0!
0%
#735875000000
1!
1%
#735880000000
0!
0%
#735885000000
1!
1%
#735890000000
0!
0%
#735895000000
1!
1%
#735900000000
0!
0%
#735905000000
1!
1%
#735910000000
0!
0%
#735915000000
1!
1%
#735920000000
0!
0%
#735925000000
1!
1%
#735930000000
0!
0%
#735935000000
1!
1%
#735940000000
0!
0%
#735945000000
1!
1%
#735950000000
0!
0%
#735955000000
1!
1%
#735960000000
0!
0%
#735965000000
1!
1%
#735970000000
0!
0%
#735975000000
1!
1%
#735980000000
0!
0%
#735985000000
1!
1%
#735990000000
0!
0%
#735995000000
1!
1%
#736000000000
0!
0%
#736005000000
1!
1%
#736010000000
0!
0%
#736015000000
1!
1%
#736020000000
0!
0%
#736025000000
1!
1%
#736030000000
0!
0%
#736035000000
1!
1%
#736040000000
0!
0%
#736045000000
1!
1%
#736050000000
0!
0%
#736055000000
1!
1%
#736060000000
0!
0%
#736065000000
1!
1%
#736070000000
0!
0%
#736075000000
1!
1%
#736080000000
0!
0%
#736085000000
1!
1%
#736090000000
0!
0%
#736095000000
1!
1%
#736100000000
0!
0%
#736105000000
1!
1%
#736110000000
0!
0%
#736115000000
1!
1%
#736120000000
0!
0%
#736125000000
1!
1%
#736130000000
0!
0%
#736135000000
1!
1%
#736140000000
0!
0%
#736145000000
1!
1%
#736150000000
0!
0%
#736155000000
1!
1%
#736160000000
0!
0%
#736165000000
1!
1%
#736170000000
0!
0%
#736175000000
1!
1%
#736180000000
0!
0%
#736185000000
1!
1%
#736190000000
0!
0%
#736195000000
1!
1%
#736200000000
0!
0%
#736205000000
1!
1%
#736210000000
0!
0%
#736215000000
1!
1%
#736220000000
0!
0%
#736225000000
1!
1%
#736230000000
0!
0%
#736235000000
1!
1%
#736240000000
0!
0%
#736245000000
1!
1%
#736250000000
0!
0%
#736255000000
1!
1%
#736260000000
0!
0%
#736265000000
1!
1%
#736270000000
0!
0%
#736275000000
1!
1%
#736280000000
0!
0%
#736285000000
1!
1%
#736290000000
0!
0%
#736295000000
1!
1%
#736300000000
0!
0%
#736305000000
1!
1%
#736310000000
0!
0%
#736315000000
1!
1%
#736320000000
0!
0%
#736325000000
1!
1%
#736330000000
0!
0%
#736335000000
1!
1%
#736340000000
0!
0%
#736345000000
1!
1%
#736350000000
0!
0%
#736355000000
1!
1%
#736360000000
0!
0%
#736365000000
1!
1%
#736370000000
0!
0%
#736375000000
1!
1%
#736380000000
0!
0%
#736385000000
1!
1%
#736390000000
0!
0%
#736395000000
1!
1%
#736400000000
0!
0%
#736405000000
1!
1%
#736410000000
0!
0%
#736415000000
1!
1%
#736420000000
0!
0%
#736425000000
1!
1%
#736430000000
0!
0%
#736435000000
1!
1%
#736440000000
0!
0%
#736445000000
1!
1%
#736450000000
0!
0%
#736455000000
1!
1%
#736460000000
0!
0%
#736465000000
1!
1%
#736470000000
0!
0%
#736475000000
1!
1%
#736480000000
0!
0%
#736485000000
1!
1%
#736490000000
0!
0%
#736495000000
1!
1%
#736500000000
0!
0%
#736505000000
1!
1%
#736510000000
0!
0%
#736515000000
1!
1%
#736520000000
0!
0%
#736525000000
1!
1%
#736530000000
0!
0%
#736535000000
1!
1%
#736540000000
0!
0%
#736545000000
1!
1%
#736550000000
0!
0%
#736555000000
1!
1%
#736560000000
0!
0%
#736565000000
1!
1%
#736570000000
0!
0%
#736575000000
1!
1%
#736580000000
0!
0%
#736585000000
1!
1%
#736590000000
0!
0%
#736595000000
1!
1%
#736600000000
0!
0%
#736605000000
1!
1%
#736610000000
0!
0%
#736615000000
1!
1%
#736620000000
0!
0%
#736625000000
1!
1%
#736630000000
0!
0%
#736635000000
1!
1%
#736640000000
0!
0%
#736645000000
1!
1%
#736650000000
0!
0%
#736655000000
1!
1%
#736660000000
0!
0%
#736665000000
1!
1%
#736670000000
0!
0%
#736675000000
1!
1%
#736680000000
0!
0%
#736685000000
1!
1%
#736690000000
0!
0%
#736695000000
1!
1%
#736700000000
0!
0%
#736705000000
1!
1%
#736710000000
0!
0%
#736715000000
1!
1%
#736720000000
0!
0%
#736725000000
1!
1%
#736730000000
0!
0%
#736735000000
1!
1%
#736740000000
0!
0%
#736745000000
1!
1%
#736750000000
0!
0%
#736755000000
1!
1%
#736760000000
0!
0%
#736765000000
1!
1%
#736770000000
0!
0%
#736775000000
1!
1%
#736780000000
0!
0%
#736785000000
1!
1%
#736790000000
0!
0%
#736795000000
1!
1%
#736800000000
0!
0%
#736805000000
1!
1%
#736810000000
0!
0%
#736815000000
1!
1%
#736820000000
0!
0%
#736825000000
1!
1%
#736830000000
0!
0%
#736835000000
1!
1%
#736840000000
0!
0%
#736845000000
1!
1%
#736850000000
0!
0%
#736855000000
1!
1%
#736860000000
0!
0%
#736865000000
1!
1%
#736870000000
0!
0%
#736875000000
1!
1%
#736880000000
0!
0%
#736885000000
1!
1%
#736890000000
0!
0%
#736895000000
1!
1%
#736900000000
0!
0%
#736905000000
1!
1%
#736910000000
0!
0%
#736915000000
1!
1%
#736920000000
0!
0%
#736925000000
1!
1%
#736930000000
0!
0%
#736935000000
1!
1%
#736940000000
0!
0%
#736945000000
1!
1%
#736950000000
0!
0%
#736955000000
1!
1%
#736960000000
0!
0%
#736965000000
1!
1%
#736970000000
0!
0%
#736975000000
1!
1%
#736980000000
0!
0%
#736985000000
1!
1%
#736990000000
0!
0%
#736995000000
1!
1%
#737000000000
0!
0%
#737005000000
1!
1%
#737010000000
0!
0%
#737015000000
1!
1%
#737020000000
0!
0%
#737025000000
1!
1%
#737030000000
0!
0%
#737035000000
1!
1%
#737040000000
0!
0%
#737045000000
1!
1%
#737050000000
0!
0%
#737055000000
1!
1%
#737060000000
0!
0%
#737065000000
1!
1%
#737070000000
0!
0%
#737075000000
1!
1%
#737080000000
0!
0%
#737085000000
1!
1%
#737090000000
0!
0%
#737095000000
1!
1%
#737100000000
0!
0%
#737105000000
1!
1%
#737110000000
0!
0%
#737115000000
1!
1%
#737120000000
0!
0%
#737125000000
1!
1%
#737130000000
0!
0%
#737135000000
1!
1%
#737140000000
0!
0%
#737145000000
1!
1%
#737150000000
0!
0%
#737155000000
1!
1%
#737160000000
0!
0%
#737165000000
1!
1%
#737170000000
0!
0%
#737175000000
1!
1%
#737180000000
0!
0%
#737185000000
1!
1%
#737190000000
0!
0%
#737195000000
1!
1%
#737200000000
0!
0%
#737205000000
1!
1%
#737210000000
0!
0%
#737215000000
1!
1%
#737220000000
0!
0%
#737225000000
1!
1%
#737230000000
0!
0%
#737235000000
1!
1%
#737240000000
0!
0%
#737245000000
1!
1%
#737250000000
0!
0%
#737255000000
1!
1%
#737260000000
0!
0%
#737265000000
1!
1%
#737270000000
0!
0%
#737275000000
1!
1%
#737280000000
0!
0%
#737285000000
1!
1%
#737290000000
0!
0%
#737295000000
1!
1%
#737300000000
0!
0%
#737305000000
1!
1%
#737310000000
0!
0%
#737315000000
1!
1%
#737320000000
0!
0%
#737325000000
1!
1%
#737330000000
0!
0%
#737335000000
1!
1%
#737340000000
0!
0%
#737345000000
1!
1%
#737350000000
0!
0%
#737355000000
1!
1%
#737360000000
0!
0%
#737365000000
1!
1%
#737370000000
0!
0%
#737375000000
1!
1%
#737380000000
0!
0%
#737385000000
1!
1%
#737390000000
0!
0%
#737395000000
1!
1%
#737400000000
0!
0%
#737405000000
1!
1%
#737410000000
0!
0%
#737415000000
1!
1%
#737420000000
0!
0%
#737425000000
1!
1%
#737430000000
0!
0%
#737435000000
1!
1%
#737440000000
0!
0%
#737445000000
1!
1%
#737450000000
0!
0%
#737455000000
1!
1%
#737460000000
0!
0%
#737465000000
1!
1%
#737470000000
0!
0%
#737475000000
1!
1%
#737480000000
0!
0%
#737485000000
1!
1%
#737490000000
0!
0%
#737495000000
1!
1%
#737500000000
0!
0%
#737505000000
1!
1%
#737510000000
0!
0%
#737515000000
1!
1%
#737520000000
0!
0%
#737525000000
1!
1%
#737530000000
0!
0%
#737535000000
1!
1%
#737540000000
0!
0%
#737545000000
1!
1%
#737550000000
0!
0%
#737555000000
1!
1%
#737560000000
0!
0%
#737565000000
1!
1%
#737570000000
0!
0%
#737575000000
1!
1%
#737580000000
0!
0%
#737585000000
1!
1%
#737590000000
0!
0%
#737595000000
1!
1%
#737600000000
0!
0%
#737605000000
1!
1%
#737610000000
0!
0%
#737615000000
1!
1%
#737620000000
0!
0%
#737625000000
1!
1%
#737630000000
0!
0%
#737635000000
1!
1%
#737640000000
0!
0%
#737645000000
1!
1%
#737650000000
0!
0%
#737655000000
1!
1%
#737660000000
0!
0%
#737665000000
1!
1%
#737670000000
0!
0%
#737675000000
1!
1%
#737680000000
0!
0%
#737685000000
1!
1%
#737690000000
0!
0%
#737695000000
1!
1%
#737700000000
0!
0%
#737705000000
1!
1%
#737710000000
0!
0%
#737715000000
1!
1%
#737720000000
0!
0%
#737725000000
1!
1%
#737730000000
0!
0%
#737735000000
1!
1%
#737740000000
0!
0%
#737745000000
1!
1%
#737750000000
0!
0%
#737755000000
1!
1%
#737760000000
0!
0%
#737765000000
1!
1%
#737770000000
0!
0%
#737775000000
1!
1%
#737780000000
0!
0%
#737785000000
1!
1%
#737790000000
0!
0%
#737795000000
1!
1%
#737800000000
0!
0%
#737805000000
1!
1%
#737810000000
0!
0%
#737815000000
1!
1%
#737820000000
0!
0%
#737825000000
1!
1%
#737830000000
0!
0%
#737835000000
1!
1%
#737840000000
0!
0%
#737845000000
1!
1%
#737850000000
0!
0%
#737855000000
1!
1%
#737860000000
0!
0%
#737865000000
1!
1%
#737870000000
0!
0%
#737875000000
1!
1%
#737880000000
0!
0%
#737885000000
1!
1%
#737890000000
0!
0%
#737895000000
1!
1%
#737900000000
0!
0%
#737905000000
1!
1%
#737910000000
0!
0%
#737915000000
1!
1%
#737920000000
0!
0%
#737925000000
1!
1%
#737930000000
0!
0%
#737935000000
1!
1%
#737940000000
0!
0%
#737945000000
1!
1%
#737950000000
0!
0%
#737955000000
1!
1%
#737960000000
0!
0%
#737965000000
1!
1%
#737970000000
0!
0%
#737975000000
1!
1%
#737980000000
0!
0%
#737985000000
1!
1%
#737990000000
0!
0%
#737995000000
1!
1%
#738000000000
0!
0%
#738005000000
1!
1%
#738010000000
0!
0%
#738015000000
1!
1%
#738020000000
0!
0%
#738025000000
1!
1%
#738030000000
0!
0%
#738035000000
1!
1%
#738040000000
0!
0%
#738045000000
1!
1%
#738050000000
0!
0%
#738055000000
1!
1%
#738060000000
0!
0%
#738065000000
1!
1%
#738070000000
0!
0%
#738075000000
1!
1%
#738080000000
0!
0%
#738085000000
1!
1%
#738090000000
0!
0%
#738095000000
1!
1%
#738100000000
0!
0%
#738105000000
1!
1%
#738110000000
0!
0%
#738115000000
1!
1%
#738120000000
0!
0%
#738125000000
1!
1%
#738130000000
0!
0%
#738135000000
1!
1%
#738140000000
0!
0%
#738145000000
1!
1%
#738150000000
0!
0%
#738155000000
1!
1%
#738160000000
0!
0%
#738165000000
1!
1%
#738170000000
0!
0%
#738175000000
1!
1%
#738180000000
0!
0%
#738185000000
1!
1%
#738190000000
0!
0%
#738195000000
1!
1%
#738200000000
0!
0%
#738205000000
1!
1%
#738210000000
0!
0%
#738215000000
1!
1%
#738220000000
0!
0%
#738225000000
1!
1%
#738230000000
0!
0%
#738235000000
1!
1%
#738240000000
0!
0%
#738245000000
1!
1%
#738250000000
0!
0%
#738255000000
1!
1%
#738260000000
0!
0%
#738265000000
1!
1%
#738270000000
0!
0%
#738275000000
1!
1%
#738280000000
0!
0%
#738285000000
1!
1%
#738290000000
0!
0%
#738295000000
1!
1%
#738300000000
0!
0%
#738305000000
1!
1%
#738310000000
0!
0%
#738315000000
1!
1%
#738320000000
0!
0%
#738325000000
1!
1%
#738330000000
0!
0%
#738335000000
1!
1%
#738340000000
0!
0%
#738345000000
1!
1%
#738350000000
0!
0%
#738355000000
1!
1%
#738360000000
0!
0%
#738365000000
1!
1%
#738370000000
0!
0%
#738375000000
1!
1%
#738380000000
0!
0%
#738385000000
1!
1%
#738390000000
0!
0%
#738395000000
1!
1%
#738400000000
0!
0%
#738405000000
1!
1%
#738410000000
0!
0%
#738415000000
1!
1%
#738420000000
0!
0%
#738425000000
1!
1%
#738430000000
0!
0%
#738435000000
1!
1%
#738440000000
0!
0%
#738445000000
1!
1%
#738450000000
0!
0%
#738455000000
1!
1%
#738460000000
0!
0%
#738465000000
1!
1%
#738470000000
0!
0%
#738475000000
1!
1%
#738480000000
0!
0%
#738485000000
1!
1%
#738490000000
0!
0%
#738495000000
1!
1%
#738500000000
0!
0%
#738505000000
1!
1%
#738510000000
0!
0%
#738515000000
1!
1%
#738520000000
0!
0%
#738525000000
1!
1%
#738530000000
0!
0%
#738535000000
1!
1%
#738540000000
0!
0%
#738545000000
1!
1%
#738550000000
0!
0%
#738555000000
1!
1%
#738560000000
0!
0%
#738565000000
1!
1%
#738570000000
0!
0%
#738575000000
1!
1%
#738580000000
0!
0%
#738585000000
1!
1%
#738590000000
0!
0%
#738595000000
1!
1%
#738600000000
0!
0%
#738605000000
1!
1%
#738610000000
0!
0%
#738615000000
1!
1%
#738620000000
0!
0%
#738625000000
1!
1%
#738630000000
0!
0%
#738635000000
1!
1%
#738640000000
0!
0%
#738645000000
1!
1%
#738650000000
0!
0%
#738655000000
1!
1%
#738660000000
0!
0%
#738665000000
1!
1%
#738670000000
0!
0%
#738675000000
1!
1%
#738680000000
0!
0%
#738685000000
1!
1%
#738690000000
0!
0%
#738695000000
1!
1%
#738700000000
0!
0%
#738705000000
1!
1%
#738710000000
0!
0%
#738715000000
1!
1%
#738720000000
0!
0%
#738725000000
1!
1%
#738730000000
0!
0%
#738735000000
1!
1%
#738740000000
0!
0%
#738745000000
1!
1%
#738750000000
0!
0%
#738755000000
1!
1%
#738760000000
0!
0%
#738765000000
1!
1%
#738770000000
0!
0%
#738775000000
1!
1%
#738780000000
0!
0%
#738785000000
1!
1%
#738790000000
0!
0%
#738795000000
1!
1%
#738800000000
0!
0%
#738805000000
1!
1%
#738810000000
0!
0%
#738815000000
1!
1%
#738820000000
0!
0%
#738825000000
1!
1%
#738830000000
0!
0%
#738835000000
1!
1%
#738840000000
0!
0%
#738845000000
1!
1%
#738850000000
0!
0%
#738855000000
1!
1%
#738860000000
0!
0%
#738865000000
1!
1%
#738870000000
0!
0%
#738875000000
1!
1%
#738880000000
0!
0%
#738885000000
1!
1%
#738890000000
0!
0%
#738895000000
1!
1%
#738900000000
0!
0%
#738905000000
1!
1%
#738910000000
0!
0%
#738915000000
1!
1%
#738920000000
0!
0%
#738925000000
1!
1%
#738930000000
0!
0%
#738935000000
1!
1%
#738940000000
0!
0%
#738945000000
1!
1%
#738950000000
0!
0%
#738955000000
1!
1%
#738960000000
0!
0%
#738965000000
1!
1%
#738970000000
0!
0%
#738975000000
1!
1%
#738980000000
0!
0%
#738985000000
1!
1%
#738990000000
0!
0%
#738995000000
1!
1%
#739000000000
0!
0%
#739005000000
1!
1%
#739010000000
0!
0%
#739015000000
1!
1%
#739020000000
0!
0%
#739025000000
1!
1%
#739030000000
0!
0%
#739035000000
1!
1%
#739040000000
0!
0%
#739045000000
1!
1%
#739050000000
0!
0%
#739055000000
1!
1%
#739060000000
0!
0%
#739065000000
1!
1%
#739070000000
0!
0%
#739075000000
1!
1%
#739080000000
0!
0%
#739085000000
1!
1%
#739090000000
0!
0%
#739095000000
1!
1%
#739100000000
0!
0%
#739105000000
1!
1%
#739110000000
0!
0%
#739115000000
1!
1%
#739120000000
0!
0%
#739125000000
1!
1%
#739130000000
0!
0%
#739135000000
1!
1%
#739140000000
0!
0%
#739145000000
1!
1%
#739150000000
0!
0%
#739155000000
1!
1%
#739160000000
0!
0%
#739165000000
1!
1%
#739170000000
0!
0%
#739175000000
1!
1%
#739180000000
0!
0%
#739185000000
1!
1%
#739190000000
0!
0%
#739195000000
1!
1%
#739200000000
0!
0%
#739205000000
1!
1%
#739210000000
0!
0%
#739215000000
1!
1%
#739220000000
0!
0%
#739225000000
1!
1%
#739230000000
0!
0%
#739235000000
1!
1%
#739240000000
0!
0%
#739245000000
1!
1%
#739250000000
0!
0%
#739255000000
1!
1%
#739260000000
0!
0%
#739265000000
1!
1%
#739270000000
0!
0%
#739275000000
1!
1%
#739280000000
0!
0%
#739285000000
1!
1%
#739290000000
0!
0%
#739295000000
1!
1%
#739300000000
0!
0%
#739305000000
1!
1%
#739310000000
0!
0%
#739315000000
1!
1%
#739320000000
0!
0%
#739325000000
1!
1%
#739330000000
0!
0%
#739335000000
1!
1%
#739340000000
0!
0%
#739345000000
1!
1%
#739350000000
0!
0%
#739355000000
1!
1%
#739360000000
0!
0%
#739365000000
1!
1%
#739370000000
0!
0%
#739375000000
1!
1%
#739380000000
0!
0%
#739385000000
1!
1%
#739390000000
0!
0%
#739395000000
1!
1%
#739400000000
0!
0%
#739405000000
1!
1%
#739410000000
0!
0%
#739415000000
1!
1%
#739420000000
0!
0%
#739425000000
1!
1%
#739430000000
0!
0%
#739435000000
1!
1%
#739440000000
0!
0%
#739445000000
1!
1%
#739450000000
0!
0%
#739455000000
1!
1%
#739460000000
0!
0%
#739465000000
1!
1%
#739470000000
0!
0%
#739475000000
1!
1%
#739480000000
0!
0%
#739485000000
1!
1%
#739490000000
0!
0%
#739495000000
1!
1%
#739500000000
0!
0%
#739505000000
1!
1%
#739510000000
0!
0%
#739515000000
1!
1%
#739520000000
0!
0%
#739525000000
1!
1%
#739530000000
0!
0%
#739535000000
1!
1%
#739540000000
0!
0%
#739545000000
1!
1%
#739550000000
0!
0%
#739555000000
1!
1%
#739560000000
0!
0%
#739565000000
1!
1%
#739570000000
0!
0%
#739575000000
1!
1%
#739580000000
0!
0%
#739585000000
1!
1%
#739590000000
0!
0%
#739595000000
1!
1%
#739600000000
0!
0%
#739605000000
1!
1%
#739610000000
0!
0%
#739615000000
1!
1%
#739620000000
0!
0%
#739625000000
1!
1%
#739630000000
0!
0%
#739635000000
1!
1%
#739640000000
0!
0%
#739645000000
1!
1%
#739650000000
0!
0%
#739655000000
1!
1%
#739660000000
0!
0%
#739665000000
1!
1%
#739670000000
0!
0%
#739675000000
1!
1%
#739680000000
0!
0%
#739685000000
1!
1%
#739690000000
0!
0%
#739695000000
1!
1%
#739700000000
0!
0%
#739705000000
1!
1%
#739710000000
0!
0%
#739715000000
1!
1%
#739720000000
0!
0%
#739725000000
1!
1%
#739730000000
0!
0%
#739735000000
1!
1%
#739740000000
0!
0%
#739745000000
1!
1%
#739750000000
0!
0%
#739755000000
1!
1%
#739760000000
0!
0%
#739765000000
1!
1%
#739770000000
0!
0%
#739775000000
1!
1%
#739780000000
0!
0%
#739785000000
1!
1%
#739790000000
0!
0%
#739795000000
1!
1%
#739800000000
0!
0%
#739805000000
1!
1%
#739810000000
0!
0%
#739815000000
1!
1%
#739820000000
0!
0%
#739825000000
1!
1%
#739830000000
0!
0%
#739835000000
1!
1%
#739840000000
0!
0%
#739845000000
1!
1%
#739850000000
0!
0%
#739855000000
1!
1%
#739860000000
0!
0%
#739865000000
1!
1%
#739870000000
0!
0%
#739875000000
1!
1%
#739880000000
0!
0%
#739885000000
1!
1%
#739890000000
0!
0%
#739895000000
1!
1%
#739900000000
0!
0%
#739905000000
1!
1%
#739910000000
0!
0%
#739915000000
1!
1%
#739920000000
0!
0%
#739925000000
1!
1%
#739930000000
0!
0%
#739935000000
1!
1%
#739940000000
0!
0%
#739945000000
1!
1%
#739950000000
0!
0%
#739955000000
1!
1%
#739960000000
0!
0%
#739965000000
1!
1%
#739970000000
0!
0%
#739975000000
1!
1%
#739980000000
0!
0%
#739985000000
1!
1%
#739990000000
0!
0%
#739995000000
1!
1%
#740000000000
0!
0%
#740005000000
1!
1%
#740010000000
0!
0%
#740015000000
1!
1%
#740020000000
0!
0%
#740025000000
1!
1%
#740030000000
0!
0%
#740035000000
1!
1%
#740040000000
0!
0%
#740045000000
1!
1%
#740050000000
0!
0%
#740055000000
1!
1%
#740060000000
0!
0%
#740065000000
1!
1%
#740070000000
0!
0%
#740075000000
1!
1%
#740080000000
0!
0%
#740085000000
1!
1%
#740090000000
0!
0%
#740095000000
1!
1%
#740100000000
0!
0%
#740105000000
1!
1%
#740110000000
0!
0%
#740115000000
1!
1%
#740120000000
0!
0%
#740125000000
1!
1%
#740130000000
0!
0%
#740135000000
1!
1%
#740140000000
0!
0%
#740145000000
1!
1%
#740150000000
0!
0%
#740155000000
1!
1%
#740160000000
0!
0%
#740165000000
1!
1%
#740170000000
0!
0%
#740175000000
1!
1%
#740180000000
0!
0%
#740185000000
1!
1%
#740190000000
0!
0%
#740195000000
1!
1%
#740200000000
0!
0%
#740205000000
1!
1%
#740210000000
0!
0%
#740215000000
1!
1%
#740220000000
0!
0%
#740225000000
1!
1%
#740230000000
0!
0%
#740235000000
1!
1%
#740240000000
0!
0%
#740245000000
1!
1%
#740250000000
0!
0%
#740255000000
1!
1%
#740260000000
0!
0%
#740265000000
1!
1%
#740270000000
0!
0%
#740275000000
1!
1%
#740280000000
0!
0%
#740285000000
1!
1%
#740290000000
0!
0%
#740295000000
1!
1%
#740300000000
0!
0%
#740305000000
1!
1%
#740310000000
0!
0%
#740315000000
1!
1%
#740320000000
0!
0%
#740325000000
1!
1%
#740330000000
0!
0%
#740335000000
1!
1%
#740340000000
0!
0%
#740345000000
1!
1%
#740350000000
0!
0%
#740355000000
1!
1%
#740360000000
0!
0%
#740365000000
1!
1%
#740370000000
0!
0%
#740375000000
1!
1%
#740380000000
0!
0%
#740385000000
1!
1%
#740390000000
0!
0%
#740395000000
1!
1%
#740400000000
0!
0%
#740405000000
1!
1%
#740410000000
0!
0%
#740415000000
1!
1%
#740420000000
0!
0%
#740425000000
1!
1%
#740430000000
0!
0%
#740435000000
1!
1%
#740440000000
0!
0%
#740445000000
1!
1%
#740450000000
0!
0%
#740455000000
1!
1%
#740460000000
0!
0%
#740465000000
1!
1%
#740470000000
0!
0%
#740475000000
1!
1%
#740480000000
0!
0%
#740485000000
1!
1%
#740490000000
0!
0%
#740495000000
1!
1%
#740500000000
0!
0%
#740505000000
1!
1%
#740510000000
0!
0%
#740515000000
1!
1%
#740520000000
0!
0%
#740525000000
1!
1%
#740530000000
0!
0%
#740535000000
1!
1%
#740540000000
0!
0%
#740545000000
1!
1%
#740550000000
0!
0%
#740555000000
1!
1%
#740560000000
0!
0%
#740565000000
1!
1%
#740570000000
0!
0%
#740575000000
1!
1%
#740580000000
0!
0%
#740585000000
1!
1%
#740590000000
0!
0%
#740595000000
1!
1%
#740600000000
0!
0%
#740605000000
1!
1%
#740610000000
0!
0%
#740615000000
1!
1%
#740620000000
0!
0%
#740625000000
1!
1%
#740630000000
0!
0%
#740635000000
1!
1%
#740640000000
0!
0%
#740645000000
1!
1%
#740650000000
0!
0%
#740655000000
1!
1%
#740660000000
0!
0%
#740665000000
1!
1%
#740670000000
0!
0%
#740675000000
1!
1%
#740680000000
0!
0%
#740685000000
1!
1%
#740690000000
0!
0%
#740695000000
1!
1%
#740700000000
0!
0%
#740705000000
1!
1%
#740710000000
0!
0%
#740715000000
1!
1%
#740720000000
0!
0%
#740725000000
1!
1%
#740730000000
0!
0%
#740735000000
1!
1%
#740740000000
0!
0%
#740745000000
1!
1%
#740750000000
0!
0%
#740755000000
1!
1%
#740760000000
0!
0%
#740765000000
1!
1%
#740770000000
0!
0%
#740775000000
1!
1%
#740780000000
0!
0%
#740785000000
1!
1%
#740790000000
0!
0%
#740795000000
1!
1%
#740800000000
0!
0%
#740805000000
1!
1%
#740810000000
0!
0%
#740815000000
1!
1%
#740820000000
0!
0%
#740825000000
1!
1%
#740830000000
0!
0%
#740835000000
1!
1%
#740840000000
0!
0%
#740845000000
1!
1%
#740850000000
0!
0%
#740855000000
1!
1%
#740860000000
0!
0%
#740865000000
1!
1%
#740870000000
0!
0%
#740875000000
1!
1%
#740880000000
0!
0%
#740885000000
1!
1%
#740890000000
0!
0%
#740895000000
1!
1%
#740900000000
0!
0%
#740905000000
1!
1%
#740910000000
0!
0%
#740915000000
1!
1%
#740920000000
0!
0%
#740925000000
1!
1%
#740930000000
0!
0%
#740935000000
1!
1%
#740940000000
0!
0%
#740945000000
1!
1%
#740950000000
0!
0%
#740955000000
1!
1%
#740960000000
0!
0%
#740965000000
1!
1%
#740970000000
0!
0%
#740975000000
1!
1%
#740980000000
0!
0%
#740985000000
1!
1%
#740990000000
0!
0%
#740995000000
1!
1%
#741000000000
0!
0%
#741005000000
1!
1%
#741010000000
0!
0%
#741015000000
1!
1%
#741020000000
0!
0%
#741025000000
1!
1%
#741030000000
0!
0%
#741035000000
1!
1%
#741040000000
0!
0%
#741045000000
1!
1%
#741050000000
0!
0%
#741055000000
1!
1%
#741060000000
0!
0%
#741065000000
1!
1%
#741070000000
0!
0%
#741075000000
1!
1%
#741080000000
0!
0%
#741085000000
1!
1%
#741090000000
0!
0%
#741095000000
1!
1%
#741100000000
0!
0%
#741105000000
1!
1%
#741110000000
0!
0%
#741115000000
1!
1%
#741120000000
0!
0%
#741125000000
1!
1%
#741130000000
0!
0%
#741135000000
1!
1%
#741140000000
0!
0%
#741145000000
1!
1%
#741150000000
0!
0%
#741155000000
1!
1%
#741160000000
0!
0%
#741165000000
1!
1%
#741170000000
0!
0%
#741175000000
1!
1%
#741180000000
0!
0%
#741185000000
1!
1%
#741190000000
0!
0%
#741195000000
1!
1%
#741200000000
0!
0%
#741205000000
1!
1%
#741210000000
0!
0%
#741215000000
1!
1%
#741220000000
0!
0%
#741225000000
1!
1%
#741230000000
0!
0%
#741235000000
1!
1%
#741240000000
0!
0%
#741245000000
1!
1%
#741250000000
0!
0%
#741255000000
1!
1%
#741260000000
0!
0%
#741265000000
1!
1%
#741270000000
0!
0%
#741275000000
1!
1%
#741280000000
0!
0%
#741285000000
1!
1%
#741290000000
0!
0%
#741295000000
1!
1%
#741300000000
0!
0%
#741305000000
1!
1%
#741310000000
0!
0%
#741315000000
1!
1%
#741320000000
0!
0%
#741325000000
1!
1%
#741330000000
0!
0%
#741335000000
1!
1%
#741340000000
0!
0%
#741345000000
1!
1%
#741350000000
0!
0%
#741355000000
1!
1%
#741360000000
0!
0%
#741365000000
1!
1%
#741370000000
0!
0%
#741375000000
1!
1%
#741380000000
0!
0%
#741385000000
1!
1%
#741390000000
0!
0%
#741395000000
1!
1%
#741400000000
0!
0%
#741405000000
1!
1%
#741410000000
0!
0%
#741415000000
1!
1%
#741420000000
0!
0%
#741425000000
1!
1%
#741430000000
0!
0%
#741435000000
1!
1%
#741440000000
0!
0%
#741445000000
1!
1%
#741450000000
0!
0%
#741455000000
1!
1%
#741460000000
0!
0%
#741465000000
1!
1%
#741470000000
0!
0%
#741475000000
1!
1%
#741480000000
0!
0%
#741485000000
1!
1%
#741490000000
0!
0%
#741495000000
1!
1%
#741500000000
0!
0%
#741505000000
1!
1%
#741510000000
0!
0%
#741515000000
1!
1%
#741520000000
0!
0%
#741525000000
1!
1%
#741530000000
0!
0%
#741535000000
1!
1%
#741540000000
0!
0%
#741545000000
1!
1%
#741550000000
0!
0%
#741555000000
1!
1%
#741560000000
0!
0%
#741565000000
1!
1%
#741570000000
0!
0%
#741575000000
1!
1%
#741580000000
0!
0%
#741585000000
1!
1%
#741590000000
0!
0%
#741595000000
1!
1%
#741600000000
0!
0%
#741605000000
1!
1%
#741610000000
0!
0%
#741615000000
1!
1%
#741620000000
0!
0%
#741625000000
1!
1%
#741630000000
0!
0%
#741635000000
1!
1%
#741640000000
0!
0%
#741645000000
1!
1%
#741650000000
0!
0%
#741655000000
1!
1%
#741660000000
0!
0%
#741665000000
1!
1%
#741670000000
0!
0%
#741675000000
1!
1%
#741680000000
0!
0%
#741685000000
1!
1%
#741690000000
0!
0%
#741695000000
1!
1%
#741700000000
0!
0%
#741705000000
1!
1%
#741710000000
0!
0%
#741715000000
1!
1%
#741720000000
0!
0%
#741725000000
1!
1%
#741730000000
0!
0%
#741735000000
1!
1%
#741740000000
0!
0%
#741745000000
1!
1%
#741750000000
0!
0%
#741755000000
1!
1%
#741760000000
0!
0%
#741765000000
1!
1%
#741770000000
0!
0%
#741775000000
1!
1%
#741780000000
0!
0%
#741785000000
1!
1%
#741790000000
0!
0%
#741795000000
1!
1%
#741800000000
0!
0%
#741805000000
1!
1%
#741810000000
0!
0%
#741815000000
1!
1%
#741820000000
0!
0%
#741825000000
1!
1%
#741830000000
0!
0%
#741835000000
1!
1%
#741840000000
0!
0%
#741845000000
1!
1%
#741850000000
0!
0%
#741855000000
1!
1%
#741860000000
0!
0%
#741865000000
1!
1%
#741870000000
0!
0%
#741875000000
1!
1%
#741880000000
0!
0%
#741885000000
1!
1%
#741890000000
0!
0%
#741895000000
1!
1%
#741900000000
0!
0%
#741905000000
1!
1%
#741910000000
0!
0%
#741915000000
1!
1%
#741920000000
0!
0%
#741925000000
1!
1%
#741930000000
0!
0%
#741935000000
1!
1%
#741940000000
0!
0%
#741945000000
1!
1%
#741950000000
0!
0%
#741955000000
1!
1%
#741960000000
0!
0%
#741965000000
1!
1%
#741970000000
0!
0%
#741975000000
1!
1%
#741980000000
0!
0%
#741985000000
1!
1%
#741990000000
0!
0%
#741995000000
1!
1%
#742000000000
0!
0%
#742005000000
1!
1%
#742010000000
0!
0%
#742015000000
1!
1%
#742020000000
0!
0%
#742025000000
1!
1%
#742030000000
0!
0%
#742035000000
1!
1%
#742040000000
0!
0%
#742045000000
1!
1%
#742050000000
0!
0%
#742055000000
1!
1%
#742060000000
0!
0%
#742065000000
1!
1%
#742070000000
0!
0%
#742075000000
1!
1%
#742080000000
0!
0%
#742085000000
1!
1%
#742090000000
0!
0%
#742095000000
1!
1%
#742100000000
0!
0%
#742105000000
1!
1%
#742110000000
0!
0%
#742115000000
1!
1%
#742120000000
0!
0%
#742125000000
1!
1%
#742130000000
0!
0%
#742135000000
1!
1%
#742140000000
0!
0%
#742145000000
1!
1%
#742150000000
0!
0%
#742155000000
1!
1%
#742160000000
0!
0%
#742165000000
1!
1%
#742170000000
0!
0%
#742175000000
1!
1%
#742180000000
0!
0%
#742185000000
1!
1%
#742190000000
0!
0%
#742195000000
1!
1%
#742200000000
0!
0%
#742205000000
1!
1%
#742210000000
0!
0%
#742215000000
1!
1%
#742220000000
0!
0%
#742225000000
1!
1%
#742230000000
0!
0%
#742235000000
1!
1%
#742240000000
0!
0%
#742245000000
1!
1%
#742250000000
0!
0%
#742255000000
1!
1%
#742260000000
0!
0%
#742265000000
1!
1%
#742270000000
0!
0%
#742275000000
1!
1%
#742280000000
0!
0%
#742285000000
1!
1%
#742290000000
0!
0%
#742295000000
1!
1%
#742300000000
0!
0%
#742305000000
1!
1%
#742310000000
0!
0%
#742315000000
1!
1%
#742320000000
0!
0%
#742325000000
1!
1%
#742330000000
0!
0%
#742335000000
1!
1%
#742340000000
0!
0%
#742345000000
1!
1%
#742350000000
0!
0%
#742355000000
1!
1%
#742360000000
0!
0%
#742365000000
1!
1%
#742370000000
0!
0%
#742375000000
1!
1%
#742380000000
0!
0%
#742385000000
1!
1%
#742390000000
0!
0%
#742395000000
1!
1%
#742400000000
0!
0%
#742405000000
1!
1%
#742410000000
0!
0%
#742415000000
1!
1%
#742420000000
0!
0%
#742425000000
1!
1%
#742430000000
0!
0%
#742435000000
1!
1%
#742440000000
0!
0%
#742445000000
1!
1%
#742450000000
0!
0%
#742455000000
1!
1%
#742460000000
0!
0%
#742465000000
1!
1%
#742470000000
0!
0%
#742475000000
1!
1%
#742480000000
0!
0%
#742485000000
1!
1%
#742490000000
0!
0%
#742495000000
1!
1%
#742500000000
0!
0%
#742505000000
1!
1%
#742510000000
0!
0%
#742515000000
1!
1%
#742520000000
0!
0%
#742525000000
1!
1%
#742530000000
0!
0%
#742535000000
1!
1%
#742540000000
0!
0%
#742545000000
1!
1%
#742550000000
0!
0%
#742555000000
1!
1%
#742560000000
0!
0%
#742565000000
1!
1%
#742570000000
0!
0%
#742575000000
1!
1%
#742580000000
0!
0%
#742585000000
1!
1%
#742590000000
0!
0%
#742595000000
1!
1%
#742600000000
0!
0%
#742605000000
1!
1%
#742610000000
0!
0%
#742615000000
1!
1%
#742620000000
0!
0%
#742625000000
1!
1%
#742630000000
0!
0%
#742635000000
1!
1%
#742640000000
0!
0%
#742645000000
1!
1%
#742650000000
0!
0%
#742655000000
1!
1%
#742660000000
0!
0%
#742665000000
1!
1%
#742670000000
0!
0%
#742675000000
1!
1%
#742680000000
0!
0%
#742685000000
1!
1%
#742690000000
0!
0%
#742695000000
1!
1%
#742700000000
0!
0%
#742705000000
1!
1%
#742710000000
0!
0%
#742715000000
1!
1%
#742720000000
0!
0%
#742725000000
1!
1%
#742730000000
0!
0%
#742735000000
1!
1%
#742740000000
0!
0%
#742745000000
1!
1%
#742750000000
0!
0%
#742755000000
1!
1%
#742760000000
0!
0%
#742765000000
1!
1%
#742770000000
0!
0%
#742775000000
1!
1%
#742780000000
0!
0%
#742785000000
1!
1%
#742790000000
0!
0%
#742795000000
1!
1%
#742800000000
0!
0%
#742805000000
1!
1%
#742810000000
0!
0%
#742815000000
1!
1%
#742820000000
0!
0%
#742825000000
1!
1%
#742830000000
0!
0%
#742835000000
1!
1%
#742840000000
0!
0%
#742845000000
1!
1%
#742850000000
0!
0%
#742855000000
1!
1%
#742860000000
0!
0%
#742865000000
1!
1%
#742870000000
0!
0%
#742875000000
1!
1%
#742880000000
0!
0%
#742885000000
1!
1%
#742890000000
0!
0%
#742895000000
1!
1%
#742900000000
0!
0%
#742905000000
1!
1%
#742910000000
0!
0%
#742915000000
1!
1%
#742920000000
0!
0%
#742925000000
1!
1%
#742930000000
0!
0%
#742935000000
1!
1%
#742940000000
0!
0%
#742945000000
1!
1%
#742950000000
0!
0%
#742955000000
1!
1%
#742960000000
0!
0%
#742965000000
1!
1%
#742970000000
0!
0%
#742975000000
1!
1%
#742980000000
0!
0%
#742985000000
1!
1%
#742990000000
0!
0%
#742995000000
1!
1%
#743000000000
0!
0%
#743005000000
1!
1%
#743010000000
0!
0%
#743015000000
1!
1%
#743020000000
0!
0%
#743025000000
1!
1%
#743030000000
0!
0%
#743035000000
1!
1%
#743040000000
0!
0%
#743045000000
1!
1%
#743050000000
0!
0%
#743055000000
1!
1%
#743060000000
0!
0%
#743065000000
1!
1%
#743070000000
0!
0%
#743075000000
1!
1%
#743080000000
0!
0%
#743085000000
1!
1%
#743090000000
0!
0%
#743095000000
1!
1%
#743100000000
0!
0%
#743105000000
1!
1%
#743110000000
0!
0%
#743115000000
1!
1%
#743120000000
0!
0%
#743125000000
1!
1%
#743130000000
0!
0%
#743135000000
1!
1%
#743140000000
0!
0%
#743145000000
1!
1%
#743150000000
0!
0%
#743155000000
1!
1%
#743160000000
0!
0%
#743165000000
1!
1%
#743170000000
0!
0%
#743175000000
1!
1%
#743180000000
0!
0%
#743185000000
1!
1%
#743190000000
0!
0%
#743195000000
1!
1%
#743200000000
0!
0%
#743205000000
1!
1%
#743210000000
0!
0%
#743215000000
1!
1%
#743220000000
0!
0%
#743225000000
1!
1%
#743230000000
0!
0%
#743235000000
1!
1%
#743240000000
0!
0%
#743245000000
1!
1%
#743250000000
0!
0%
#743255000000
1!
1%
#743260000000
0!
0%
#743265000000
1!
1%
#743270000000
0!
0%
#743275000000
1!
1%
#743280000000
0!
0%
#743285000000
1!
1%
#743290000000
0!
0%
#743295000000
1!
1%
#743300000000
0!
0%
#743305000000
1!
1%
#743310000000
0!
0%
#743315000000
1!
1%
#743320000000
0!
0%
#743325000000
1!
1%
#743330000000
0!
0%
#743335000000
1!
1%
#743340000000
0!
0%
#743345000000
1!
1%
#743350000000
0!
0%
#743355000000
1!
1%
#743360000000
0!
0%
#743365000000
1!
1%
#743370000000
0!
0%
#743375000000
1!
1%
#743380000000
0!
0%
#743385000000
1!
1%
#743390000000
0!
0%
#743395000000
1!
1%
#743400000000
0!
0%
#743405000000
1!
1%
#743410000000
0!
0%
#743415000000
1!
1%
#743420000000
0!
0%
#743425000000
1!
1%
#743430000000
0!
0%
#743435000000
1!
1%
#743440000000
0!
0%
#743445000000
1!
1%
#743450000000
0!
0%
#743455000000
1!
1%
#743460000000
0!
0%
#743465000000
1!
1%
#743470000000
0!
0%
#743475000000
1!
1%
#743480000000
0!
0%
#743485000000
1!
1%
#743490000000
0!
0%
#743495000000
1!
1%
#743500000000
0!
0%
#743505000000
1!
1%
#743510000000
0!
0%
#743515000000
1!
1%
#743520000000
0!
0%
#743525000000
1!
1%
#743530000000
0!
0%
#743535000000
1!
1%
#743540000000
0!
0%
#743545000000
1!
1%
#743550000000
0!
0%
#743555000000
1!
1%
#743560000000
0!
0%
#743565000000
1!
1%
#743570000000
0!
0%
#743575000000
1!
1%
#743580000000
0!
0%
#743585000000
1!
1%
#743590000000
0!
0%
#743595000000
1!
1%
#743600000000
0!
0%
#743605000000
1!
1%
#743610000000
0!
0%
#743615000000
1!
1%
#743620000000
0!
0%
#743625000000
1!
1%
#743630000000
0!
0%
#743635000000
1!
1%
#743640000000
0!
0%
#743645000000
1!
1%
#743650000000
0!
0%
#743655000000
1!
1%
#743660000000
0!
0%
#743665000000
1!
1%
#743670000000
0!
0%
#743675000000
1!
1%
#743680000000
0!
0%
#743685000000
1!
1%
#743690000000
0!
0%
#743695000000
1!
1%
#743700000000
0!
0%
#743705000000
1!
1%
#743710000000
0!
0%
#743715000000
1!
1%
#743720000000
0!
0%
#743725000000
1!
1%
#743730000000
0!
0%
#743735000000
1!
1%
#743740000000
0!
0%
#743745000000
1!
1%
#743750000000
0!
0%
#743755000000
1!
1%
#743760000000
0!
0%
#743765000000
1!
1%
#743770000000
0!
0%
#743775000000
1!
1%
#743780000000
0!
0%
#743785000000
1!
1%
#743790000000
0!
0%
#743795000000
1!
1%
#743800000000
0!
0%
#743805000000
1!
1%
#743810000000
0!
0%
#743815000000
1!
1%
#743820000000
0!
0%
#743825000000
1!
1%
#743830000000
0!
0%
#743835000000
1!
1%
#743840000000
0!
0%
#743845000000
1!
1%
#743850000000
0!
0%
#743855000000
1!
1%
#743860000000
0!
0%
#743865000000
1!
1%
#743870000000
0!
0%
#743875000000
1!
1%
#743880000000
0!
0%
#743885000000
1!
1%
#743890000000
0!
0%
#743895000000
1!
1%
#743900000000
0!
0%
#743905000000
1!
1%
#743910000000
0!
0%
#743915000000
1!
1%
#743920000000
0!
0%
#743925000000
1!
1%
#743930000000
0!
0%
#743935000000
1!
1%
#743940000000
0!
0%
#743945000000
1!
1%
#743950000000
0!
0%
#743955000000
1!
1%
#743960000000
0!
0%
#743965000000
1!
1%
#743970000000
0!
0%
#743975000000
1!
1%
#743980000000
0!
0%
#743985000000
1!
1%
#743990000000
0!
0%
#743995000000
1!
1%
#744000000000
0!
0%
#744005000000
1!
1%
#744010000000
0!
0%
#744015000000
1!
1%
#744020000000
0!
0%
#744025000000
1!
1%
#744030000000
0!
0%
#744035000000
1!
1%
#744040000000
0!
0%
#744045000000
1!
1%
#744050000000
0!
0%
#744055000000
1!
1%
#744060000000
0!
0%
#744065000000
1!
1%
#744070000000
0!
0%
#744075000000
1!
1%
#744080000000
0!
0%
#744085000000
1!
1%
#744090000000
0!
0%
#744095000000
1!
1%
#744100000000
0!
0%
#744105000000
1!
1%
#744110000000
0!
0%
#744115000000
1!
1%
#744120000000
0!
0%
#744125000000
1!
1%
#744130000000
0!
0%
#744135000000
1!
1%
#744140000000
0!
0%
#744145000000
1!
1%
#744150000000
0!
0%
#744155000000
1!
1%
#744160000000
0!
0%
#744165000000
1!
1%
#744170000000
0!
0%
#744175000000
1!
1%
#744180000000
0!
0%
#744185000000
1!
1%
#744190000000
0!
0%
#744195000000
1!
1%
#744200000000
0!
0%
#744205000000
1!
1%
#744210000000
0!
0%
#744215000000
1!
1%
#744220000000
0!
0%
#744225000000
1!
1%
#744230000000
0!
0%
#744235000000
1!
1%
#744240000000
0!
0%
#744245000000
1!
1%
#744250000000
0!
0%
#744255000000
1!
1%
#744260000000
0!
0%
#744265000000
1!
1%
#744270000000
0!
0%
#744275000000
1!
1%
#744280000000
0!
0%
#744285000000
1!
1%
#744290000000
0!
0%
#744295000000
1!
1%
#744300000000
0!
0%
#744305000000
1!
1%
#744310000000
0!
0%
#744315000000
1!
1%
#744320000000
0!
0%
#744325000000
1!
1%
#744330000000
0!
0%
#744335000000
1!
1%
#744340000000
0!
0%
#744345000000
1!
1%
#744350000000
0!
0%
#744355000000
1!
1%
#744360000000
0!
0%
#744365000000
1!
1%
#744370000000
0!
0%
#744375000000
1!
1%
#744380000000
0!
0%
#744385000000
1!
1%
#744390000000
0!
0%
#744395000000
1!
1%
#744400000000
0!
0%
#744405000000
1!
1%
#744410000000
0!
0%
#744415000000
1!
1%
#744420000000
0!
0%
#744425000000
1!
1%
#744430000000
0!
0%
#744435000000
1!
1%
#744440000000
0!
0%
#744445000000
1!
1%
#744450000000
0!
0%
#744455000000
1!
1%
#744460000000
0!
0%
#744465000000
1!
1%
#744470000000
0!
0%
#744475000000
1!
1%
#744480000000
0!
0%
#744485000000
1!
1%
#744490000000
0!
0%
#744495000000
1!
1%
#744500000000
0!
0%
#744505000000
1!
1%
#744510000000
0!
0%
#744515000000
1!
1%
#744520000000
0!
0%
#744525000000
1!
1%
#744530000000
0!
0%
#744535000000
1!
1%
#744540000000
0!
0%
#744545000000
1!
1%
#744550000000
0!
0%
#744555000000
1!
1%
#744560000000
0!
0%
#744565000000
1!
1%
#744570000000
0!
0%
#744575000000
1!
1%
#744580000000
0!
0%
#744585000000
1!
1%
#744590000000
0!
0%
#744595000000
1!
1%
#744600000000
0!
0%
#744605000000
1!
1%
#744610000000
0!
0%
#744615000000
1!
1%
#744620000000
0!
0%
#744625000000
1!
1%
#744630000000
0!
0%
#744635000000
1!
1%
#744640000000
0!
0%
#744645000000
1!
1%
#744650000000
0!
0%
#744655000000
1!
1%
#744660000000
0!
0%
#744665000000
1!
1%
#744670000000
0!
0%
#744675000000
1!
1%
#744680000000
0!
0%
#744685000000
1!
1%
#744690000000
0!
0%
#744695000000
1!
1%
#744700000000
0!
0%
#744705000000
1!
1%
#744710000000
0!
0%
#744715000000
1!
1%
#744720000000
0!
0%
#744725000000
1!
1%
#744730000000
0!
0%
#744735000000
1!
1%
#744740000000
0!
0%
#744745000000
1!
1%
#744750000000
0!
0%
#744755000000
1!
1%
#744760000000
0!
0%
#744765000000
1!
1%
#744770000000
0!
0%
#744775000000
1!
1%
#744780000000
0!
0%
#744785000000
1!
1%
#744790000000
0!
0%
#744795000000
1!
1%
#744800000000
0!
0%
#744805000000
1!
1%
#744810000000
0!
0%
#744815000000
1!
1%
#744820000000
0!
0%
#744825000000
1!
1%
#744830000000
0!
0%
#744835000000
1!
1%
#744840000000
0!
0%
#744845000000
1!
1%
#744850000000
0!
0%
#744855000000
1!
1%
#744860000000
0!
0%
#744865000000
1!
1%
#744870000000
0!
0%
#744875000000
1!
1%
#744880000000
0!
0%
#744885000000
1!
1%
#744890000000
0!
0%
#744895000000
1!
1%
#744900000000
0!
0%
#744905000000
1!
1%
#744910000000
0!
0%
#744915000000
1!
1%
#744920000000
0!
0%
#744925000000
1!
1%
#744930000000
0!
0%
#744935000000
1!
1%
#744940000000
0!
0%
#744945000000
1!
1%
#744950000000
0!
0%
#744955000000
1!
1%
#744960000000
0!
0%
#744965000000
1!
1%
#744970000000
0!
0%
#744975000000
1!
1%
#744980000000
0!
0%
#744985000000
1!
1%
#744990000000
0!
0%
#744995000000
1!
1%
#745000000000
0!
0%
#745005000000
1!
1%
#745010000000
0!
0%
#745015000000
1!
1%
#745020000000
0!
0%
#745025000000
1!
1%
#745030000000
0!
0%
#745035000000
1!
1%
#745040000000
0!
0%
#745045000000
1!
1%
#745050000000
0!
0%
#745055000000
1!
1%
#745060000000
0!
0%
#745065000000
1!
1%
#745070000000
0!
0%
#745075000000
1!
1%
#745080000000
0!
0%
#745085000000
1!
1%
#745090000000
0!
0%
#745095000000
1!
1%
#745100000000
0!
0%
#745105000000
1!
1%
#745110000000
0!
0%
#745115000000
1!
1%
#745120000000
0!
0%
#745125000000
1!
1%
#745130000000
0!
0%
#745135000000
1!
1%
#745140000000
0!
0%
#745145000000
1!
1%
#745150000000
0!
0%
#745155000000
1!
1%
#745160000000
0!
0%
#745165000000
1!
1%
#745170000000
0!
0%
#745175000000
1!
1%
#745180000000
0!
0%
#745185000000
1!
1%
#745190000000
0!
0%
#745195000000
1!
1%
#745200000000
0!
0%
#745205000000
1!
1%
#745210000000
0!
0%
#745215000000
1!
1%
#745220000000
0!
0%
#745225000000
1!
1%
#745230000000
0!
0%
#745235000000
1!
1%
#745240000000
0!
0%
#745245000000
1!
1%
#745250000000
0!
0%
#745255000000
1!
1%
#745260000000
0!
0%
#745265000000
1!
1%
#745270000000
0!
0%
#745275000000
1!
1%
#745280000000
0!
0%
#745285000000
1!
1%
#745290000000
0!
0%
#745295000000
1!
1%
#745300000000
0!
0%
#745305000000
1!
1%
#745310000000
0!
0%
#745315000000
1!
1%
#745320000000
0!
0%
#745325000000
1!
1%
#745330000000
0!
0%
#745335000000
1!
1%
#745340000000
0!
0%
#745345000000
1!
1%
#745350000000
0!
0%
#745355000000
1!
1%
#745360000000
0!
0%
#745365000000
1!
1%
#745370000000
0!
0%
#745375000000
1!
1%
#745380000000
0!
0%
#745385000000
1!
1%
#745390000000
0!
0%
#745395000000
1!
1%
#745400000000
0!
0%
#745405000000
1!
1%
#745410000000
0!
0%
#745415000000
1!
1%
#745420000000
0!
0%
#745425000000
1!
1%
#745430000000
0!
0%
#745435000000
1!
1%
#745440000000
0!
0%
#745445000000
1!
1%
#745450000000
0!
0%
#745455000000
1!
1%
#745460000000
0!
0%
#745465000000
1!
1%
#745470000000
0!
0%
#745475000000
1!
1%
#745480000000
0!
0%
#745485000000
1!
1%
#745490000000
0!
0%
#745495000000
1!
1%
#745500000000
0!
0%
#745505000000
1!
1%
#745510000000
0!
0%
#745515000000
1!
1%
#745520000000
0!
0%
#745525000000
1!
1%
#745530000000
0!
0%
#745535000000
1!
1%
#745540000000
0!
0%
#745545000000
1!
1%
#745550000000
0!
0%
#745555000000
1!
1%
#745560000000
0!
0%
#745565000000
1!
1%
#745570000000
0!
0%
#745575000000
1!
1%
#745580000000
0!
0%
#745585000000
1!
1%
#745590000000
0!
0%
#745595000000
1!
1%
#745600000000
0!
0%
#745605000000
1!
1%
#745610000000
0!
0%
#745615000000
1!
1%
#745620000000
0!
0%
#745625000000
1!
1%
#745630000000
0!
0%
#745635000000
1!
1%
#745640000000
0!
0%
#745645000000
1!
1%
#745650000000
0!
0%
#745655000000
1!
1%
#745660000000
0!
0%
#745665000000
1!
1%
#745670000000
0!
0%
#745675000000
1!
1%
#745680000000
0!
0%
#745685000000
1!
1%
#745690000000
0!
0%
#745695000000
1!
1%
#745700000000
0!
0%
#745705000000
1!
1%
#745710000000
0!
0%
#745715000000
1!
1%
#745720000000
0!
0%
#745725000000
1!
1%
#745730000000
0!
0%
#745735000000
1!
1%
#745740000000
0!
0%
#745745000000
1!
1%
#745750000000
0!
0%
#745755000000
1!
1%
#745760000000
0!
0%
#745765000000
1!
1%
#745770000000
0!
0%
#745775000000
1!
1%
#745780000000
0!
0%
#745785000000
1!
1%
#745790000000
0!
0%
#745795000000
1!
1%
#745800000000
0!
0%
#745805000000
1!
1%
#745810000000
0!
0%
#745815000000
1!
1%
#745820000000
0!
0%
#745825000000
1!
1%
#745830000000
0!
0%
#745835000000
1!
1%
#745840000000
0!
0%
#745845000000
1!
1%
#745850000000
0!
0%
#745855000000
1!
1%
#745860000000
0!
0%
#745865000000
1!
1%
#745870000000
0!
0%
#745875000000
1!
1%
#745880000000
0!
0%
#745885000000
1!
1%
#745890000000
0!
0%
#745895000000
1!
1%
#745900000000
0!
0%
#745905000000
1!
1%
#745910000000
0!
0%
#745915000000
1!
1%
#745920000000
0!
0%
#745925000000
1!
1%
#745930000000
0!
0%
#745935000000
1!
1%
#745940000000
0!
0%
#745945000000
1!
1%
#745950000000
0!
0%
#745955000000
1!
1%
#745960000000
0!
0%
#745965000000
1!
1%
#745970000000
0!
0%
#745975000000
1!
1%
#745980000000
0!
0%
#745985000000
1!
1%
#745990000000
0!
0%
#745995000000
1!
1%
#746000000000
0!
0%
#746005000000
1!
1%
#746010000000
0!
0%
#746015000000
1!
1%
#746020000000
0!
0%
#746025000000
1!
1%
#746030000000
0!
0%
#746035000000
1!
1%
#746040000000
0!
0%
#746045000000
1!
1%
#746050000000
0!
0%
#746055000000
1!
1%
#746060000000
0!
0%
#746065000000
1!
1%
#746070000000
0!
0%
#746075000000
1!
1%
#746080000000
0!
0%
#746085000000
1!
1%
#746090000000
0!
0%
#746095000000
1!
1%
#746100000000
0!
0%
#746105000000
1!
1%
#746110000000
0!
0%
#746115000000
1!
1%
#746120000000
0!
0%
#746125000000
1!
1%
#746130000000
0!
0%
#746135000000
1!
1%
#746140000000
0!
0%
#746145000000
1!
1%
#746150000000
0!
0%
#746155000000
1!
1%
#746160000000
0!
0%
#746165000000
1!
1%
#746170000000
0!
0%
#746175000000
1!
1%
#746180000000
0!
0%
#746185000000
1!
1%
#746190000000
0!
0%
#746195000000
1!
1%
#746200000000
0!
0%
#746205000000
1!
1%
#746210000000
0!
0%
#746215000000
1!
1%
#746220000000
0!
0%
#746225000000
1!
1%
#746230000000
0!
0%
#746235000000
1!
1%
#746240000000
0!
0%
#746245000000
1!
1%
#746250000000
0!
0%
#746255000000
1!
1%
#746260000000
0!
0%
#746265000000
1!
1%
#746270000000
0!
0%
#746275000000
1!
1%
#746280000000
0!
0%
#746285000000
1!
1%
#746290000000
0!
0%
#746295000000
1!
1%
#746300000000
0!
0%
#746305000000
1!
1%
#746310000000
0!
0%
#746315000000
1!
1%
#746320000000
0!
0%
#746325000000
1!
1%
#746330000000
0!
0%
#746335000000
1!
1%
#746340000000
0!
0%
#746345000000
1!
1%
#746350000000
0!
0%
#746355000000
1!
1%
#746360000000
0!
0%
#746365000000
1!
1%
#746370000000
0!
0%
#746375000000
1!
1%
#746380000000
0!
0%
#746385000000
1!
1%
#746390000000
0!
0%
#746395000000
1!
1%
#746400000000
0!
0%
#746405000000
1!
1%
#746410000000
0!
0%
#746415000000
1!
1%
#746420000000
0!
0%
#746425000000
1!
1%
#746430000000
0!
0%
#746435000000
1!
1%
#746440000000
0!
0%
#746445000000
1!
1%
#746450000000
0!
0%
#746455000000
1!
1%
#746460000000
0!
0%
#746465000000
1!
1%
#746470000000
0!
0%
#746475000000
1!
1%
#746480000000
0!
0%
#746485000000
1!
1%
#746490000000
0!
0%
#746495000000
1!
1%
#746500000000
0!
0%
#746505000000
1!
1%
#746510000000
0!
0%
#746515000000
1!
1%
#746520000000
0!
0%
#746525000000
1!
1%
#746530000000
0!
0%
#746535000000
1!
1%
#746540000000
0!
0%
#746545000000
1!
1%
#746550000000
0!
0%
#746555000000
1!
1%
#746560000000
0!
0%
#746565000000
1!
1%
#746570000000
0!
0%
#746575000000
1!
1%
#746580000000
0!
0%
#746585000000
1!
1%
#746590000000
0!
0%
#746595000000
1!
1%
#746600000000
0!
0%
#746605000000
1!
1%
#746610000000
0!
0%
#746615000000
1!
1%
#746620000000
0!
0%
#746625000000
1!
1%
#746630000000
0!
0%
#746635000000
1!
1%
#746640000000
0!
0%
#746645000000
1!
1%
#746650000000
0!
0%
#746655000000
1!
1%
#746660000000
0!
0%
#746665000000
1!
1%
#746670000000
0!
0%
#746675000000
1!
1%
#746680000000
0!
0%
#746685000000
1!
1%
#746690000000
0!
0%
#746695000000
1!
1%
#746700000000
0!
0%
#746705000000
1!
1%
#746710000000
0!
0%
#746715000000
1!
1%
#746720000000
0!
0%
#746725000000
1!
1%
#746730000000
0!
0%
#746735000000
1!
1%
#746740000000
0!
0%
#746745000000
1!
1%
#746750000000
0!
0%
#746755000000
1!
1%
#746760000000
0!
0%
#746765000000
1!
1%
#746770000000
0!
0%
#746775000000
1!
1%
#746780000000
0!
0%
#746785000000
1!
1%
#746790000000
0!
0%
#746795000000
1!
1%
#746800000000
0!
0%
#746805000000
1!
1%
#746810000000
0!
0%
#746815000000
1!
1%
#746820000000
0!
0%
#746825000000
1!
1%
#746830000000
0!
0%
#746835000000
1!
1%
#746840000000
0!
0%
#746845000000
1!
1%
#746850000000
0!
0%
#746855000000
1!
1%
#746860000000
0!
0%
#746865000000
1!
1%
#746870000000
0!
0%
#746875000000
1!
1%
#746880000000
0!
0%
#746885000000
1!
1%
#746890000000
0!
0%
#746895000000
1!
1%
#746900000000
0!
0%
#746905000000
1!
1%
#746910000000
0!
0%
#746915000000
1!
1%
#746920000000
0!
0%
#746925000000
1!
1%
#746930000000
0!
0%
#746935000000
1!
1%
#746940000000
0!
0%
#746945000000
1!
1%
#746950000000
0!
0%
#746955000000
1!
1%
#746960000000
0!
0%
#746965000000
1!
1%
#746970000000
0!
0%
#746975000000
1!
1%
#746980000000
0!
0%
#746985000000
1!
1%
#746990000000
0!
0%
#746995000000
1!
1%
#747000000000
0!
0%
#747005000000
1!
1%
#747010000000
0!
0%
#747015000000
1!
1%
#747020000000
0!
0%
#747025000000
1!
1%
#747030000000
0!
0%
#747035000000
1!
1%
#747040000000
0!
0%
#747045000000
1!
1%
#747050000000
0!
0%
#747055000000
1!
1%
#747060000000
0!
0%
#747065000000
1!
1%
#747070000000
0!
0%
#747075000000
1!
1%
#747080000000
0!
0%
#747085000000
1!
1%
#747090000000
0!
0%
#747095000000
1!
1%
#747100000000
0!
0%
#747105000000
1!
1%
#747110000000
0!
0%
#747115000000
1!
1%
#747120000000
0!
0%
#747125000000
1!
1%
#747130000000
0!
0%
#747135000000
1!
1%
#747140000000
0!
0%
#747145000000
1!
1%
#747150000000
0!
0%
#747155000000
1!
1%
#747160000000
0!
0%
#747165000000
1!
1%
#747170000000
0!
0%
#747175000000
1!
1%
#747180000000
0!
0%
#747185000000
1!
1%
#747190000000
0!
0%
#747195000000
1!
1%
#747200000000
0!
0%
#747205000000
1!
1%
#747210000000
0!
0%
#747215000000
1!
1%
#747220000000
0!
0%
#747225000000
1!
1%
#747230000000
0!
0%
#747235000000
1!
1%
#747240000000
0!
0%
#747245000000
1!
1%
#747250000000
0!
0%
#747255000000
1!
1%
#747260000000
0!
0%
#747265000000
1!
1%
#747270000000
0!
0%
#747275000000
1!
1%
#747280000000
0!
0%
#747285000000
1!
1%
#747290000000
0!
0%
#747295000000
1!
1%
#747300000000
0!
0%
#747305000000
1!
1%
#747310000000
0!
0%
#747315000000
1!
1%
#747320000000
0!
0%
#747325000000
1!
1%
#747330000000
0!
0%
#747335000000
1!
1%
#747340000000
0!
0%
#747345000000
1!
1%
#747350000000
0!
0%
#747355000000
1!
1%
#747360000000
0!
0%
#747365000000
1!
1%
#747370000000
0!
0%
#747375000000
1!
1%
#747380000000
0!
0%
#747385000000
1!
1%
#747390000000
0!
0%
#747395000000
1!
1%
#747400000000
0!
0%
#747405000000
1!
1%
#747410000000
0!
0%
#747415000000
1!
1%
#747420000000
0!
0%
#747425000000
1!
1%
#747430000000
0!
0%
#747435000000
1!
1%
#747440000000
0!
0%
#747445000000
1!
1%
#747450000000
0!
0%
#747455000000
1!
1%
#747460000000
0!
0%
#747465000000
1!
1%
#747470000000
0!
0%
#747475000000
1!
1%
#747480000000
0!
0%
#747485000000
1!
1%
#747490000000
0!
0%
#747495000000
1!
1%
#747500000000
0!
0%
#747505000000
1!
1%
#747510000000
0!
0%
#747515000000
1!
1%
#747520000000
0!
0%
#747525000000
1!
1%
#747530000000
0!
0%
#747535000000
1!
1%
#747540000000
0!
0%
#747545000000
1!
1%
#747550000000
0!
0%
#747555000000
1!
1%
#747560000000
0!
0%
#747565000000
1!
1%
#747570000000
0!
0%
#747575000000
1!
1%
#747580000000
0!
0%
#747585000000
1!
1%
#747590000000
0!
0%
#747595000000
1!
1%
#747600000000
0!
0%
#747605000000
1!
1%
#747610000000
0!
0%
#747615000000
1!
1%
#747620000000
0!
0%
#747625000000
1!
1%
#747630000000
0!
0%
#747635000000
1!
1%
#747640000000
0!
0%
#747645000000
1!
1%
#747650000000
0!
0%
#747655000000
1!
1%
#747660000000
0!
0%
#747665000000
1!
1%
#747670000000
0!
0%
#747675000000
1!
1%
#747680000000
0!
0%
#747685000000
1!
1%
#747690000000
0!
0%
#747695000000
1!
1%
#747700000000
0!
0%
#747705000000
1!
1%
#747710000000
0!
0%
#747715000000
1!
1%
#747720000000
0!
0%
#747725000000
1!
1%
#747730000000
0!
0%
#747735000000
1!
1%
#747740000000
0!
0%
#747745000000
1!
1%
#747750000000
0!
0%
#747755000000
1!
1%
#747760000000
0!
0%
#747765000000
1!
1%
#747770000000
0!
0%
#747775000000
1!
1%
#747780000000
0!
0%
#747785000000
1!
1%
#747790000000
0!
0%
#747795000000
1!
1%
#747800000000
0!
0%
#747805000000
1!
1%
#747810000000
0!
0%
#747815000000
1!
1%
#747820000000
0!
0%
#747825000000
1!
1%
#747830000000
0!
0%
#747835000000
1!
1%
#747840000000
0!
0%
#747845000000
1!
1%
#747850000000
0!
0%
#747855000000
1!
1%
#747860000000
0!
0%
#747865000000
1!
1%
#747870000000
0!
0%
#747875000000
1!
1%
#747880000000
0!
0%
#747885000000
1!
1%
#747890000000
0!
0%
#747895000000
1!
1%
#747900000000
0!
0%
#747905000000
1!
1%
#747910000000
0!
0%
#747915000000
1!
1%
#747920000000
0!
0%
#747925000000
1!
1%
#747930000000
0!
0%
#747935000000
1!
1%
#747940000000
0!
0%
#747945000000
1!
1%
#747950000000
0!
0%
#747955000000
1!
1%
#747960000000
0!
0%
#747965000000
1!
1%
#747970000000
0!
0%
#747975000000
1!
1%
#747980000000
0!
0%
#747985000000
1!
1%
#747990000000
0!
0%
#747995000000
1!
1%
#748000000000
0!
0%
#748005000000
1!
1%
#748010000000
0!
0%
#748015000000
1!
1%
#748020000000
0!
0%
#748025000000
1!
1%
#748030000000
0!
0%
#748035000000
1!
1%
#748040000000
0!
0%
#748045000000
1!
1%
#748050000000
0!
0%
#748055000000
1!
1%
#748060000000
0!
0%
#748065000000
1!
1%
#748070000000
0!
0%
#748075000000
1!
1%
#748080000000
0!
0%
#748085000000
1!
1%
#748090000000
0!
0%
#748095000000
1!
1%
#748100000000
0!
0%
#748105000000
1!
1%
#748110000000
0!
0%
#748115000000
1!
1%
#748120000000
0!
0%
#748125000000
1!
1%
#748130000000
0!
0%
#748135000000
1!
1%
#748140000000
0!
0%
#748145000000
1!
1%
#748150000000
0!
0%
#748155000000
1!
1%
#748160000000
0!
0%
#748165000000
1!
1%
#748170000000
0!
0%
#748175000000
1!
1%
#748180000000
0!
0%
#748185000000
1!
1%
#748190000000
0!
0%
#748195000000
1!
1%
#748200000000
0!
0%
#748205000000
1!
1%
#748210000000
0!
0%
#748215000000
1!
1%
#748220000000
0!
0%
#748225000000
1!
1%
#748230000000
0!
0%
#748235000000
1!
1%
#748240000000
0!
0%
#748245000000
1!
1%
#748250000000
0!
0%
#748255000000
1!
1%
#748260000000
0!
0%
#748265000000
1!
1%
#748270000000
0!
0%
#748275000000
1!
1%
#748280000000
0!
0%
#748285000000
1!
1%
#748290000000
0!
0%
#748295000000
1!
1%
#748300000000
0!
0%
#748305000000
1!
1%
#748310000000
0!
0%
#748315000000
1!
1%
#748320000000
0!
0%
#748325000000
1!
1%
#748330000000
0!
0%
#748335000000
1!
1%
#748340000000
0!
0%
#748345000000
1!
1%
#748350000000
0!
0%
#748355000000
1!
1%
#748360000000
0!
0%
#748365000000
1!
1%
#748370000000
0!
0%
#748375000000
1!
1%
#748380000000
0!
0%
#748385000000
1!
1%
#748390000000
0!
0%
#748395000000
1!
1%
#748400000000
0!
0%
#748405000000
1!
1%
#748410000000
0!
0%
#748415000000
1!
1%
#748420000000
0!
0%
#748425000000
1!
1%
#748430000000
0!
0%
#748435000000
1!
1%
#748440000000
0!
0%
#748445000000
1!
1%
#748450000000
0!
0%
#748455000000
1!
1%
#748460000000
0!
0%
#748465000000
1!
1%
#748470000000
0!
0%
#748475000000
1!
1%
#748480000000
0!
0%
#748485000000
1!
1%
#748490000000
0!
0%
#748495000000
1!
1%
#748500000000
0!
0%
#748505000000
1!
1%
#748510000000
0!
0%
#748515000000
1!
1%
#748520000000
0!
0%
#748525000000
1!
1%
#748530000000
0!
0%
#748535000000
1!
1%
#748540000000
0!
0%
#748545000000
1!
1%
#748550000000
0!
0%
#748555000000
1!
1%
#748560000000
0!
0%
#748565000000
1!
1%
#748570000000
0!
0%
#748575000000
1!
1%
#748580000000
0!
0%
#748585000000
1!
1%
#748590000000
0!
0%
#748595000000
1!
1%
#748600000000
0!
0%
#748605000000
1!
1%
#748610000000
0!
0%
#748615000000
1!
1%
#748620000000
0!
0%
#748625000000
1!
1%
#748630000000
0!
0%
#748635000000
1!
1%
#748640000000
0!
0%
#748645000000
1!
1%
#748650000000
0!
0%
#748655000000
1!
1%
#748660000000
0!
0%
#748665000000
1!
1%
#748670000000
0!
0%
#748675000000
1!
1%
#748680000000
0!
0%
#748685000000
1!
1%
#748690000000
0!
0%
#748695000000
1!
1%
#748700000000
0!
0%
#748705000000
1!
1%
#748710000000
0!
0%
#748715000000
1!
1%
#748720000000
0!
0%
#748725000000
1!
1%
#748730000000
0!
0%
#748735000000
1!
1%
#748740000000
0!
0%
#748745000000
1!
1%
#748750000000
0!
0%
#748755000000
1!
1%
#748760000000
0!
0%
#748765000000
1!
1%
#748770000000
0!
0%
#748775000000
1!
1%
#748780000000
0!
0%
#748785000000
1!
1%
#748790000000
0!
0%
#748795000000
1!
1%
#748800000000
0!
0%
#748805000000
1!
1%
#748810000000
0!
0%
#748815000000
1!
1%
#748820000000
0!
0%
#748825000000
1!
1%
#748830000000
0!
0%
#748835000000
1!
1%
#748840000000
0!
0%
#748845000000
1!
1%
#748850000000
0!
0%
#748855000000
1!
1%
#748860000000
0!
0%
#748865000000
1!
1%
#748870000000
0!
0%
#748875000000
1!
1%
#748880000000
0!
0%
#748885000000
1!
1%
#748890000000
0!
0%
#748895000000
1!
1%
#748900000000
0!
0%
#748905000000
1!
1%
#748910000000
0!
0%
#748915000000
1!
1%
#748920000000
0!
0%
#748925000000
1!
1%
#748930000000
0!
0%
#748935000000
1!
1%
#748940000000
0!
0%
#748945000000
1!
1%
#748950000000
0!
0%
#748955000000
1!
1%
#748960000000
0!
0%
#748965000000
1!
1%
#748970000000
0!
0%
#748975000000
1!
1%
#748980000000
0!
0%
#748985000000
1!
1%
#748990000000
0!
0%
#748995000000
1!
1%
#749000000000
0!
0%
#749005000000
1!
1%
#749010000000
0!
0%
#749015000000
1!
1%
#749020000000
0!
0%
#749025000000
1!
1%
#749030000000
0!
0%
#749035000000
1!
1%
#749040000000
0!
0%
#749045000000
1!
1%
#749050000000
0!
0%
#749055000000
1!
1%
#749060000000
0!
0%
#749065000000
1!
1%
#749070000000
0!
0%
#749075000000
1!
1%
#749080000000
0!
0%
#749085000000
1!
1%
#749090000000
0!
0%
#749095000000
1!
1%
#749100000000
0!
0%
#749105000000
1!
1%
#749110000000
0!
0%
#749115000000
1!
1%
#749120000000
0!
0%
#749125000000
1!
1%
#749130000000
0!
0%
#749135000000
1!
1%
#749140000000
0!
0%
#749145000000
1!
1%
#749150000000
0!
0%
#749155000000
1!
1%
#749160000000
0!
0%
#749165000000
1!
1%
#749170000000
0!
0%
#749175000000
1!
1%
#749180000000
0!
0%
#749185000000
1!
1%
#749190000000
0!
0%
#749195000000
1!
1%
#749200000000
0!
0%
#749205000000
1!
1%
#749210000000
0!
0%
#749215000000
1!
1%
#749220000000
0!
0%
#749225000000
1!
1%
#749230000000
0!
0%
#749235000000
1!
1%
#749240000000
0!
0%
#749245000000
1!
1%
#749250000000
0!
0%
#749255000000
1!
1%
#749260000000
0!
0%
#749265000000
1!
1%
#749270000000
0!
0%
#749275000000
1!
1%
#749280000000
0!
0%
#749285000000
1!
1%
#749290000000
0!
0%
#749295000000
1!
1%
#749300000000
0!
0%
#749305000000
1!
1%
#749310000000
0!
0%
#749315000000
1!
1%
#749320000000
0!
0%
#749325000000
1!
1%
#749330000000
0!
0%
#749335000000
1!
1%
#749340000000
0!
0%
#749345000000
1!
1%
#749350000000
0!
0%
#749355000000
1!
1%
#749360000000
0!
0%
#749365000000
1!
1%
#749370000000
0!
0%
#749375000000
1!
1%
#749380000000
0!
0%
#749385000000
1!
1%
#749390000000
0!
0%
#749395000000
1!
1%
#749400000000
0!
0%
#749405000000
1!
1%
#749410000000
0!
0%
#749415000000
1!
1%
#749420000000
0!
0%
#749425000000
1!
1%
#749430000000
0!
0%
#749435000000
1!
1%
#749440000000
0!
0%
#749445000000
1!
1%
#749450000000
0!
0%
#749455000000
1!
1%
#749460000000
0!
0%
#749465000000
1!
1%
#749470000000
0!
0%
#749475000000
1!
1%
#749480000000
0!
0%
#749485000000
1!
1%
#749490000000
0!
0%
#749495000000
1!
1%
#749500000000
0!
0%
#749505000000
1!
1%
#749510000000
0!
0%
#749515000000
1!
1%
#749520000000
0!
0%
#749525000000
1!
1%
#749530000000
0!
0%
#749535000000
1!
1%
#749540000000
0!
0%
#749545000000
1!
1%
#749550000000
0!
0%
#749555000000
1!
1%
#749560000000
0!
0%
#749565000000
1!
1%
#749570000000
0!
0%
#749575000000
1!
1%
#749580000000
0!
0%
#749585000000
1!
1%
#749590000000
0!
0%
#749595000000
1!
1%
#749600000000
0!
0%
#749605000000
1!
1%
#749610000000
0!
0%
#749615000000
1!
1%
#749620000000
0!
0%
#749625000000
1!
1%
#749630000000
0!
0%
#749635000000
1!
1%
#749640000000
0!
0%
#749645000000
1!
1%
#749650000000
0!
0%
#749655000000
1!
1%
#749660000000
0!
0%
#749665000000
1!
1%
#749670000000
0!
0%
#749675000000
1!
1%
#749680000000
0!
0%
#749685000000
1!
1%
#749690000000
0!
0%
#749695000000
1!
1%
#749700000000
0!
0%
#749705000000
1!
1%
#749710000000
0!
0%
#749715000000
1!
1%
#749720000000
0!
0%
#749725000000
1!
1%
#749730000000
0!
0%
#749735000000
1!
1%
#749740000000
0!
0%
#749745000000
1!
1%
#749750000000
0!
0%
#749755000000
1!
1%
#749760000000
0!
0%
#749765000000
1!
1%
#749770000000
0!
0%
#749775000000
1!
1%
#749780000000
0!
0%
#749785000000
1!
1%
#749790000000
0!
0%
#749795000000
1!
1%
#749800000000
0!
0%
#749805000000
1!
1%
#749810000000
0!
0%
#749815000000
1!
1%
#749820000000
0!
0%
#749825000000
1!
1%
#749830000000
0!
0%
#749835000000
1!
1%
#749840000000
0!
0%
#749845000000
1!
1%
#749850000000
0!
0%
#749855000000
1!
1%
#749860000000
0!
0%
#749865000000
1!
1%
#749870000000
0!
0%
#749875000000
1!
1%
#749880000000
0!
0%
#749885000000
1!
1%
#749890000000
0!
0%
#749895000000
1!
1%
#749900000000
0!
0%
#749905000000
1!
1%
#749910000000
0!
0%
#749915000000
1!
1%
#749920000000
0!
0%
#749925000000
1!
1%
#749930000000
0!
0%
#749935000000
1!
1%
#749940000000
0!
0%
#749945000000
1!
1%
#749950000000
0!
0%
#749955000000
1!
1%
#749960000000
0!
0%
#749965000000
1!
1%
#749970000000
0!
0%
#749975000000
1!
1%
#749980000000
0!
0%
#749985000000
1!
1%
#749990000000
0!
0%
#749995000000
1!
1%
#750000000000
0!
0%
#750005000000
1!
1%
#750010000000
0!
0%
#750015000000
1!
1%
#750020000000
0!
0%
#750025000000
1!
1%
#750030000000
0!
0%
#750035000000
1!
1%
#750040000000
0!
0%
#750045000000
1!
1%
#750050000000
0!
0%
#750055000000
1!
1%
#750060000000
0!
0%
#750065000000
1!
1%
#750070000000
0!
0%
#750075000000
1!
1%
#750080000000
0!
0%
#750085000000
1!
1%
#750090000000
0!
0%
#750095000000
1!
1%
#750100000000
0!
0%
#750105000000
1!
1%
#750110000000
0!
0%
#750115000000
1!
1%
#750120000000
0!
0%
#750125000000
1!
1%
#750130000000
0!
0%
#750135000000
1!
1%
#750140000000
0!
0%
#750145000000
1!
1%
#750150000000
0!
0%
#750155000000
1!
1%
#750160000000
0!
0%
#750165000000
1!
1%
#750170000000
0!
0%
#750175000000
1!
1%
#750180000000
0!
0%
#750185000000
1!
1%
#750190000000
0!
0%
#750195000000
1!
1%
#750200000000
0!
0%
#750205000000
1!
1%
#750210000000
0!
0%
#750215000000
1!
1%
#750220000000
0!
0%
#750225000000
1!
1%
#750230000000
0!
0%
#750235000000
1!
1%
#750240000000
0!
0%
#750245000000
1!
1%
#750250000000
0!
0%
#750255000000
1!
1%
#750260000000
0!
0%
#750265000000
1!
1%
#750270000000
0!
0%
#750275000000
1!
1%
#750280000000
0!
0%
#750285000000
1!
1%
#750290000000
0!
0%
#750295000000
1!
1%
#750300000000
0!
0%
#750305000000
1!
1%
#750310000000
0!
0%
#750315000000
1!
1%
#750320000000
0!
0%
#750325000000
1!
1%
#750330000000
0!
0%
#750335000000
1!
1%
#750340000000
0!
0%
#750345000000
1!
1%
#750350000000
0!
0%
#750355000000
1!
1%
#750360000000
0!
0%
#750365000000
1!
1%
#750370000000
0!
0%
#750375000000
1!
1%
#750380000000
0!
0%
#750385000000
1!
1%
#750390000000
0!
0%
#750395000000
1!
1%
#750400000000
0!
0%
#750405000000
1!
1%
#750410000000
0!
0%
#750415000000
1!
1%
#750420000000
0!
0%
#750425000000
1!
1%
#750430000000
0!
0%
#750435000000
1!
1%
#750440000000
0!
0%
#750445000000
1!
1%
#750450000000
0!
0%
#750455000000
1!
1%
#750460000000
0!
0%
#750465000000
1!
1%
#750470000000
0!
0%
#750475000000
1!
1%
#750480000000
0!
0%
#750485000000
1!
1%
#750490000000
0!
0%
#750495000000
1!
1%
#750500000000
0!
0%
#750505000000
1!
1%
#750510000000
0!
0%
#750515000000
1!
1%
#750520000000
0!
0%
#750525000000
1!
1%
#750530000000
0!
0%
#750535000000
1!
1%
#750540000000
0!
0%
#750545000000
1!
1%
#750550000000
0!
0%
#750555000000
1!
1%
#750560000000
0!
0%
#750565000000
1!
1%
#750570000000
0!
0%
#750575000000
1!
1%
#750580000000
0!
0%
#750585000000
1!
1%
#750590000000
0!
0%
#750595000000
1!
1%
#750600000000
0!
0%
#750605000000
1!
1%
#750610000000
0!
0%
#750615000000
1!
1%
#750620000000
0!
0%
#750625000000
1!
1%
#750630000000
0!
0%
#750635000000
1!
1%
#750640000000
0!
0%
#750645000000
1!
1%
#750650000000
0!
0%
#750655000000
1!
1%
#750660000000
0!
0%
#750665000000
1!
1%
#750670000000
0!
0%
#750675000000
1!
1%
#750680000000
0!
0%
#750685000000
1!
1%
#750690000000
0!
0%
#750695000000
1!
1%
#750700000000
0!
0%
#750705000000
1!
1%
#750710000000
0!
0%
#750715000000
1!
1%
#750720000000
0!
0%
#750725000000
1!
1%
#750730000000
0!
0%
#750735000000
1!
1%
#750740000000
0!
0%
#750745000000
1!
1%
#750750000000
0!
0%
#750755000000
1!
1%
#750760000000
0!
0%
#750765000000
1!
1%
#750770000000
0!
0%
#750775000000
1!
1%
#750780000000
0!
0%
#750785000000
1!
1%
#750790000000
0!
0%
#750795000000
1!
1%
#750800000000
0!
0%
#750805000000
1!
1%
#750810000000
0!
0%
#750815000000
1!
1%
#750820000000
0!
0%
#750825000000
1!
1%
#750830000000
0!
0%
#750835000000
1!
1%
#750840000000
0!
0%
#750845000000
1!
1%
#750850000000
0!
0%
#750855000000
1!
1%
#750860000000
0!
0%
#750865000000
1!
1%
#750870000000
0!
0%
#750875000000
1!
1%
#750880000000
0!
0%
#750885000000
1!
1%
#750890000000
0!
0%
#750895000000
1!
1%
#750900000000
0!
0%
#750905000000
1!
1%
#750910000000
0!
0%
#750915000000
1!
1%
#750920000000
0!
0%
#750925000000
1!
1%
#750930000000
0!
0%
#750935000000
1!
1%
#750940000000
0!
0%
#750945000000
1!
1%
#750950000000
0!
0%
#750955000000
1!
1%
#750960000000
0!
0%
#750965000000
1!
1%
#750970000000
0!
0%
#750975000000
1!
1%
#750980000000
0!
0%
#750985000000
1!
1%
#750990000000
0!
0%
#750995000000
1!
1%
#751000000000
0!
0%
#751005000000
1!
1%
#751010000000
0!
0%
#751015000000
1!
1%
#751020000000
0!
0%
#751025000000
1!
1%
#751030000000
0!
0%
#751035000000
1!
1%
#751040000000
0!
0%
#751045000000
1!
1%
#751050000000
0!
0%
#751055000000
1!
1%
#751060000000
0!
0%
#751065000000
1!
1%
#751070000000
0!
0%
#751075000000
1!
1%
#751080000000
0!
0%
#751085000000
1!
1%
#751090000000
0!
0%
#751095000000
1!
1%
#751100000000
0!
0%
#751105000000
1!
1%
#751110000000
0!
0%
#751115000000
1!
1%
#751120000000
0!
0%
#751125000000
1!
1%
#751130000000
0!
0%
#751135000000
1!
1%
#751140000000
0!
0%
#751145000000
1!
1%
#751150000000
0!
0%
#751155000000
1!
1%
#751160000000
0!
0%
#751165000000
1!
1%
#751170000000
0!
0%
#751175000000
1!
1%
#751180000000
0!
0%
#751185000000
1!
1%
#751190000000
0!
0%
#751195000000
1!
1%
#751200000000
0!
0%
#751205000000
1!
1%
#751210000000
0!
0%
#751215000000
1!
1%
#751220000000
0!
0%
#751225000000
1!
1%
#751230000000
0!
0%
#751235000000
1!
1%
#751240000000
0!
0%
#751245000000
1!
1%
#751250000000
0!
0%
#751255000000
1!
1%
#751260000000
0!
0%
#751265000000
1!
1%
#751270000000
0!
0%
#751275000000
1!
1%
#751280000000
0!
0%
#751285000000
1!
1%
#751290000000
0!
0%
#751295000000
1!
1%
#751300000000
0!
0%
#751305000000
1!
1%
#751310000000
0!
0%
#751315000000
1!
1%
#751320000000
0!
0%
#751325000000
1!
1%
#751330000000
0!
0%
#751335000000
1!
1%
#751340000000
0!
0%
#751345000000
1!
1%
#751350000000
0!
0%
#751355000000
1!
1%
#751360000000
0!
0%
#751365000000
1!
1%
#751370000000
0!
0%
#751375000000
1!
1%
#751380000000
0!
0%
#751385000000
1!
1%
#751390000000
0!
0%
#751395000000
1!
1%
#751400000000
0!
0%
#751405000000
1!
1%
#751410000000
0!
0%
#751415000000
1!
1%
#751420000000
0!
0%
#751425000000
1!
1%
#751430000000
0!
0%
#751435000000
1!
1%
#751440000000
0!
0%
#751445000000
1!
1%
#751450000000
0!
0%
#751455000000
1!
1%
#751460000000
0!
0%
#751465000000
1!
1%
#751470000000
0!
0%
#751475000000
1!
1%
#751480000000
0!
0%
#751485000000
1!
1%
#751490000000
0!
0%
#751495000000
1!
1%
#751500000000
0!
0%
#751505000000
1!
1%
#751510000000
0!
0%
#751515000000
1!
1%
#751520000000
0!
0%
#751525000000
1!
1%
#751530000000
0!
0%
#751535000000
1!
1%
#751540000000
0!
0%
#751545000000
1!
1%
#751550000000
0!
0%
#751555000000
1!
1%
#751560000000
0!
0%
#751565000000
1!
1%
#751570000000
0!
0%
#751575000000
1!
1%
#751580000000
0!
0%
#751585000000
1!
1%
#751590000000
0!
0%
#751595000000
1!
1%
#751600000000
0!
0%
#751605000000
1!
1%
#751610000000
0!
0%
#751615000000
1!
1%
#751620000000
0!
0%
#751625000000
1!
1%
#751630000000
0!
0%
#751635000000
1!
1%
#751640000000
0!
0%
#751645000000
1!
1%
#751650000000
0!
0%
#751655000000
1!
1%
#751660000000
0!
0%
#751665000000
1!
1%
#751670000000
0!
0%
#751675000000
1!
1%
#751680000000
0!
0%
#751685000000
1!
1%
#751690000000
0!
0%
#751695000000
1!
1%
#751700000000
0!
0%
#751705000000
1!
1%
#751710000000
0!
0%
#751715000000
1!
1%
#751720000000
0!
0%
#751725000000
1!
1%
#751730000000
0!
0%
#751735000000
1!
1%
#751740000000
0!
0%
#751745000000
1!
1%
#751750000000
0!
0%
#751755000000
1!
1%
#751760000000
0!
0%
#751765000000
1!
1%
#751770000000
0!
0%
#751775000000
1!
1%
#751780000000
0!
0%
#751785000000
1!
1%
#751790000000
0!
0%
#751795000000
1!
1%
#751800000000
0!
0%
#751805000000
1!
1%
#751810000000
0!
0%
#751815000000
1!
1%
#751820000000
0!
0%
#751825000000
1!
1%
#751830000000
0!
0%
#751835000000
1!
1%
#751840000000
0!
0%
#751845000000
1!
1%
#751850000000
0!
0%
#751855000000
1!
1%
#751860000000
0!
0%
#751865000000
1!
1%
#751870000000
0!
0%
#751875000000
1!
1%
#751880000000
0!
0%
#751885000000
1!
1%
#751890000000
0!
0%
#751895000000
1!
1%
#751900000000
0!
0%
#751905000000
1!
1%
#751910000000
0!
0%
#751915000000
1!
1%
#751920000000
0!
0%
#751925000000
1!
1%
#751930000000
0!
0%
#751935000000
1!
1%
#751940000000
0!
0%
#751945000000
1!
1%
#751950000000
0!
0%
#751955000000
1!
1%
#751960000000
0!
0%
#751965000000
1!
1%
#751970000000
0!
0%
#751975000000
1!
1%
#751980000000
0!
0%
#751985000000
1!
1%
#751990000000
0!
0%
#751995000000
1!
1%
#752000000000
0!
0%
#752005000000
1!
1%
#752010000000
0!
0%
#752015000000
1!
1%
#752020000000
0!
0%
#752025000000
1!
1%
#752030000000
0!
0%
#752035000000
1!
1%
#752040000000
0!
0%
#752045000000
1!
1%
#752050000000
0!
0%
#752055000000
1!
1%
#752060000000
0!
0%
#752065000000
1!
1%
#752070000000
0!
0%
#752075000000
1!
1%
#752080000000
0!
0%
#752085000000
1!
1%
#752090000000
0!
0%
#752095000000
1!
1%
#752100000000
0!
0%
#752105000000
1!
1%
#752110000000
0!
0%
#752115000000
1!
1%
#752120000000
0!
0%
#752125000000
1!
1%
#752130000000
0!
0%
#752135000000
1!
1%
#752140000000
0!
0%
#752145000000
1!
1%
#752150000000
0!
0%
#752155000000
1!
1%
#752160000000
0!
0%
#752165000000
1!
1%
#752170000000
0!
0%
#752175000000
1!
1%
#752180000000
0!
0%
#752185000000
1!
1%
#752190000000
0!
0%
#752195000000
1!
1%
#752200000000
0!
0%
#752205000000
1!
1%
#752210000000
0!
0%
#752215000000
1!
1%
#752220000000
0!
0%
#752225000000
1!
1%
#752230000000
0!
0%
#752235000000
1!
1%
#752240000000
0!
0%
#752245000000
1!
1%
#752250000000
0!
0%
#752255000000
1!
1%
#752260000000
0!
0%
#752265000000
1!
1%
#752270000000
0!
0%
#752275000000
1!
1%
#752280000000
0!
0%
#752285000000
1!
1%
#752290000000
0!
0%
#752295000000
1!
1%
#752300000000
0!
0%
#752305000000
1!
1%
#752310000000
0!
0%
#752315000000
1!
1%
#752320000000
0!
0%
#752325000000
1!
1%
#752330000000
0!
0%
#752335000000
1!
1%
#752340000000
0!
0%
#752345000000
1!
1%
#752350000000
0!
0%
#752355000000
1!
1%
#752360000000
0!
0%
#752365000000
1!
1%
#752370000000
0!
0%
#752375000000
1!
1%
#752380000000
0!
0%
#752385000000
1!
1%
#752390000000
0!
0%
#752395000000
1!
1%
#752400000000
0!
0%
#752405000000
1!
1%
#752410000000
0!
0%
#752415000000
1!
1%
#752420000000
0!
0%
#752425000000
1!
1%
#752430000000
0!
0%
#752435000000
1!
1%
#752440000000
0!
0%
#752445000000
1!
1%
#752450000000
0!
0%
#752455000000
1!
1%
#752460000000
0!
0%
#752465000000
1!
1%
#752470000000
0!
0%
#752475000000
1!
1%
#752480000000
0!
0%
#752485000000
1!
1%
#752490000000
0!
0%
#752495000000
1!
1%
#752500000000
0!
0%
#752505000000
1!
1%
#752510000000
0!
0%
#752515000000
1!
1%
#752520000000
0!
0%
#752525000000
1!
1%
#752530000000
0!
0%
#752535000000
1!
1%
#752540000000
0!
0%
#752545000000
1!
1%
#752550000000
0!
0%
#752555000000
1!
1%
#752560000000
0!
0%
#752565000000
1!
1%
#752570000000
0!
0%
#752575000000
1!
1%
#752580000000
0!
0%
#752585000000
1!
1%
#752590000000
0!
0%
#752595000000
1!
1%
#752600000000
0!
0%
#752605000000
1!
1%
#752610000000
0!
0%
#752615000000
1!
1%
#752620000000
0!
0%
#752625000000
1!
1%
#752630000000
0!
0%
#752635000000
1!
1%
#752640000000
0!
0%
#752645000000
1!
1%
#752650000000
0!
0%
#752655000000
1!
1%
#752660000000
0!
0%
#752665000000
1!
1%
#752670000000
0!
0%
#752675000000
1!
1%
#752680000000
0!
0%
#752685000000
1!
1%
#752690000000
0!
0%
#752695000000
1!
1%
#752700000000
0!
0%
#752705000000
1!
1%
#752710000000
0!
0%
#752715000000
1!
1%
#752720000000
0!
0%
#752725000000
1!
1%
#752730000000
0!
0%
#752735000000
1!
1%
#752740000000
0!
0%
#752745000000
1!
1%
#752750000000
0!
0%
#752755000000
1!
1%
#752760000000
0!
0%
#752765000000
1!
1%
#752770000000
0!
0%
#752775000000
1!
1%
#752780000000
0!
0%
#752785000000
1!
1%
#752790000000
0!
0%
#752795000000
1!
1%
#752800000000
0!
0%
#752805000000
1!
1%
#752810000000
0!
0%
#752815000000
1!
1%
#752820000000
0!
0%
#752825000000
1!
1%
#752830000000
0!
0%
#752835000000
1!
1%
#752840000000
0!
0%
#752845000000
1!
1%
#752850000000
0!
0%
#752855000000
1!
1%
#752860000000
0!
0%
#752865000000
1!
1%
#752870000000
0!
0%
#752875000000
1!
1%
#752880000000
0!
0%
#752885000000
1!
1%
#752890000000
0!
0%
#752895000000
1!
1%
#752900000000
0!
0%
#752905000000
1!
1%
#752910000000
0!
0%
#752915000000
1!
1%
#752920000000
0!
0%
#752925000000
1!
1%
#752930000000
0!
0%
#752935000000
1!
1%
#752940000000
0!
0%
#752945000000
1!
1%
#752950000000
0!
0%
#752955000000
1!
1%
#752960000000
0!
0%
#752965000000
1!
1%
#752970000000
0!
0%
#752975000000
1!
1%
#752980000000
0!
0%
#752985000000
1!
1%
#752990000000
0!
0%
#752995000000
1!
1%
#753000000000
0!
0%
#753005000000
1!
1%
#753010000000
0!
0%
#753015000000
1!
1%
#753020000000
0!
0%
#753025000000
1!
1%
#753030000000
0!
0%
#753035000000
1!
1%
#753040000000
0!
0%
#753045000000
1!
1%
#753050000000
0!
0%
#753055000000
1!
1%
#753060000000
0!
0%
#753065000000
1!
1%
#753070000000
0!
0%
#753075000000
1!
1%
#753080000000
0!
0%
#753085000000
1!
1%
#753090000000
0!
0%
#753095000000
1!
1%
#753100000000
0!
0%
#753105000000
1!
1%
#753110000000
0!
0%
#753115000000
1!
1%
#753120000000
0!
0%
#753125000000
1!
1%
#753130000000
0!
0%
#753135000000
1!
1%
#753140000000
0!
0%
#753145000000
1!
1%
#753150000000
0!
0%
#753155000000
1!
1%
#753160000000
0!
0%
#753165000000
1!
1%
#753170000000
0!
0%
#753175000000
1!
1%
#753180000000
0!
0%
#753185000000
1!
1%
#753190000000
0!
0%
#753195000000
1!
1%
#753200000000
0!
0%
#753205000000
1!
1%
#753210000000
0!
0%
#753215000000
1!
1%
#753220000000
0!
0%
#753225000000
1!
1%
#753230000000
0!
0%
#753235000000
1!
1%
#753240000000
0!
0%
#753245000000
1!
1%
#753250000000
0!
0%
#753255000000
1!
1%
#753260000000
0!
0%
#753265000000
1!
1%
#753270000000
0!
0%
#753275000000
1!
1%
#753280000000
0!
0%
#753285000000
1!
1%
#753290000000
0!
0%
#753295000000
1!
1%
#753300000000
0!
0%
#753305000000
1!
1%
#753310000000
0!
0%
#753315000000
1!
1%
#753320000000
0!
0%
#753325000000
1!
1%
#753330000000
0!
0%
#753335000000
1!
1%
#753340000000
0!
0%
#753345000000
1!
1%
#753350000000
0!
0%
#753355000000
1!
1%
#753360000000
0!
0%
#753365000000
1!
1%
#753370000000
0!
0%
#753375000000
1!
1%
#753380000000
0!
0%
#753385000000
1!
1%
#753390000000
0!
0%
#753395000000
1!
1%
#753400000000
0!
0%
#753405000000
1!
1%
#753410000000
0!
0%
#753415000000
1!
1%
#753420000000
0!
0%
#753425000000
1!
1%
#753430000000
0!
0%
#753435000000
1!
1%
#753440000000
0!
0%
#753445000000
1!
1%
#753450000000
0!
0%
#753455000000
1!
1%
#753460000000
0!
0%
#753465000000
1!
1%
#753470000000
0!
0%
#753475000000
1!
1%
#753480000000
0!
0%
#753485000000
1!
1%
#753490000000
0!
0%
#753495000000
1!
1%
#753500000000
0!
0%
#753505000000
1!
1%
#753510000000
0!
0%
#753515000000
1!
1%
#753520000000
0!
0%
#753525000000
1!
1%
#753530000000
0!
0%
#753535000000
1!
1%
#753540000000
0!
0%
#753545000000
1!
1%
#753550000000
0!
0%
#753555000000
1!
1%
#753560000000
0!
0%
#753565000000
1!
1%
#753570000000
0!
0%
#753575000000
1!
1%
#753580000000
0!
0%
#753585000000
1!
1%
#753590000000
0!
0%
#753595000000
1!
1%
#753600000000
0!
0%
#753605000000
1!
1%
#753610000000
0!
0%
#753615000000
1!
1%
#753620000000
0!
0%
#753625000000
1!
1%
#753630000000
0!
0%
#753635000000
1!
1%
#753640000000
0!
0%
#753645000000
1!
1%
#753650000000
0!
0%
#753655000000
1!
1%
#753660000000
0!
0%
#753665000000
1!
1%
#753670000000
0!
0%
#753675000000
1!
1%
#753680000000
0!
0%
#753685000000
1!
1%
#753690000000
0!
0%
#753695000000
1!
1%
#753700000000
0!
0%
#753705000000
1!
1%
#753710000000
0!
0%
#753715000000
1!
1%
#753720000000
0!
0%
#753725000000
1!
1%
#753730000000
0!
0%
#753735000000
1!
1%
#753740000000
0!
0%
#753745000000
1!
1%
#753750000000
0!
0%
#753755000000
1!
1%
#753760000000
0!
0%
#753765000000
1!
1%
#753770000000
0!
0%
#753775000000
1!
1%
#753780000000
0!
0%
#753785000000
1!
1%
#753790000000
0!
0%
#753795000000
1!
1%
#753800000000
0!
0%
#753805000000
1!
1%
#753810000000
0!
0%
#753815000000
1!
1%
#753820000000
0!
0%
#753825000000
1!
1%
#753830000000
0!
0%
#753835000000
1!
1%
#753840000000
0!
0%
#753845000000
1!
1%
#753850000000
0!
0%
#753855000000
1!
1%
#753860000000
0!
0%
#753865000000
1!
1%
#753870000000
0!
0%
#753875000000
1!
1%
#753880000000
0!
0%
#753885000000
1!
1%
#753890000000
0!
0%
#753895000000
1!
1%
#753900000000
0!
0%
#753905000000
1!
1%
#753910000000
0!
0%
#753915000000
1!
1%
#753920000000
0!
0%
#753925000000
1!
1%
#753930000000
0!
0%
#753935000000
1!
1%
#753940000000
0!
0%
#753945000000
1!
1%
#753950000000
0!
0%
#753955000000
1!
1%
#753960000000
0!
0%
#753965000000
1!
1%
#753970000000
0!
0%
#753975000000
1!
1%
#753980000000
0!
0%
#753985000000
1!
1%
#753990000000
0!
0%
#753995000000
1!
1%
#754000000000
0!
0%
#754005000000
1!
1%
#754010000000
0!
0%
#754015000000
1!
1%
#754020000000
0!
0%
#754025000000
1!
1%
#754030000000
0!
0%
#754035000000
1!
1%
#754040000000
0!
0%
#754045000000
1!
1%
#754050000000
0!
0%
#754055000000
1!
1%
#754060000000
0!
0%
#754065000000
1!
1%
#754070000000
0!
0%
#754075000000
1!
1%
#754080000000
0!
0%
#754085000000
1!
1%
#754090000000
0!
0%
#754095000000
1!
1%
#754100000000
0!
0%
#754105000000
1!
1%
#754110000000
0!
0%
#754115000000
1!
1%
#754120000000
0!
0%
#754125000000
1!
1%
#754130000000
0!
0%
#754135000000
1!
1%
#754140000000
0!
0%
#754145000000
1!
1%
#754150000000
0!
0%
#754155000000
1!
1%
#754160000000
0!
0%
#754165000000
1!
1%
#754170000000
0!
0%
#754175000000
1!
1%
#754180000000
0!
0%
#754185000000
1!
1%
#754190000000
0!
0%
#754195000000
1!
1%
#754200000000
0!
0%
#754205000000
1!
1%
#754210000000
0!
0%
#754215000000
1!
1%
#754220000000
0!
0%
#754225000000
1!
1%
#754230000000
0!
0%
#754235000000
1!
1%
#754240000000
0!
0%
#754245000000
1!
1%
#754250000000
0!
0%
#754255000000
1!
1%
#754260000000
0!
0%
#754265000000
1!
1%
#754270000000
0!
0%
#754275000000
1!
1%
#754280000000
0!
0%
#754285000000
1!
1%
#754290000000
0!
0%
#754295000000
1!
1%
#754300000000
0!
0%
#754305000000
1!
1%
#754310000000
0!
0%
#754315000000
1!
1%
#754320000000
0!
0%
#754325000000
1!
1%
#754330000000
0!
0%
#754335000000
1!
1%
#754340000000
0!
0%
#754345000000
1!
1%
#754350000000
0!
0%
#754355000000
1!
1%
#754360000000
0!
0%
#754365000000
1!
1%
#754370000000
0!
0%
#754375000000
1!
1%
#754380000000
0!
0%
#754385000000
1!
1%
#754390000000
0!
0%
#754395000000
1!
1%
#754400000000
0!
0%
#754405000000
1!
1%
#754410000000
0!
0%
#754415000000
1!
1%
#754420000000
0!
0%
#754425000000
1!
1%
#754430000000
0!
0%
#754435000000
1!
1%
#754440000000
0!
0%
#754445000000
1!
1%
#754450000000
0!
0%
#754455000000
1!
1%
#754460000000
0!
0%
#754465000000
1!
1%
#754470000000
0!
0%
#754475000000
1!
1%
#754480000000
0!
0%
#754485000000
1!
1%
#754490000000
0!
0%
#754495000000
1!
1%
#754500000000
0!
0%
#754505000000
1!
1%
#754510000000
0!
0%
#754515000000
1!
1%
#754520000000
0!
0%
#754525000000
1!
1%
#754530000000
0!
0%
#754535000000
1!
1%
#754540000000
0!
0%
#754545000000
1!
1%
#754550000000
0!
0%
#754555000000
1!
1%
#754560000000
0!
0%
#754565000000
1!
1%
#754570000000
0!
0%
#754575000000
1!
1%
#754580000000
0!
0%
#754585000000
1!
1%
#754590000000
0!
0%
#754595000000
1!
1%
#754600000000
0!
0%
#754605000000
1!
1%
#754610000000
0!
0%
#754615000000
1!
1%
#754620000000
0!
0%
#754625000000
1!
1%
#754630000000
0!
0%
#754635000000
1!
1%
#754640000000
0!
0%
#754645000000
1!
1%
#754650000000
0!
0%
#754655000000
1!
1%
#754660000000
0!
0%
#754665000000
1!
1%
#754670000000
0!
0%
#754675000000
1!
1%
#754680000000
0!
0%
#754685000000
1!
1%
#754690000000
0!
0%
#754695000000
1!
1%
#754700000000
0!
0%
#754705000000
1!
1%
#754710000000
0!
0%
#754715000000
1!
1%
#754720000000
0!
0%
#754725000000
1!
1%
#754730000000
0!
0%
#754735000000
1!
1%
#754740000000
0!
0%
#754745000000
1!
1%
#754750000000
0!
0%
#754755000000
1!
1%
#754760000000
0!
0%
#754765000000
1!
1%
#754770000000
0!
0%
#754775000000
1!
1%
#754780000000
0!
0%
#754785000000
1!
1%
#754790000000
0!
0%
#754795000000
1!
1%
#754800000000
0!
0%
#754805000000
1!
1%
#754810000000
0!
0%
#754815000000
1!
1%
#754820000000
0!
0%
#754825000000
1!
1%
#754830000000
0!
0%
#754835000000
1!
1%
#754840000000
0!
0%
#754845000000
1!
1%
#754850000000
0!
0%
#754855000000
1!
1%
#754860000000
0!
0%
#754865000000
1!
1%
#754870000000
0!
0%
#754875000000
1!
1%
#754880000000
0!
0%
#754885000000
1!
1%
#754890000000
0!
0%
#754895000000
1!
1%
#754900000000
0!
0%
#754905000000
1!
1%
#754910000000
0!
0%
#754915000000
1!
1%
#754920000000
0!
0%
#754925000000
1!
1%
#754930000000
0!
0%
#754935000000
1!
1%
#754940000000
0!
0%
#754945000000
1!
1%
#754950000000
0!
0%
#754955000000
1!
1%
#754960000000
0!
0%
#754965000000
1!
1%
#754970000000
0!
0%
#754975000000
1!
1%
#754980000000
0!
0%
#754985000000
1!
1%
#754990000000
0!
0%
#754995000000
1!
1%
#755000000000
0!
0%
#755005000000
1!
1%
#755010000000
0!
0%
#755015000000
1!
1%
#755020000000
0!
0%
#755025000000
1!
1%
#755030000000
0!
0%
#755035000000
1!
1%
#755040000000
0!
0%
#755045000000
1!
1%
#755050000000
0!
0%
#755055000000
1!
1%
#755060000000
0!
0%
#755065000000
1!
1%
#755070000000
0!
0%
#755075000000
1!
1%
#755080000000
0!
0%
#755085000000
1!
1%
#755090000000
0!
0%
#755095000000
1!
1%
#755100000000
0!
0%
#755105000000
1!
1%
#755110000000
0!
0%
#755115000000
1!
1%
#755120000000
0!
0%
#755125000000
1!
1%
#755130000000
0!
0%
#755135000000
1!
1%
#755140000000
0!
0%
#755145000000
1!
1%
#755150000000
0!
0%
#755155000000
1!
1%
#755160000000
0!
0%
#755165000000
1!
1%
#755170000000
0!
0%
#755175000000
1!
1%
#755180000000
0!
0%
#755185000000
1!
1%
#755190000000
0!
0%
#755195000000
1!
1%
#755200000000
0!
0%
#755205000000
1!
1%
#755210000000
0!
0%
#755215000000
1!
1%
#755220000000
0!
0%
#755225000000
1!
1%
#755230000000
0!
0%
#755235000000
1!
1%
#755240000000
0!
0%
#755245000000
1!
1%
#755250000000
0!
0%
#755255000000
1!
1%
#755260000000
0!
0%
#755265000000
1!
1%
#755270000000
0!
0%
#755275000000
1!
1%
#755280000000
0!
0%
#755285000000
1!
1%
#755290000000
0!
0%
#755295000000
1!
1%
#755300000000
0!
0%
#755305000000
1!
1%
#755310000000
0!
0%
#755315000000
1!
1%
#755320000000
0!
0%
#755325000000
1!
1%
#755330000000
0!
0%
#755335000000
1!
1%
#755340000000
0!
0%
#755345000000
1!
1%
#755350000000
0!
0%
#755355000000
1!
1%
#755360000000
0!
0%
#755365000000
1!
1%
#755370000000
0!
0%
#755375000000
1!
1%
#755380000000
0!
0%
#755385000000
1!
1%
#755390000000
0!
0%
#755395000000
1!
1%
#755400000000
0!
0%
#755405000000
1!
1%
#755410000000
0!
0%
#755415000000
1!
1%
#755420000000
0!
0%
#755425000000
1!
1%
#755430000000
0!
0%
#755435000000
1!
1%
#755440000000
0!
0%
#755445000000
1!
1%
#755450000000
0!
0%
#755455000000
1!
1%
#755460000000
0!
0%
#755465000000
1!
1%
#755470000000
0!
0%
#755475000000
1!
1%
#755480000000
0!
0%
#755485000000
1!
1%
#755490000000
0!
0%
#755495000000
1!
1%
#755500000000
0!
0%
#755505000000
1!
1%
#755510000000
0!
0%
#755515000000
1!
1%
#755520000000
0!
0%
#755525000000
1!
1%
#755530000000
0!
0%
#755535000000
1!
1%
#755540000000
0!
0%
#755545000000
1!
1%
#755550000000
0!
0%
#755555000000
1!
1%
#755560000000
0!
0%
#755565000000
1!
1%
#755570000000
0!
0%
#755575000000
1!
1%
#755580000000
0!
0%
#755585000000
1!
1%
#755590000000
0!
0%
#755595000000
1!
1%
#755600000000
0!
0%
#755605000000
1!
1%
#755610000000
0!
0%
#755615000000
1!
1%
#755620000000
0!
0%
#755625000000
1!
1%
#755630000000
0!
0%
#755635000000
1!
1%
#755640000000
0!
0%
#755645000000
1!
1%
#755650000000
0!
0%
#755655000000
1!
1%
#755660000000
0!
0%
#755665000000
1!
1%
#755670000000
0!
0%
#755675000000
1!
1%
#755680000000
0!
0%
#755685000000
1!
1%
#755690000000
0!
0%
#755695000000
1!
1%
#755700000000
0!
0%
#755705000000
1!
1%
#755710000000
0!
0%
#755715000000
1!
1%
#755720000000
0!
0%
#755725000000
1!
1%
#755730000000
0!
0%
#755735000000
1!
1%
#755740000000
0!
0%
#755745000000
1!
1%
#755750000000
0!
0%
#755755000000
1!
1%
#755760000000
0!
0%
#755765000000
1!
1%
#755770000000
0!
0%
#755775000000
1!
1%
#755780000000
0!
0%
#755785000000
1!
1%
#755790000000
0!
0%
#755795000000
1!
1%
#755800000000
0!
0%
#755805000000
1!
1%
#755810000000
0!
0%
#755815000000
1!
1%
#755820000000
0!
0%
#755825000000
1!
1%
#755830000000
0!
0%
#755835000000
1!
1%
#755840000000
0!
0%
#755845000000
1!
1%
#755850000000
0!
0%
#755855000000
1!
1%
#755860000000
0!
0%
#755865000000
1!
1%
#755870000000
0!
0%
#755875000000
1!
1%
#755880000000
0!
0%
#755885000000
1!
1%
#755890000000
0!
0%
#755895000000
1!
1%
#755900000000
0!
0%
#755905000000
1!
1%
#755910000000
0!
0%
#755915000000
1!
1%
#755920000000
0!
0%
#755925000000
1!
1%
#755930000000
0!
0%
#755935000000
1!
1%
#755940000000
0!
0%
#755945000000
1!
1%
#755950000000
0!
0%
#755955000000
1!
1%
#755960000000
0!
0%
#755965000000
1!
1%
#755970000000
0!
0%
#755975000000
1!
1%
#755980000000
0!
0%
#755985000000
1!
1%
#755990000000
0!
0%
#755995000000
1!
1%
#756000000000
0!
0%
#756005000000
1!
1%
#756010000000
0!
0%
#756015000000
1!
1%
#756020000000
0!
0%
#756025000000
1!
1%
#756030000000
0!
0%
#756035000000
1!
1%
#756040000000
0!
0%
#756045000000
1!
1%
#756050000000
0!
0%
#756055000000
1!
1%
#756060000000
0!
0%
#756065000000
1!
1%
#756070000000
0!
0%
#756075000000
1!
1%
#756080000000
0!
0%
#756085000000
1!
1%
#756090000000
0!
0%
#756095000000
1!
1%
#756100000000
0!
0%
#756105000000
1!
1%
#756110000000
0!
0%
#756115000000
1!
1%
#756120000000
0!
0%
#756125000000
1!
1%
#756130000000
0!
0%
#756135000000
1!
1%
#756140000000
0!
0%
#756145000000
1!
1%
#756150000000
0!
0%
#756155000000
1!
1%
#756160000000
0!
0%
#756165000000
1!
1%
#756170000000
0!
0%
#756175000000
1!
1%
#756180000000
0!
0%
#756185000000
1!
1%
#756190000000
0!
0%
#756195000000
1!
1%
#756200000000
0!
0%
#756205000000
1!
1%
#756210000000
0!
0%
#756215000000
1!
1%
#756220000000
0!
0%
#756225000000
1!
1%
#756230000000
0!
0%
#756235000000
1!
1%
#756240000000
0!
0%
#756245000000
1!
1%
#756250000000
0!
0%
#756255000000
1!
1%
#756260000000
0!
0%
#756265000000
1!
1%
#756270000000
0!
0%
#756275000000
1!
1%
#756280000000
0!
0%
#756285000000
1!
1%
#756290000000
0!
0%
#756295000000
1!
1%
#756300000000
0!
0%
#756305000000
1!
1%
#756310000000
0!
0%
#756315000000
1!
1%
#756320000000
0!
0%
#756325000000
1!
1%
#756330000000
0!
0%
#756335000000
1!
1%
#756340000000
0!
0%
#756345000000
1!
1%
#756350000000
0!
0%
#756355000000
1!
1%
#756360000000
0!
0%
#756365000000
1!
1%
#756370000000
0!
0%
#756375000000
1!
1%
#756380000000
0!
0%
#756385000000
1!
1%
#756390000000
0!
0%
#756395000000
1!
1%
#756400000000
0!
0%
#756405000000
1!
1%
#756410000000
0!
0%
#756415000000
1!
1%
#756420000000
0!
0%
#756425000000
1!
1%
#756430000000
0!
0%
#756435000000
1!
1%
#756440000000
0!
0%
#756445000000
1!
1%
#756450000000
0!
0%
#756455000000
1!
1%
#756460000000
0!
0%
#756465000000
1!
1%
#756470000000
0!
0%
#756475000000
1!
1%
#756480000000
0!
0%
#756485000000
1!
1%
#756490000000
0!
0%
#756495000000
1!
1%
#756500000000
0!
0%
#756505000000
1!
1%
#756510000000
0!
0%
#756515000000
1!
1%
#756520000000
0!
0%
#756525000000
1!
1%
#756530000000
0!
0%
#756535000000
1!
1%
#756540000000
0!
0%
#756545000000
1!
1%
#756550000000
0!
0%
#756555000000
1!
1%
#756560000000
0!
0%
#756565000000
1!
1%
#756570000000
0!
0%
#756575000000
1!
1%
#756580000000
0!
0%
#756585000000
1!
1%
#756590000000
0!
0%
#756595000000
1!
1%
#756600000000
0!
0%
#756605000000
1!
1%
#756610000000
0!
0%
#756615000000
1!
1%
#756620000000
0!
0%
#756625000000
1!
1%
#756630000000
0!
0%
#756635000000
1!
1%
#756640000000
0!
0%
#756645000000
1!
1%
#756650000000
0!
0%
#756655000000
1!
1%
#756660000000
0!
0%
#756665000000
1!
1%
#756670000000
0!
0%
#756675000000
1!
1%
#756680000000
0!
0%
#756685000000
1!
1%
#756690000000
0!
0%
#756695000000
1!
1%
#756700000000
0!
0%
#756705000000
1!
1%
#756710000000
0!
0%
#756715000000
1!
1%
#756720000000
0!
0%
#756725000000
1!
1%
#756730000000
0!
0%
#756735000000
1!
1%
#756740000000
0!
0%
#756745000000
1!
1%
#756750000000
0!
0%
#756755000000
1!
1%
#756760000000
0!
0%
#756765000000
1!
1%
#756770000000
0!
0%
#756775000000
1!
1%
#756780000000
0!
0%
#756785000000
1!
1%
#756790000000
0!
0%
#756795000000
1!
1%
#756800000000
0!
0%
#756805000000
1!
1%
#756810000000
0!
0%
#756815000000
1!
1%
#756820000000
0!
0%
#756825000000
1!
1%
#756830000000
0!
0%
#756835000000
1!
1%
#756840000000
0!
0%
#756845000000
1!
1%
#756850000000
0!
0%
#756855000000
1!
1%
#756860000000
0!
0%
#756865000000
1!
1%
#756870000000
0!
0%
#756875000000
1!
1%
#756880000000
0!
0%
#756885000000
1!
1%
#756890000000
0!
0%
#756895000000
1!
1%
#756900000000
0!
0%
#756905000000
1!
1%
#756910000000
0!
0%
#756915000000
1!
1%
#756920000000
0!
0%
#756925000000
1!
1%
#756930000000
0!
0%
#756935000000
1!
1%
#756940000000
0!
0%
#756945000000
1!
1%
#756950000000
0!
0%
#756955000000
1!
1%
#756960000000
0!
0%
#756965000000
1!
1%
#756970000000
0!
0%
#756975000000
1!
1%
#756980000000
0!
0%
#756985000000
1!
1%
#756990000000
0!
0%
#756995000000
1!
1%
#757000000000
0!
0%
#757005000000
1!
1%
#757010000000
0!
0%
#757015000000
1!
1%
#757020000000
0!
0%
#757025000000
1!
1%
#757030000000
0!
0%
#757035000000
1!
1%
#757040000000
0!
0%
#757045000000
1!
1%
#757050000000
0!
0%
#757055000000
1!
1%
#757060000000
0!
0%
#757065000000
1!
1%
#757070000000
0!
0%
#757075000000
1!
1%
#757080000000
0!
0%
#757085000000
1!
1%
#757090000000
0!
0%
#757095000000
1!
1%
#757100000000
0!
0%
#757105000000
1!
1%
#757110000000
0!
0%
#757115000000
1!
1%
#757120000000
0!
0%
#757125000000
1!
1%
#757130000000
0!
0%
#757135000000
1!
1%
#757140000000
0!
0%
#757145000000
1!
1%
#757150000000
0!
0%
#757155000000
1!
1%
#757160000000
0!
0%
#757165000000
1!
1%
#757170000000
0!
0%
#757175000000
1!
1%
#757180000000
0!
0%
#757185000000
1!
1%
#757190000000
0!
0%
#757195000000
1!
1%
#757200000000
0!
0%
#757205000000
1!
1%
#757210000000
0!
0%
#757215000000
1!
1%
#757220000000
0!
0%
#757225000000
1!
1%
#757230000000
0!
0%
#757235000000
1!
1%
#757240000000
0!
0%
#757245000000
1!
1%
#757250000000
0!
0%
#757255000000
1!
1%
#757260000000
0!
0%
#757265000000
1!
1%
#757270000000
0!
0%
#757275000000
1!
1%
#757280000000
0!
0%
#757285000000
1!
1%
#757290000000
0!
0%
#757295000000
1!
1%
#757300000000
0!
0%
#757305000000
1!
1%
#757310000000
0!
0%
#757315000000
1!
1%
#757320000000
0!
0%
#757325000000
1!
1%
#757330000000
0!
0%
#757335000000
1!
1%
#757340000000
0!
0%
#757345000000
1!
1%
#757350000000
0!
0%
#757355000000
1!
1%
#757360000000
0!
0%
#757365000000
1!
1%
#757370000000
0!
0%
#757375000000
1!
1%
#757380000000
0!
0%
#757385000000
1!
1%
#757390000000
0!
0%
#757395000000
1!
1%
#757400000000
0!
0%
#757405000000
1!
1%
#757410000000
0!
0%
#757415000000
1!
1%
#757420000000
0!
0%
#757425000000
1!
1%
#757430000000
0!
0%
#757435000000
1!
1%
#757440000000
0!
0%
#757445000000
1!
1%
#757450000000
0!
0%
#757455000000
1!
1%
#757460000000
0!
0%
#757465000000
1!
1%
#757470000000
0!
0%
#757475000000
1!
1%
#757480000000
0!
0%
#757485000000
1!
1%
#757490000000
0!
0%
#757495000000
1!
1%
#757500000000
0!
0%
#757505000000
1!
1%
#757510000000
0!
0%
#757515000000
1!
1%
#757520000000
0!
0%
#757525000000
1!
1%
#757530000000
0!
0%
#757535000000
1!
1%
#757540000000
0!
0%
#757545000000
1!
1%
#757550000000
0!
0%
#757555000000
1!
1%
#757560000000
0!
0%
#757565000000
1!
1%
#757570000000
0!
0%
#757575000000
1!
1%
#757580000000
0!
0%
#757585000000
1!
1%
#757590000000
0!
0%
#757595000000
1!
1%
#757600000000
0!
0%
#757605000000
1!
1%
#757610000000
0!
0%
#757615000000
1!
1%
#757620000000
0!
0%
#757625000000
1!
1%
#757630000000
0!
0%
#757635000000
1!
1%
#757640000000
0!
0%
#757645000000
1!
1%
#757650000000
0!
0%
#757655000000
1!
1%
#757660000000
0!
0%
#757665000000
1!
1%
#757670000000
0!
0%
#757675000000
1!
1%
#757680000000
0!
0%
#757685000000
1!
1%
#757690000000
0!
0%
#757695000000
1!
1%
#757700000000
0!
0%
#757705000000
1!
1%
#757710000000
0!
0%
#757715000000
1!
1%
#757720000000
0!
0%
#757725000000
1!
1%
#757730000000
0!
0%
#757735000000
1!
1%
#757740000000
0!
0%
#757745000000
1!
1%
#757750000000
0!
0%
#757755000000
1!
1%
#757760000000
0!
0%
#757765000000
1!
1%
#757770000000
0!
0%
#757775000000
1!
1%
#757780000000
0!
0%
#757785000000
1!
1%
#757790000000
0!
0%
#757795000000
1!
1%
#757800000000
0!
0%
#757805000000
1!
1%
#757810000000
0!
0%
#757815000000
1!
1%
#757820000000
0!
0%
#757825000000
1!
1%
#757830000000
0!
0%
#757835000000
1!
1%
#757840000000
0!
0%
#757845000000
1!
1%
#757850000000
0!
0%
#757855000000
1!
1%
#757860000000
0!
0%
#757865000000
1!
1%
#757870000000
0!
0%
#757875000000
1!
1%
#757880000000
0!
0%
#757885000000
1!
1%
#757890000000
0!
0%
#757895000000
1!
1%
#757900000000
0!
0%
#757905000000
1!
1%
#757910000000
0!
0%
#757915000000
1!
1%
#757920000000
0!
0%
#757925000000
1!
1%
#757930000000
0!
0%
#757935000000
1!
1%
#757940000000
0!
0%
#757945000000
1!
1%
#757950000000
0!
0%
#757955000000
1!
1%
#757960000000
0!
0%
#757965000000
1!
1%
#757970000000
0!
0%
#757975000000
1!
1%
#757980000000
0!
0%
#757985000000
1!
1%
#757990000000
0!
0%
#757995000000
1!
1%
#758000000000
0!
0%
#758005000000
1!
1%
#758010000000
0!
0%
#758015000000
1!
1%
#758020000000
0!
0%
#758025000000
1!
1%
#758030000000
0!
0%
#758035000000
1!
1%
#758040000000
0!
0%
#758045000000
1!
1%
#758050000000
0!
0%
#758055000000
1!
1%
#758060000000
0!
0%
#758065000000
1!
1%
#758070000000
0!
0%
#758075000000
1!
1%
#758080000000
0!
0%
#758085000000
1!
1%
#758090000000
0!
0%
#758095000000
1!
1%
#758100000000
0!
0%
#758105000000
1!
1%
#758110000000
0!
0%
#758115000000
1!
1%
#758120000000
0!
0%
#758125000000
1!
1%
#758130000000
0!
0%
#758135000000
1!
1%
#758140000000
0!
0%
#758145000000
1!
1%
#758150000000
0!
0%
#758155000000
1!
1%
#758160000000
0!
0%
#758165000000
1!
1%
#758170000000
0!
0%
#758175000000
1!
1%
#758180000000
0!
0%
#758185000000
1!
1%
#758190000000
0!
0%
#758195000000
1!
1%
#758200000000
0!
0%
#758205000000
1!
1%
#758210000000
0!
0%
#758215000000
1!
1%
#758220000000
0!
0%
#758225000000
1!
1%
#758230000000
0!
0%
#758235000000
1!
1%
#758240000000
0!
0%
#758245000000
1!
1%
#758250000000
0!
0%
#758255000000
1!
1%
#758260000000
0!
0%
#758265000000
1!
1%
#758270000000
0!
0%
#758275000000
1!
1%
#758280000000
0!
0%
#758285000000
1!
1%
#758290000000
0!
0%
#758295000000
1!
1%
#758300000000
0!
0%
#758305000000
1!
1%
#758310000000
0!
0%
#758315000000
1!
1%
#758320000000
0!
0%
#758325000000
1!
1%
#758330000000
0!
0%
#758335000000
1!
1%
#758340000000
0!
0%
#758345000000
1!
1%
#758350000000
0!
0%
#758355000000
1!
1%
#758360000000
0!
0%
#758365000000
1!
1%
#758370000000
0!
0%
#758375000000
1!
1%
#758380000000
0!
0%
#758385000000
1!
1%
#758390000000
0!
0%
#758395000000
1!
1%
#758400000000
0!
0%
#758405000000
1!
1%
#758410000000
0!
0%
#758415000000
1!
1%
#758420000000
0!
0%
#758425000000
1!
1%
#758430000000
0!
0%
#758435000000
1!
1%
#758440000000
0!
0%
#758445000000
1!
1%
#758450000000
0!
0%
#758455000000
1!
1%
#758460000000
0!
0%
#758465000000
1!
1%
#758470000000
0!
0%
#758475000000
1!
1%
#758480000000
0!
0%
#758485000000
1!
1%
#758490000000
0!
0%
#758495000000
1!
1%
#758500000000
0!
0%
#758505000000
1!
1%
#758510000000
0!
0%
#758515000000
1!
1%
#758520000000
0!
0%
#758525000000
1!
1%
#758530000000
0!
0%
#758535000000
1!
1%
#758540000000
0!
0%
#758545000000
1!
1%
#758550000000
0!
0%
#758555000000
1!
1%
#758560000000
0!
0%
#758565000000
1!
1%
#758570000000
0!
0%
#758575000000
1!
1%
#758580000000
0!
0%
#758585000000
1!
1%
#758590000000
0!
0%
#758595000000
1!
1%
#758600000000
0!
0%
#758605000000
1!
1%
#758610000000
0!
0%
#758615000000
1!
1%
#758620000000
0!
0%
#758625000000
1!
1%
#758630000000
0!
0%
#758635000000
1!
1%
#758640000000
0!
0%
#758645000000
1!
1%
#758650000000
0!
0%
#758655000000
1!
1%
#758660000000
0!
0%
#758665000000
1!
1%
#758670000000
0!
0%
#758675000000
1!
1%
#758680000000
0!
0%
#758685000000
1!
1%
#758690000000
0!
0%
#758695000000
1!
1%
#758700000000
0!
0%
#758705000000
1!
1%
#758710000000
0!
0%
#758715000000
1!
1%
#758720000000
0!
0%
#758725000000
1!
1%
#758730000000
0!
0%
#758735000000
1!
1%
#758740000000
0!
0%
#758745000000
1!
1%
#758750000000
0!
0%
#758755000000
1!
1%
#758760000000
0!
0%
#758765000000
1!
1%
#758770000000
0!
0%
#758775000000
1!
1%
#758780000000
0!
0%
#758785000000
1!
1%
#758790000000
0!
0%
#758795000000
1!
1%
#758800000000
0!
0%
#758805000000
1!
1%
#758810000000
0!
0%
#758815000000
1!
1%
#758820000000
0!
0%
#758825000000
1!
1%
#758830000000
0!
0%
#758835000000
1!
1%
#758840000000
0!
0%
#758845000000
1!
1%
#758850000000
0!
0%
#758855000000
1!
1%
#758860000000
0!
0%
#758865000000
1!
1%
#758870000000
0!
0%
#758875000000
1!
1%
#758880000000
0!
0%
#758885000000
1!
1%
#758890000000
0!
0%
#758895000000
1!
1%
#758900000000
0!
0%
#758905000000
1!
1%
#758910000000
0!
0%
#758915000000
1!
1%
#758920000000
0!
0%
#758925000000
1!
1%
#758930000000
0!
0%
#758935000000
1!
1%
#758940000000
0!
0%
#758945000000
1!
1%
#758950000000
0!
0%
#758955000000
1!
1%
#758960000000
0!
0%
#758965000000
1!
1%
#758970000000
0!
0%
#758975000000
1!
1%
#758980000000
0!
0%
#758985000000
1!
1%
#758990000000
0!
0%
#758995000000
1!
1%
#759000000000
0!
0%
#759005000000
1!
1%
#759010000000
0!
0%
#759015000000
1!
1%
#759020000000
0!
0%
#759025000000
1!
1%
#759030000000
0!
0%
#759035000000
1!
1%
#759040000000
0!
0%
#759045000000
1!
1%
#759050000000
0!
0%
#759055000000
1!
1%
#759060000000
0!
0%
#759065000000
1!
1%
#759070000000
0!
0%
#759075000000
1!
1%
#759080000000
0!
0%
#759085000000
1!
1%
#759090000000
0!
0%
#759095000000
1!
1%
#759100000000
0!
0%
#759105000000
1!
1%
#759110000000
0!
0%
#759115000000
1!
1%
#759120000000
0!
0%
#759125000000
1!
1%
#759130000000
0!
0%
#759135000000
1!
1%
#759140000000
0!
0%
#759145000000
1!
1%
#759150000000
0!
0%
#759155000000
1!
1%
#759160000000
0!
0%
#759165000000
1!
1%
#759170000000
0!
0%
#759175000000
1!
1%
#759180000000
0!
0%
#759185000000
1!
1%
#759190000000
0!
0%
#759195000000
1!
1%
#759200000000
0!
0%
#759205000000
1!
1%
#759210000000
0!
0%
#759215000000
1!
1%
#759220000000
0!
0%
#759225000000
1!
1%
#759230000000
0!
0%
#759235000000
1!
1%
#759240000000
0!
0%
#759245000000
1!
1%
#759250000000
0!
0%
#759255000000
1!
1%
#759260000000
0!
0%
#759265000000
1!
1%
#759270000000
0!
0%
#759275000000
1!
1%
#759280000000
0!
0%
#759285000000
1!
1%
#759290000000
0!
0%
#759295000000
1!
1%
#759300000000
0!
0%
#759305000000
1!
1%
#759310000000
0!
0%
#759315000000
1!
1%
#759320000000
0!
0%
#759325000000
1!
1%
#759330000000
0!
0%
#759335000000
1!
1%
#759340000000
0!
0%
#759345000000
1!
1%
#759350000000
0!
0%
#759355000000
1!
1%
#759360000000
0!
0%
#759365000000
1!
1%
#759370000000
0!
0%
#759375000000
1!
1%
#759380000000
0!
0%
#759385000000
1!
1%
#759390000000
0!
0%
#759395000000
1!
1%
#759400000000
0!
0%
#759405000000
1!
1%
#759410000000
0!
0%
#759415000000
1!
1%
#759420000000
0!
0%
#759425000000
1!
1%
#759430000000
0!
0%
#759435000000
1!
1%
#759440000000
0!
0%
#759445000000
1!
1%
#759450000000
0!
0%
#759455000000
1!
1%
#759460000000
0!
0%
#759465000000
1!
1%
#759470000000
0!
0%
#759475000000
1!
1%
#759480000000
0!
0%
#759485000000
1!
1%
#759490000000
0!
0%
#759495000000
1!
1%
#759500000000
0!
0%
#759505000000
1!
1%
#759510000000
0!
0%
#759515000000
1!
1%
#759520000000
0!
0%
#759525000000
1!
1%
#759530000000
0!
0%
#759535000000
1!
1%
#759540000000
0!
0%
#759545000000
1!
1%
#759550000000
0!
0%
#759555000000
1!
1%
#759560000000
0!
0%
#759565000000
1!
1%
#759570000000
0!
0%
#759575000000
1!
1%
#759580000000
0!
0%
#759585000000
1!
1%
#759590000000
0!
0%
#759595000000
1!
1%
#759600000000
0!
0%
#759605000000
1!
1%
#759610000000
0!
0%
#759615000000
1!
1%
#759620000000
0!
0%
#759625000000
1!
1%
#759630000000
0!
0%
#759635000000
1!
1%
#759640000000
0!
0%
#759645000000
1!
1%
#759650000000
0!
0%
#759655000000
1!
1%
#759660000000
0!
0%
#759665000000
1!
1%
#759670000000
0!
0%
#759675000000
1!
1%
#759680000000
0!
0%
#759685000000
1!
1%
#759690000000
0!
0%
#759695000000
1!
1%
#759700000000
0!
0%
#759705000000
1!
1%
#759710000000
0!
0%
#759715000000
1!
1%
#759720000000
0!
0%
#759725000000
1!
1%
#759730000000
0!
0%
#759735000000
1!
1%
#759740000000
0!
0%
#759745000000
1!
1%
#759750000000
0!
0%
#759755000000
1!
1%
#759760000000
0!
0%
#759765000000
1!
1%
#759770000000
0!
0%
#759775000000
1!
1%
#759780000000
0!
0%
#759785000000
1!
1%
#759790000000
0!
0%
#759795000000
1!
1%
#759800000000
0!
0%
#759805000000
1!
1%
#759810000000
0!
0%
#759815000000
1!
1%
#759820000000
0!
0%
#759825000000
1!
1%
#759830000000
0!
0%
#759835000000
1!
1%
#759840000000
0!
0%
#759845000000
1!
1%
#759850000000
0!
0%
#759855000000
1!
1%
#759860000000
0!
0%
#759865000000
1!
1%
#759870000000
0!
0%
#759875000000
1!
1%
#759880000000
0!
0%
#759885000000
1!
1%
#759890000000
0!
0%
#759895000000
1!
1%
#759900000000
0!
0%
#759905000000
1!
1%
#759910000000
0!
0%
#759915000000
1!
1%
#759920000000
0!
0%
#759925000000
1!
1%
#759930000000
0!
0%
#759935000000
1!
1%
#759940000000
0!
0%
#759945000000
1!
1%
#759950000000
0!
0%
#759955000000
1!
1%
#759960000000
0!
0%
#759965000000
1!
1%
#759970000000
0!
0%
#759975000000
1!
1%
#759980000000
0!
0%
#759985000000
1!
1%
#759990000000
0!
0%
#759995000000
1!
1%
#760000000000
0!
0%
#760005000000
1!
1%
#760010000000
0!
0%
#760015000000
1!
1%
#760020000000
0!
0%
#760025000000
1!
1%
#760030000000
0!
0%
#760035000000
1!
1%
#760040000000
0!
0%
#760045000000
1!
1%
#760050000000
0!
0%
#760055000000
1!
1%
#760060000000
0!
0%
#760065000000
1!
1%
#760070000000
0!
0%
#760075000000
1!
1%
#760080000000
0!
0%
#760085000000
1!
1%
#760090000000
0!
0%
#760095000000
1!
1%
#760100000000
0!
0%
#760105000000
1!
1%
#760110000000
0!
0%
#760115000000
1!
1%
#760120000000
0!
0%
#760125000000
1!
1%
#760130000000
0!
0%
#760135000000
1!
1%
#760140000000
0!
0%
#760145000000
1!
1%
#760150000000
0!
0%
#760155000000
1!
1%
#760160000000
0!
0%
#760165000000
1!
1%
#760170000000
0!
0%
#760175000000
1!
1%
#760180000000
0!
0%
#760185000000
1!
1%
#760190000000
0!
0%
#760195000000
1!
1%
#760200000000
0!
0%
#760205000000
1!
1%
#760210000000
0!
0%
#760215000000
1!
1%
#760220000000
0!
0%
#760225000000
1!
1%
#760230000000
0!
0%
#760235000000
1!
1%
#760240000000
0!
0%
#760245000000
1!
1%
#760250000000
0!
0%
#760255000000
1!
1%
#760260000000
0!
0%
#760265000000
1!
1%
#760270000000
0!
0%
#760275000000
1!
1%
#760280000000
0!
0%
#760285000000
1!
1%
#760290000000
0!
0%
#760295000000
1!
1%
#760300000000
0!
0%
#760305000000
1!
1%
#760310000000
0!
0%
#760315000000
1!
1%
#760320000000
0!
0%
#760325000000
1!
1%
#760330000000
0!
0%
#760335000000
1!
1%
#760340000000
0!
0%
#760345000000
1!
1%
#760350000000
0!
0%
#760355000000
1!
1%
#760360000000
0!
0%
#760365000000
1!
1%
#760370000000
0!
0%
#760375000000
1!
1%
#760380000000
0!
0%
#760385000000
1!
1%
#760390000000
0!
0%
#760395000000
1!
1%
#760400000000
0!
0%
#760405000000
1!
1%
#760410000000
0!
0%
#760415000000
1!
1%
#760420000000
0!
0%
#760425000000
1!
1%
#760430000000
0!
0%
#760435000000
1!
1%
#760440000000
0!
0%
#760445000000
1!
1%
#760450000000
0!
0%
#760455000000
1!
1%
#760460000000
0!
0%
#760465000000
1!
1%
#760470000000
0!
0%
#760475000000
1!
1%
#760480000000
0!
0%
#760485000000
1!
1%
#760490000000
0!
0%
#760495000000
1!
1%
#760500000000
0!
0%
#760505000000
1!
1%
#760510000000
0!
0%
#760515000000
1!
1%
#760520000000
0!
0%
#760525000000
1!
1%
#760530000000
0!
0%
#760535000000
1!
1%
#760540000000
0!
0%
#760545000000
1!
1%
#760550000000
0!
0%
#760555000000
1!
1%
#760560000000
0!
0%
#760565000000
1!
1%
#760570000000
0!
0%
#760575000000
1!
1%
#760580000000
0!
0%
#760585000000
1!
1%
#760590000000
0!
0%
#760595000000
1!
1%
#760600000000
0!
0%
#760605000000
1!
1%
#760610000000
0!
0%
#760615000000
1!
1%
#760620000000
0!
0%
#760625000000
1!
1%
#760630000000
0!
0%
#760635000000
1!
1%
#760640000000
0!
0%
#760645000000
1!
1%
#760650000000
0!
0%
#760655000000
1!
1%
#760660000000
0!
0%
#760665000000
1!
1%
#760670000000
0!
0%
#760675000000
1!
1%
#760680000000
0!
0%
#760685000000
1!
1%
#760690000000
0!
0%
#760695000000
1!
1%
#760700000000
0!
0%
#760705000000
1!
1%
#760710000000
0!
0%
#760715000000
1!
1%
#760720000000
0!
0%
#760725000000
1!
1%
#760730000000
0!
0%
#760735000000
1!
1%
#760740000000
0!
0%
#760745000000
1!
1%
#760750000000
0!
0%
#760755000000
1!
1%
#760760000000
0!
0%
#760765000000
1!
1%
#760770000000
0!
0%
#760775000000
1!
1%
#760780000000
0!
0%
#760785000000
1!
1%
#760790000000
0!
0%
#760795000000
1!
1%
#760800000000
0!
0%
#760805000000
1!
1%
#760810000000
0!
0%
#760815000000
1!
1%
#760820000000
0!
0%
#760825000000
1!
1%
#760830000000
0!
0%
#760835000000
1!
1%
#760840000000
0!
0%
#760845000000
1!
1%
#760850000000
0!
0%
#760855000000
1!
1%
#760860000000
0!
0%
#760865000000
1!
1%
#760870000000
0!
0%
#760875000000
1!
1%
#760880000000
0!
0%
#760885000000
1!
1%
#760890000000
0!
0%
#760895000000
1!
1%
#760900000000
0!
0%
#760905000000
1!
1%
#760910000000
0!
0%
#760915000000
1!
1%
#760920000000
0!
0%
#760925000000
1!
1%
#760930000000
0!
0%
#760935000000
1!
1%
#760940000000
0!
0%
#760945000000
1!
1%
#760950000000
0!
0%
#760955000000
1!
1%
#760960000000
0!
0%
#760965000000
1!
1%
#760970000000
0!
0%
#760975000000
1!
1%
#760980000000
0!
0%
#760985000000
1!
1%
#760990000000
0!
0%
#760995000000
1!
1%
#761000000000
0!
0%
#761005000000
1!
1%
#761010000000
0!
0%
#761015000000
1!
1%
#761020000000
0!
0%
#761025000000
1!
1%
#761030000000
0!
0%
#761035000000
1!
1%
#761040000000
0!
0%
#761045000000
1!
1%
#761050000000
0!
0%
#761055000000
1!
1%
#761060000000
0!
0%
#761065000000
1!
1%
#761070000000
0!
0%
#761075000000
1!
1%
#761080000000
0!
0%
#761085000000
1!
1%
#761090000000
0!
0%
#761095000000
1!
1%
#761100000000
0!
0%
#761105000000
1!
1%
#761110000000
0!
0%
#761115000000
1!
1%
#761120000000
0!
0%
#761125000000
1!
1%
#761130000000
0!
0%
#761135000000
1!
1%
#761140000000
0!
0%
#761145000000
1!
1%
#761150000000
0!
0%
#761155000000
1!
1%
#761160000000
0!
0%
#761165000000
1!
1%
#761170000000
0!
0%
#761175000000
1!
1%
#761180000000
0!
0%
#761185000000
1!
1%
#761190000000
0!
0%
#761195000000
1!
1%
#761200000000
0!
0%
#761205000000
1!
1%
#761210000000
0!
0%
#761215000000
1!
1%
#761220000000
0!
0%
#761225000000
1!
1%
#761230000000
0!
0%
#761235000000
1!
1%
#761240000000
0!
0%
#761245000000
1!
1%
#761250000000
0!
0%
#761255000000
1!
1%
#761260000000
0!
0%
#761265000000
1!
1%
#761270000000
0!
0%
#761275000000
1!
1%
#761280000000
0!
0%
#761285000000
1!
1%
#761290000000
0!
0%
#761295000000
1!
1%
#761300000000
0!
0%
#761305000000
1!
1%
#761310000000
0!
0%
#761315000000
1!
1%
#761320000000
0!
0%
#761325000000
1!
1%
#761330000000
0!
0%
#761335000000
1!
1%
#761340000000
0!
0%
#761345000000
1!
1%
#761350000000
0!
0%
#761355000000
1!
1%
#761360000000
0!
0%
#761365000000
1!
1%
#761370000000
0!
0%
#761375000000
1!
1%
#761380000000
0!
0%
#761385000000
1!
1%
#761390000000
0!
0%
#761395000000
1!
1%
#761400000000
0!
0%
#761405000000
1!
1%
#761410000000
0!
0%
#761415000000
1!
1%
#761420000000
0!
0%
#761425000000
1!
1%
#761430000000
0!
0%
#761435000000
1!
1%
#761440000000
0!
0%
#761445000000
1!
1%
#761450000000
0!
0%
#761455000000
1!
1%
#761460000000
0!
0%
#761465000000
1!
1%
#761470000000
0!
0%
#761475000000
1!
1%
#761480000000
0!
0%
#761485000000
1!
1%
#761490000000
0!
0%
#761495000000
1!
1%
#761500000000
0!
0%
#761505000000
1!
1%
#761510000000
0!
0%
#761515000000
1!
1%
#761520000000
0!
0%
#761525000000
1!
1%
#761530000000
0!
0%
#761535000000
1!
1%
#761540000000
0!
0%
#761545000000
1!
1%
#761550000000
0!
0%
#761555000000
1!
1%
#761560000000
0!
0%
#761565000000
1!
1%
#761570000000
0!
0%
#761575000000
1!
1%
#761580000000
0!
0%
#761585000000
1!
1%
#761590000000
0!
0%
#761595000000
1!
1%
#761600000000
0!
0%
#761605000000
1!
1%
#761610000000
0!
0%
#761615000000
1!
1%
#761620000000
0!
0%
#761625000000
1!
1%
#761630000000
0!
0%
#761635000000
1!
1%
#761640000000
0!
0%
#761645000000
1!
1%
#761650000000
0!
0%
#761655000000
1!
1%
#761660000000
0!
0%
#761665000000
1!
1%
#761670000000
0!
0%
#761675000000
1!
1%
#761680000000
0!
0%
#761685000000
1!
1%
#761690000000
0!
0%
#761695000000
1!
1%
#761700000000
0!
0%
#761705000000
1!
1%
#761710000000
0!
0%
#761715000000
1!
1%
#761720000000
0!
0%
#761725000000
1!
1%
#761730000000
0!
0%
#761735000000
1!
1%
#761740000000
0!
0%
#761745000000
1!
1%
#761750000000
0!
0%
#761755000000
1!
1%
#761760000000
0!
0%
#761765000000
1!
1%
#761770000000
0!
0%
#761775000000
1!
1%
#761780000000
0!
0%
#761785000000
1!
1%
#761790000000
0!
0%
#761795000000
1!
1%
#761800000000
0!
0%
#761805000000
1!
1%
#761810000000
0!
0%
#761815000000
1!
1%
#761820000000
0!
0%
#761825000000
1!
1%
#761830000000
0!
0%
#761835000000
1!
1%
#761840000000
0!
0%
#761845000000
1!
1%
#761850000000
0!
0%
#761855000000
1!
1%
#761860000000
0!
0%
#761865000000
1!
1%
#761870000000
0!
0%
#761875000000
1!
1%
#761880000000
0!
0%
#761885000000
1!
1%
#761890000000
0!
0%
#761895000000
1!
1%
#761900000000
0!
0%
#761905000000
1!
1%
#761910000000
0!
0%
#761915000000
1!
1%
#761920000000
0!
0%
#761925000000
1!
1%
#761930000000
0!
0%
#761935000000
1!
1%
#761940000000
0!
0%
#761945000000
1!
1%
#761950000000
0!
0%
#761955000000
1!
1%
#761960000000
0!
0%
#761965000000
1!
1%
#761970000000
0!
0%
#761975000000
1!
1%
#761980000000
0!
0%
#761985000000
1!
1%
#761990000000
0!
0%
#761995000000
1!
1%
#762000000000
0!
0%
#762005000000
1!
1%
#762010000000
0!
0%
#762015000000
1!
1%
#762020000000
0!
0%
#762025000000
1!
1%
#762030000000
0!
0%
#762035000000
1!
1%
#762040000000
0!
0%
#762045000000
1!
1%
#762050000000
0!
0%
#762055000000
1!
1%
#762060000000
0!
0%
#762065000000
1!
1%
#762070000000
0!
0%
#762075000000
1!
1%
#762080000000
0!
0%
#762085000000
1!
1%
#762090000000
0!
0%
#762095000000
1!
1%
#762100000000
0!
0%
#762105000000
1!
1%
#762110000000
0!
0%
#762115000000
1!
1%
#762120000000
0!
0%
#762125000000
1!
1%
#762130000000
0!
0%
#762135000000
1!
1%
#762140000000
0!
0%
#762145000000
1!
1%
#762150000000
0!
0%
#762155000000
1!
1%
#762160000000
0!
0%
#762165000000
1!
1%
#762170000000
0!
0%
#762175000000
1!
1%
#762180000000
0!
0%
#762185000000
1!
1%
#762190000000
0!
0%
#762195000000
1!
1%
#762200000000
0!
0%
#762205000000
1!
1%
#762210000000
0!
0%
#762215000000
1!
1%
#762220000000
0!
0%
#762225000000
1!
1%
#762230000000
0!
0%
#762235000000
1!
1%
#762240000000
0!
0%
#762245000000
1!
1%
#762250000000
0!
0%
#762255000000
1!
1%
#762260000000
0!
0%
#762265000000
1!
1%
#762270000000
0!
0%
#762275000000
1!
1%
#762280000000
0!
0%
#762285000000
1!
1%
#762290000000
0!
0%
#762295000000
1!
1%
#762300000000
0!
0%
#762305000000
1!
1%
#762310000000
0!
0%
#762315000000
1!
1%
#762320000000
0!
0%
#762325000000
1!
1%
#762330000000
0!
0%
#762335000000
1!
1%
#762340000000
0!
0%
#762345000000
1!
1%
#762350000000
0!
0%
#762355000000
1!
1%
#762360000000
0!
0%
#762365000000
1!
1%
#762370000000
0!
0%
#762375000000
1!
1%
#762380000000
0!
0%
#762385000000
1!
1%
#762390000000
0!
0%
#762395000000
1!
1%
#762400000000
0!
0%
#762405000000
1!
1%
#762410000000
0!
0%
#762415000000
1!
1%
#762420000000
0!
0%
#762425000000
1!
1%
#762430000000
0!
0%
#762435000000
1!
1%
#762440000000
0!
0%
#762445000000
1!
1%
#762450000000
0!
0%
#762455000000
1!
1%
#762460000000
0!
0%
#762465000000
1!
1%
#762470000000
0!
0%
#762475000000
1!
1%
#762480000000
0!
0%
#762485000000
1!
1%
#762490000000
0!
0%
#762495000000
1!
1%
#762500000000
0!
0%
#762505000000
1!
1%
#762510000000
0!
0%
#762515000000
1!
1%
#762520000000
0!
0%
#762525000000
1!
1%
#762530000000
0!
0%
#762535000000
1!
1%
#762540000000
0!
0%
#762545000000
1!
1%
#762550000000
0!
0%
#762555000000
1!
1%
#762560000000
0!
0%
#762565000000
1!
1%
#762570000000
0!
0%
#762575000000
1!
1%
#762580000000
0!
0%
#762585000000
1!
1%
#762590000000
0!
0%
#762595000000
1!
1%
#762600000000
0!
0%
#762605000000
1!
1%
#762610000000
0!
0%
#762615000000
1!
1%
#762620000000
0!
0%
#762625000000
1!
1%
#762630000000
0!
0%
#762635000000
1!
1%
#762640000000
0!
0%
#762645000000
1!
1%
#762650000000
0!
0%
#762655000000
1!
1%
#762660000000
0!
0%
#762665000000
1!
1%
#762670000000
0!
0%
#762675000000
1!
1%
#762680000000
0!
0%
#762685000000
1!
1%
#762690000000
0!
0%
#762695000000
1!
1%
#762700000000
0!
0%
#762705000000
1!
1%
#762710000000
0!
0%
#762715000000
1!
1%
#762720000000
0!
0%
#762725000000
1!
1%
#762730000000
0!
0%
#762735000000
1!
1%
#762740000000
0!
0%
#762745000000
1!
1%
#762750000000
0!
0%
#762755000000
1!
1%
#762760000000
0!
0%
#762765000000
1!
1%
#762770000000
0!
0%
#762775000000
1!
1%
#762780000000
0!
0%
#762785000000
1!
1%
#762790000000
0!
0%
#762795000000
1!
1%
#762800000000
0!
0%
#762805000000
1!
1%
#762810000000
0!
0%
#762815000000
1!
1%
#762820000000
0!
0%
#762825000000
1!
1%
#762830000000
0!
0%
#762835000000
1!
1%
#762840000000
0!
0%
#762845000000
1!
1%
#762850000000
0!
0%
#762855000000
1!
1%
#762860000000
0!
0%
#762865000000
1!
1%
#762870000000
0!
0%
#762875000000
1!
1%
#762880000000
0!
0%
#762885000000
1!
1%
#762890000000
0!
0%
#762895000000
1!
1%
#762900000000
0!
0%
#762905000000
1!
1%
#762910000000
0!
0%
#762915000000
1!
1%
#762920000000
0!
0%
#762925000000
1!
1%
#762930000000
0!
0%
#762935000000
1!
1%
#762940000000
0!
0%
#762945000000
1!
1%
#762950000000
0!
0%
#762955000000
1!
1%
#762960000000
0!
0%
#762965000000
1!
1%
#762970000000
0!
0%
#762975000000
1!
1%
#762980000000
0!
0%
#762985000000
1!
1%
#762990000000
0!
0%
#762995000000
1!
1%
#763000000000
0!
0%
#763005000000
1!
1%
#763010000000
0!
0%
#763015000000
1!
1%
#763020000000
0!
0%
#763025000000
1!
1%
#763030000000
0!
0%
#763035000000
1!
1%
#763040000000
0!
0%
#763045000000
1!
1%
#763050000000
0!
0%
#763055000000
1!
1%
#763060000000
0!
0%
#763065000000
1!
1%
#763070000000
0!
0%
#763075000000
1!
1%
#763080000000
0!
0%
#763085000000
1!
1%
#763090000000
0!
0%
#763095000000
1!
1%
#763100000000
0!
0%
#763105000000
1!
1%
#763110000000
0!
0%
#763115000000
1!
1%
#763120000000
0!
0%
#763125000000
1!
1%
#763130000000
0!
0%
#763135000000
1!
1%
#763140000000
0!
0%
#763145000000
1!
1%
#763150000000
0!
0%
#763155000000
1!
1%
#763160000000
0!
0%
#763165000000
1!
1%
#763170000000
0!
0%
#763175000000
1!
1%
#763180000000
0!
0%
#763185000000
1!
1%
#763190000000
0!
0%
#763195000000
1!
1%
#763200000000
0!
0%
#763205000000
1!
1%
#763210000000
0!
0%
#763215000000
1!
1%
#763220000000
0!
0%
#763225000000
1!
1%
#763230000000
0!
0%
#763235000000
1!
1%
#763240000000
0!
0%
#763245000000
1!
1%
#763250000000
0!
0%
#763255000000
1!
1%
#763260000000
0!
0%
#763265000000
1!
1%
#763270000000
0!
0%
#763275000000
1!
1%
#763280000000
0!
0%
#763285000000
1!
1%
#763290000000
0!
0%
#763295000000
1!
1%
#763300000000
0!
0%
#763305000000
1!
1%
#763310000000
0!
0%
#763315000000
1!
1%
#763320000000
0!
0%
#763325000000
1!
1%
#763330000000
0!
0%
#763335000000
1!
1%
#763340000000
0!
0%
#763345000000
1!
1%
#763350000000
0!
0%
#763355000000
1!
1%
#763360000000
0!
0%
#763365000000
1!
1%
#763370000000
0!
0%
#763375000000
1!
1%
#763380000000
0!
0%
#763385000000
1!
1%
#763390000000
0!
0%
#763395000000
1!
1%
#763400000000
0!
0%
#763405000000
1!
1%
#763410000000
0!
0%
#763415000000
1!
1%
#763420000000
0!
0%
#763425000000
1!
1%
#763430000000
0!
0%
#763435000000
1!
1%
#763440000000
0!
0%
#763445000000
1!
1%
#763450000000
0!
0%
#763455000000
1!
1%
#763460000000
0!
0%
#763465000000
1!
1%
#763470000000
0!
0%
#763475000000
1!
1%
#763480000000
0!
0%
#763485000000
1!
1%
#763490000000
0!
0%
#763495000000
1!
1%
#763500000000
0!
0%
#763505000000
1!
1%
#763510000000
0!
0%
#763515000000
1!
1%
#763520000000
0!
0%
#763525000000
1!
1%
#763530000000
0!
0%
#763535000000
1!
1%
#763540000000
0!
0%
#763545000000
1!
1%
#763550000000
0!
0%
#763555000000
1!
1%
#763560000000
0!
0%
#763565000000
1!
1%
#763570000000
0!
0%
#763575000000
1!
1%
#763580000000
0!
0%
#763585000000
1!
1%
#763590000000
0!
0%
#763595000000
1!
1%
#763600000000
0!
0%
#763605000000
1!
1%
#763610000000
0!
0%
#763615000000
1!
1%
#763620000000
0!
0%
#763625000000
1!
1%
#763630000000
0!
0%
#763635000000
1!
1%
#763640000000
0!
0%
#763645000000
1!
1%
#763650000000
0!
0%
#763655000000
1!
1%
#763660000000
0!
0%
#763665000000
1!
1%
#763670000000
0!
0%
#763675000000
1!
1%
#763680000000
0!
0%
#763685000000
1!
1%
#763690000000
0!
0%
#763695000000
1!
1%
#763700000000
0!
0%
#763705000000
1!
1%
#763710000000
0!
0%
#763715000000
1!
1%
#763720000000
0!
0%
#763725000000
1!
1%
#763730000000
0!
0%
#763735000000
1!
1%
#763740000000
0!
0%
#763745000000
1!
1%
#763750000000
0!
0%
#763755000000
1!
1%
#763760000000
0!
0%
#763765000000
1!
1%
#763770000000
0!
0%
#763775000000
1!
1%
#763780000000
0!
0%
#763785000000
1!
1%
#763790000000
0!
0%
#763795000000
1!
1%
#763800000000
0!
0%
#763805000000
1!
1%
#763810000000
0!
0%
#763815000000
1!
1%
#763820000000
0!
0%
#763825000000
1!
1%
#763830000000
0!
0%
#763835000000
1!
1%
#763840000000
0!
0%
#763845000000
1!
1%
#763850000000
0!
0%
#763855000000
1!
1%
#763860000000
0!
0%
#763865000000
1!
1%
#763870000000
0!
0%
#763875000000
1!
1%
#763880000000
0!
0%
#763885000000
1!
1%
#763890000000
0!
0%
#763895000000
1!
1%
#763900000000
0!
0%
#763905000000
1!
1%
#763910000000
0!
0%
#763915000000
1!
1%
#763920000000
0!
0%
#763925000000
1!
1%
#763930000000
0!
0%
#763935000000
1!
1%
#763940000000
0!
0%
#763945000000
1!
1%
#763950000000
0!
0%
#763955000000
1!
1%
#763960000000
0!
0%
#763965000000
1!
1%
#763970000000
0!
0%
#763975000000
1!
1%
#763980000000
0!
0%
#763985000000
1!
1%
#763990000000
0!
0%
#763995000000
1!
1%
#764000000000
0!
0%
#764005000000
1!
1%
#764010000000
0!
0%
#764015000000
1!
1%
#764020000000
0!
0%
#764025000000
1!
1%
#764030000000
0!
0%
#764035000000
1!
1%
#764040000000
0!
0%
#764045000000
1!
1%
#764050000000
0!
0%
#764055000000
1!
1%
#764060000000
0!
0%
#764065000000
1!
1%
#764070000000
0!
0%
#764075000000
1!
1%
#764080000000
0!
0%
#764085000000
1!
1%
#764090000000
0!
0%
#764095000000
1!
1%
#764100000000
0!
0%
#764105000000
1!
1%
#764110000000
0!
0%
#764115000000
1!
1%
#764120000000
0!
0%
#764125000000
1!
1%
#764130000000
0!
0%
#764135000000
1!
1%
#764140000000
0!
0%
#764145000000
1!
1%
#764150000000
0!
0%
#764155000000
1!
1%
#764160000000
0!
0%
#764165000000
1!
1%
#764170000000
0!
0%
#764175000000
1!
1%
#764180000000
0!
0%
#764185000000
1!
1%
#764190000000
0!
0%
#764195000000
1!
1%
#764200000000
0!
0%
#764205000000
1!
1%
#764210000000
0!
0%
#764215000000
1!
1%
#764220000000
0!
0%
#764225000000
1!
1%
#764230000000
0!
0%
#764235000000
1!
1%
#764240000000
0!
0%
#764245000000
1!
1%
#764250000000
0!
0%
#764255000000
1!
1%
#764260000000
0!
0%
#764265000000
1!
1%
#764270000000
0!
0%
#764275000000
1!
1%
#764280000000
0!
0%
#764285000000
1!
1%
#764290000000
0!
0%
#764295000000
1!
1%
#764300000000
0!
0%
#764305000000
1!
1%
#764310000000
0!
0%
#764315000000
1!
1%
#764320000000
0!
0%
#764325000000
1!
1%
#764330000000
0!
0%
#764335000000
1!
1%
#764340000000
0!
0%
#764345000000
1!
1%
#764350000000
0!
0%
#764355000000
1!
1%
#764360000000
0!
0%
#764365000000
1!
1%
#764370000000
0!
0%
#764375000000
1!
1%
#764380000000
0!
0%
#764385000000
1!
1%
#764390000000
0!
0%
#764395000000
1!
1%
#764400000000
0!
0%
#764405000000
1!
1%
#764410000000
0!
0%
#764415000000
1!
1%
#764420000000
0!
0%
#764425000000
1!
1%
#764430000000
0!
0%
#764435000000
1!
1%
#764440000000
0!
0%
#764445000000
1!
1%
#764450000000
0!
0%
#764455000000
1!
1%
#764460000000
0!
0%
#764465000000
1!
1%
#764470000000
0!
0%
#764475000000
1!
1%
#764480000000
0!
0%
#764485000000
1!
1%
#764490000000
0!
0%
#764495000000
1!
1%
#764500000000
0!
0%
#764505000000
1!
1%
#764510000000
0!
0%
#764515000000
1!
1%
#764520000000
0!
0%
#764525000000
1!
1%
#764530000000
0!
0%
#764535000000
1!
1%
#764540000000
0!
0%
#764545000000
1!
1%
#764550000000
0!
0%
#764555000000
1!
1%
#764560000000
0!
0%
#764565000000
1!
1%
#764570000000
0!
0%
#764575000000
1!
1%
#764580000000
0!
0%
#764585000000
1!
1%
#764590000000
0!
0%
#764595000000
1!
1%
#764600000000
0!
0%
#764605000000
1!
1%
#764610000000
0!
0%
#764615000000
1!
1%
#764620000000
0!
0%
#764625000000
1!
1%
#764630000000
0!
0%
#764635000000
1!
1%
#764640000000
0!
0%
#764645000000
1!
1%
#764650000000
0!
0%
#764655000000
1!
1%
#764660000000
0!
0%
#764665000000
1!
1%
#764670000000
0!
0%
#764675000000
1!
1%
#764680000000
0!
0%
#764685000000
1!
1%
#764690000000
0!
0%
#764695000000
1!
1%
#764700000000
0!
0%
#764705000000
1!
1%
#764710000000
0!
0%
#764715000000
1!
1%
#764720000000
0!
0%
#764725000000
1!
1%
#764730000000
0!
0%
#764735000000
1!
1%
#764740000000
0!
0%
#764745000000
1!
1%
#764750000000
0!
0%
#764755000000
1!
1%
#764760000000
0!
0%
#764765000000
1!
1%
#764770000000
0!
0%
#764775000000
1!
1%
#764780000000
0!
0%
#764785000000
1!
1%
#764790000000
0!
0%
#764795000000
1!
1%
#764800000000
0!
0%
#764805000000
1!
1%
#764810000000
0!
0%
#764815000000
1!
1%
#764820000000
0!
0%
#764825000000
1!
1%
#764830000000
0!
0%
#764835000000
1!
1%
#764840000000
0!
0%
#764845000000
1!
1%
#764850000000
0!
0%
#764855000000
1!
1%
#764860000000
0!
0%
#764865000000
1!
1%
#764870000000
0!
0%
#764875000000
1!
1%
#764880000000
0!
0%
#764885000000
1!
1%
#764890000000
0!
0%
#764895000000
1!
1%
#764900000000
0!
0%
#764905000000
1!
1%
#764910000000
0!
0%
#764915000000
1!
1%
#764920000000
0!
0%
#764925000000
1!
1%
#764930000000
0!
0%
#764935000000
1!
1%
#764940000000
0!
0%
#764945000000
1!
1%
#764950000000
0!
0%
#764955000000
1!
1%
#764960000000
0!
0%
#764965000000
1!
1%
#764970000000
0!
0%
#764975000000
1!
1%
#764980000000
0!
0%
#764985000000
1!
1%
#764990000000
0!
0%
#764995000000
1!
1%
#765000000000
0!
0%
#765005000000
1!
1%
#765010000000
0!
0%
#765015000000
1!
1%
#765020000000
0!
0%
#765025000000
1!
1%
#765030000000
0!
0%
#765035000000
1!
1%
#765040000000
0!
0%
#765045000000
1!
1%
#765050000000
0!
0%
#765055000000
1!
1%
#765060000000
0!
0%
#765065000000
1!
1%
#765070000000
0!
0%
#765075000000
1!
1%
#765080000000
0!
0%
#765085000000
1!
1%
#765090000000
0!
0%
#765095000000
1!
1%
#765100000000
0!
0%
#765105000000
1!
1%
#765110000000
0!
0%
#765115000000
1!
1%
#765120000000
0!
0%
#765125000000
1!
1%
#765130000000
0!
0%
#765135000000
1!
1%
#765140000000
0!
0%
#765145000000
1!
1%
#765150000000
0!
0%
#765155000000
1!
1%
#765160000000
0!
0%
#765165000000
1!
1%
#765170000000
0!
0%
#765175000000
1!
1%
#765180000000
0!
0%
#765185000000
1!
1%
#765190000000
0!
0%
#765195000000
1!
1%
#765200000000
0!
0%
#765205000000
1!
1%
#765210000000
0!
0%
#765215000000
1!
1%
#765220000000
0!
0%
#765225000000
1!
1%
#765230000000
0!
0%
#765235000000
1!
1%
#765240000000
0!
0%
#765245000000
1!
1%
#765250000000
0!
0%
#765255000000
1!
1%
#765260000000
0!
0%
#765265000000
1!
1%
#765270000000
0!
0%
#765275000000
1!
1%
#765280000000
0!
0%
#765285000000
1!
1%
#765290000000
0!
0%
#765295000000
1!
1%
#765300000000
0!
0%
#765305000000
1!
1%
#765310000000
0!
0%
#765315000000
1!
1%
#765320000000
0!
0%
#765325000000
1!
1%
#765330000000
0!
0%
#765335000000
1!
1%
#765340000000
0!
0%
#765345000000
1!
1%
#765350000000
0!
0%
#765355000000
1!
1%
#765360000000
0!
0%
#765365000000
1!
1%
#765370000000
0!
0%
#765375000000
1!
1%
#765380000000
0!
0%
#765385000000
1!
1%
#765390000000
0!
0%
#765395000000
1!
1%
#765400000000
0!
0%
#765405000000
1!
1%
#765410000000
0!
0%
#765415000000
1!
1%
#765420000000
0!
0%
#765425000000
1!
1%
#765430000000
0!
0%
#765435000000
1!
1%
#765440000000
0!
0%
#765445000000
1!
1%
#765450000000
0!
0%
#765455000000
1!
1%
#765460000000
0!
0%
#765465000000
1!
1%
#765470000000
0!
0%
#765475000000
1!
1%
#765480000000
0!
0%
#765485000000
1!
1%
#765490000000
0!
0%
#765495000000
1!
1%
#765500000000
0!
0%
#765505000000
1!
1%
#765510000000
0!
0%
#765515000000
1!
1%
#765520000000
0!
0%
#765525000000
1!
1%
#765530000000
0!
0%
#765535000000
1!
1%
#765540000000
0!
0%
#765545000000
1!
1%
#765550000000
0!
0%
#765555000000
1!
1%
#765560000000
0!
0%
#765565000000
1!
1%
#765570000000
0!
0%
#765575000000
1!
1%
#765580000000
0!
0%
#765585000000
1!
1%
#765590000000
0!
0%
#765595000000
1!
1%
#765600000000
0!
0%
#765605000000
1!
1%
#765610000000
0!
0%
#765615000000
1!
1%
#765620000000
0!
0%
#765625000000
1!
1%
#765630000000
0!
0%
#765635000000
1!
1%
#765640000000
0!
0%
#765645000000
1!
1%
#765650000000
0!
0%
#765655000000
1!
1%
#765660000000
0!
0%
#765665000000
1!
1%
#765670000000
0!
0%
#765675000000
1!
1%
#765680000000
0!
0%
#765685000000
1!
1%
#765690000000
0!
0%
#765695000000
1!
1%
#765700000000
0!
0%
#765705000000
1!
1%
#765710000000
0!
0%
#765715000000
1!
1%
#765720000000
0!
0%
#765725000000
1!
1%
#765730000000
0!
0%
#765735000000
1!
1%
#765740000000
0!
0%
#765745000000
1!
1%
#765750000000
0!
0%
#765755000000
1!
1%
#765760000000
0!
0%
#765765000000
1!
1%
#765770000000
0!
0%
#765775000000
1!
1%
#765780000000
0!
0%
#765785000000
1!
1%
#765790000000
0!
0%
#765795000000
1!
1%
#765800000000
0!
0%
#765805000000
1!
1%
#765810000000
0!
0%
#765815000000
1!
1%
#765820000000
0!
0%
#765825000000
1!
1%
#765830000000
0!
0%
#765835000000
1!
1%
#765840000000
0!
0%
#765845000000
1!
1%
#765850000000
0!
0%
#765855000000
1!
1%
#765860000000
0!
0%
#765865000000
1!
1%
#765870000000
0!
0%
#765875000000
1!
1%
#765880000000
0!
0%
#765885000000
1!
1%
#765890000000
0!
0%
#765895000000
1!
1%
#765900000000
0!
0%
#765905000000
1!
1%
#765910000000
0!
0%
#765915000000
1!
1%
#765920000000
0!
0%
#765925000000
1!
1%
#765930000000
0!
0%
#765935000000
1!
1%
#765940000000
0!
0%
#765945000000
1!
1%
#765950000000
0!
0%
#765955000000
1!
1%
#765960000000
0!
0%
#765965000000
1!
1%
#765970000000
0!
0%
#765975000000
1!
1%
#765980000000
0!
0%
#765985000000
1!
1%
#765990000000
0!
0%
#765995000000
1!
1%
#766000000000
0!
0%
#766005000000
1!
1%
#766010000000
0!
0%
#766015000000
1!
1%
#766020000000
0!
0%
#766025000000
1!
1%
#766030000000
0!
0%
#766035000000
1!
1%
#766040000000
0!
0%
#766045000000
1!
1%
#766050000000
0!
0%
#766055000000
1!
1%
#766060000000
0!
0%
#766065000000
1!
1%
#766070000000
0!
0%
#766075000000
1!
1%
#766080000000
0!
0%
#766085000000
1!
1%
#766090000000
0!
0%
#766095000000
1!
1%
#766100000000
0!
0%
#766105000000
1!
1%
#766110000000
0!
0%
#766115000000
1!
1%
#766120000000
0!
0%
#766125000000
1!
1%
#766130000000
0!
0%
#766135000000
1!
1%
#766140000000
0!
0%
#766145000000
1!
1%
#766150000000
0!
0%
#766155000000
1!
1%
#766160000000
0!
0%
#766165000000
1!
1%
#766170000000
0!
0%
#766175000000
1!
1%
#766180000000
0!
0%
#766185000000
1!
1%
#766190000000
0!
0%
#766195000000
1!
1%
#766200000000
0!
0%
#766205000000
1!
1%
#766210000000
0!
0%
#766215000000
1!
1%
#766220000000
0!
0%
#766225000000
1!
1%
#766230000000
0!
0%
#766235000000
1!
1%
#766240000000
0!
0%
#766245000000
1!
1%
#766250000000
0!
0%
#766255000000
1!
1%
#766260000000
0!
0%
#766265000000
1!
1%
#766270000000
0!
0%
#766275000000
1!
1%
#766280000000
0!
0%
#766285000000
1!
1%
#766290000000
0!
0%
#766295000000
1!
1%
#766300000000
0!
0%
#766305000000
1!
1%
#766310000000
0!
0%
#766315000000
1!
1%
#766320000000
0!
0%
#766325000000
1!
1%
#766330000000
0!
0%
#766335000000
1!
1%
#766340000000
0!
0%
#766345000000
1!
1%
#766350000000
0!
0%
#766355000000
1!
1%
#766360000000
0!
0%
#766365000000
1!
1%
#766370000000
0!
0%
#766375000000
1!
1%
#766380000000
0!
0%
#766385000000
1!
1%
#766390000000
0!
0%
#766395000000
1!
1%
#766400000000
0!
0%
#766405000000
1!
1%
#766410000000
0!
0%
#766415000000
1!
1%
#766420000000
0!
0%
#766425000000
1!
1%
#766430000000
0!
0%
#766435000000
1!
1%
#766440000000
0!
0%
#766445000000
1!
1%
#766450000000
0!
0%
#766455000000
1!
1%
#766460000000
0!
0%
#766465000000
1!
1%
#766470000000
0!
0%
#766475000000
1!
1%
#766480000000
0!
0%
#766485000000
1!
1%
#766490000000
0!
0%
#766495000000
1!
1%
#766500000000
0!
0%
#766505000000
1!
1%
#766510000000
0!
0%
#766515000000
1!
1%
#766520000000
0!
0%
#766525000000
1!
1%
#766530000000
0!
0%
#766535000000
1!
1%
#766540000000
0!
0%
#766545000000
1!
1%
#766550000000
0!
0%
#766555000000
1!
1%
#766560000000
0!
0%
#766565000000
1!
1%
#766570000000
0!
0%
#766575000000
1!
1%
#766580000000
0!
0%
#766585000000
1!
1%
#766590000000
0!
0%
#766595000000
1!
1%
#766600000000
0!
0%
#766605000000
1!
1%
#766610000000
0!
0%
#766615000000
1!
1%
#766620000000
0!
0%
#766625000000
1!
1%
#766630000000
0!
0%
#766635000000
1!
1%
#766640000000
0!
0%
#766645000000
1!
1%
#766650000000
0!
0%
#766655000000
1!
1%
#766660000000
0!
0%
#766665000000
1!
1%
#766670000000
0!
0%
#766675000000
1!
1%
#766680000000
0!
0%
#766685000000
1!
1%
#766690000000
0!
0%
#766695000000
1!
1%
#766700000000
0!
0%
#766705000000
1!
1%
#766710000000
0!
0%
#766715000000
1!
1%
#766720000000
0!
0%
#766725000000
1!
1%
#766730000000
0!
0%
#766735000000
1!
1%
#766740000000
0!
0%
#766745000000
1!
1%
#766750000000
0!
0%
#766755000000
1!
1%
#766760000000
0!
0%
#766765000000
1!
1%
#766770000000
0!
0%
#766775000000
1!
1%
#766780000000
0!
0%
#766785000000
1!
1%
#766790000000
0!
0%
#766795000000
1!
1%
#766800000000
0!
0%
#766805000000
1!
1%
#766810000000
0!
0%
#766815000000
1!
1%
#766820000000
0!
0%
#766825000000
1!
1%
#766830000000
0!
0%
#766835000000
1!
1%
#766840000000
0!
0%
#766845000000
1!
1%
#766850000000
0!
0%
#766855000000
1!
1%
#766860000000
0!
0%
#766865000000
1!
1%
#766870000000
0!
0%
#766875000000
1!
1%
#766880000000
0!
0%
#766885000000
1!
1%
#766890000000
0!
0%
#766895000000
1!
1%
#766900000000
0!
0%
#766905000000
1!
1%
#766910000000
0!
0%
#766915000000
1!
1%
#766920000000
0!
0%
#766925000000
1!
1%
#766930000000
0!
0%
#766935000000
1!
1%
#766940000000
0!
0%
#766945000000
1!
1%
#766950000000
0!
0%
#766955000000
1!
1%
#766960000000
0!
0%
#766965000000
1!
1%
#766970000000
0!
0%
#766975000000
1!
1%
#766980000000
0!
0%
#766985000000
1!
1%
#766990000000
0!
0%
#766995000000
1!
1%
#767000000000
0!
0%
#767005000000
1!
1%
#767010000000
0!
0%
#767015000000
1!
1%
#767020000000
0!
0%
#767025000000
1!
1%
#767030000000
0!
0%
#767035000000
1!
1%
#767040000000
0!
0%
#767045000000
1!
1%
#767050000000
0!
0%
#767055000000
1!
1%
#767060000000
0!
0%
#767065000000
1!
1%
#767070000000
0!
0%
#767075000000
1!
1%
#767080000000
0!
0%
#767085000000
1!
1%
#767090000000
0!
0%
#767095000000
1!
1%
#767100000000
0!
0%
#767105000000
1!
1%
#767110000000
0!
0%
#767115000000
1!
1%
#767120000000
0!
0%
#767125000000
1!
1%
#767130000000
0!
0%
#767135000000
1!
1%
#767140000000
0!
0%
#767145000000
1!
1%
#767150000000
0!
0%
#767155000000
1!
1%
#767160000000
0!
0%
#767165000000
1!
1%
#767170000000
0!
0%
#767175000000
1!
1%
#767180000000
0!
0%
#767185000000
1!
1%
#767190000000
0!
0%
#767195000000
1!
1%
#767200000000
0!
0%
#767205000000
1!
1%
#767210000000
0!
0%
#767215000000
1!
1%
#767220000000
0!
0%
#767225000000
1!
1%
#767230000000
0!
0%
#767235000000
1!
1%
#767240000000
0!
0%
#767245000000
1!
1%
#767250000000
0!
0%
#767255000000
1!
1%
#767260000000
0!
0%
#767265000000
1!
1%
#767270000000
0!
0%
#767275000000
1!
1%
#767280000000
0!
0%
#767285000000
1!
1%
#767290000000
0!
0%
#767295000000
1!
1%
#767300000000
0!
0%
#767305000000
1!
1%
#767310000000
0!
0%
#767315000000
1!
1%
#767320000000
0!
0%
#767325000000
1!
1%
#767330000000
0!
0%
#767335000000
1!
1%
#767340000000
0!
0%
#767345000000
1!
1%
#767350000000
0!
0%
#767355000000
1!
1%
#767360000000
0!
0%
#767365000000
1!
1%
#767370000000
0!
0%
#767375000000
1!
1%
#767380000000
0!
0%
#767385000000
1!
1%
#767390000000
0!
0%
#767395000000
1!
1%
#767400000000
0!
0%
#767405000000
1!
1%
#767410000000
0!
0%
#767415000000
1!
1%
#767420000000
0!
0%
#767425000000
1!
1%
#767430000000
0!
0%
#767435000000
1!
1%
#767440000000
0!
0%
#767445000000
1!
1%
#767450000000
0!
0%
#767455000000
1!
1%
#767460000000
0!
0%
#767465000000
1!
1%
#767470000000
0!
0%
#767475000000
1!
1%
#767480000000
0!
0%
#767485000000
1!
1%
#767490000000
0!
0%
#767495000000
1!
1%
#767500000000
0!
0%
#767505000000
1!
1%
#767510000000
0!
0%
#767515000000
1!
1%
#767520000000
0!
0%
#767525000000
1!
1%
#767530000000
0!
0%
#767535000000
1!
1%
#767540000000
0!
0%
#767545000000
1!
1%
#767550000000
0!
0%
#767555000000
1!
1%
#767560000000
0!
0%
#767565000000
1!
1%
#767570000000
0!
0%
#767575000000
1!
1%
#767580000000
0!
0%
#767585000000
1!
1%
#767590000000
0!
0%
#767595000000
1!
1%
#767600000000
0!
0%
#767605000000
1!
1%
#767610000000
0!
0%
#767615000000
1!
1%
#767620000000
0!
0%
#767625000000
1!
1%
#767630000000
0!
0%
#767635000000
1!
1%
#767640000000
0!
0%
#767645000000
1!
1%
#767650000000
0!
0%
#767655000000
1!
1%
#767660000000
0!
0%
#767665000000
1!
1%
#767670000000
0!
0%
#767675000000
1!
1%
#767680000000
0!
0%
#767685000000
1!
1%
#767690000000
0!
0%
#767695000000
1!
1%
#767700000000
0!
0%
#767705000000
1!
1%
#767710000000
0!
0%
#767715000000
1!
1%
#767720000000
0!
0%
#767725000000
1!
1%
#767730000000
0!
0%
#767735000000
1!
1%
#767740000000
0!
0%
#767745000000
1!
1%
#767750000000
0!
0%
#767755000000
1!
1%
#767760000000
0!
0%
#767765000000
1!
1%
#767770000000
0!
0%
#767775000000
1!
1%
#767780000000
0!